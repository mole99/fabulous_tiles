magic
tech sky130A
magscale 1 2
timestamp 1740383649
<< viali >>
rect 1777 8585 1811 8619
rect 2145 8585 2179 8619
rect 2513 8585 2547 8619
rect 3065 8585 3099 8619
rect 3433 8585 3467 8619
rect 4169 8585 4203 8619
rect 4537 8585 4571 8619
rect 4905 8585 4939 8619
rect 5273 8585 5307 8619
rect 5641 8585 5675 8619
rect 6009 8585 6043 8619
rect 6745 8585 6779 8619
rect 7113 8585 7147 8619
rect 7481 8585 7515 8619
rect 7849 8585 7883 8619
rect 8217 8585 8251 8619
rect 8585 8585 8619 8619
rect 9321 8585 9355 8619
rect 9689 8585 9723 8619
rect 10057 8585 10091 8619
rect 10425 8585 10459 8619
rect 10793 8585 10827 8619
rect 11161 8585 11195 8619
rect 11897 8585 11931 8619
rect 12265 8585 12299 8619
rect 12633 8585 12667 8619
rect 13001 8585 13035 8619
rect 13461 8585 13495 8619
rect 13829 8585 13863 8619
rect 14565 8585 14599 8619
rect 14933 8585 14967 8619
rect 15301 8585 15335 8619
rect 15669 8585 15703 8619
rect 16037 8585 16071 8619
rect 16405 8585 16439 8619
rect 17141 8585 17175 8619
rect 17785 8585 17819 8619
rect 18153 8585 18187 8619
rect 18889 8585 18923 8619
rect 19625 8585 19659 8619
rect 20177 8585 20211 8619
rect 20545 8585 20579 8619
rect 39957 8585 39991 8619
rect 40509 8585 40543 8619
rect 40877 8585 40911 8619
rect 41245 8585 41279 8619
rect 41613 8585 41647 8619
rect 41981 8585 42015 8619
rect 42625 8585 42659 8619
rect 43361 8585 43395 8619
rect 44465 8585 44499 8619
rect 45569 8585 45603 8619
rect 45937 8585 45971 8619
rect 46673 8585 46707 8619
rect 6561 8517 6595 8551
rect 1961 8449 1995 8483
rect 2329 8449 2363 8483
rect 2697 8449 2731 8483
rect 2881 8449 2915 8483
rect 3249 8449 3283 8483
rect 3617 8449 3651 8483
rect 4353 8449 4387 8483
rect 4721 8449 4755 8483
rect 5089 8449 5123 8483
rect 5457 8449 5491 8483
rect 5825 8449 5859 8483
rect 6193 8449 6227 8483
rect 6929 8449 6963 8483
rect 7297 8449 7331 8483
rect 7665 8449 7699 8483
rect 8033 8449 8067 8483
rect 8401 8449 8435 8483
rect 8769 8449 8803 8483
rect 9505 8449 9539 8483
rect 9873 8449 9907 8483
rect 10241 8449 10275 8483
rect 10609 8449 10643 8483
rect 10977 8449 11011 8483
rect 11345 8449 11379 8483
rect 12081 8449 12115 8483
rect 12449 8449 12483 8483
rect 12817 8449 12851 8483
rect 13185 8449 13219 8483
rect 13277 8449 13311 8483
rect 13645 8449 13679 8483
rect 14381 8449 14415 8483
rect 14749 8449 14783 8483
rect 15117 8449 15151 8483
rect 15485 8449 15519 8483
rect 15853 8449 15887 8483
rect 16221 8449 16255 8483
rect 16957 8449 16991 8483
rect 17601 8449 17635 8483
rect 17969 8449 18003 8483
rect 18337 8449 18371 8483
rect 18705 8449 18739 8483
rect 19085 8449 19119 8483
rect 19809 8449 19843 8483
rect 19993 8449 20027 8483
rect 20361 8449 20395 8483
rect 20729 8449 20763 8483
rect 20913 8449 20947 8483
rect 40141 8449 40175 8483
rect 40325 8449 40359 8483
rect 40693 8449 40727 8483
rect 41061 8449 41095 8483
rect 41429 8449 41463 8483
rect 41797 8449 41831 8483
rect 42441 8449 42475 8483
rect 42809 8449 42843 8483
rect 43177 8449 43211 8483
rect 43545 8449 43579 8483
rect 43913 8449 43947 8483
rect 44281 8449 44315 8483
rect 45017 8449 45051 8483
rect 45385 8449 45419 8483
rect 45753 8449 45787 8483
rect 46121 8449 46155 8483
rect 46489 8449 46523 8483
rect 46857 8449 46891 8483
rect 17417 8313 17451 8347
rect 18521 8313 18555 8347
rect 19993 8313 20027 8347
rect 42993 8313 43027 8347
rect 43729 8313 43763 8347
rect 44097 8313 44131 8347
rect 45201 8313 45235 8347
rect 46305 8313 46339 8347
rect 47041 8313 47075 8347
rect 1593 8041 1627 8075
rect 3985 8041 4019 8075
rect 6561 8041 6595 8075
rect 9137 8041 9171 8075
rect 10793 8041 10827 8075
rect 11345 8041 11379 8075
rect 12357 8041 12391 8075
rect 13093 8041 13127 8075
rect 14381 8041 14415 8075
rect 14749 8041 14783 8075
rect 16957 8041 16991 8075
rect 17325 8041 17359 8075
rect 17785 8041 17819 8075
rect 18153 8041 18187 8075
rect 19441 8041 19475 8075
rect 20177 8041 20211 8075
rect 29837 8041 29871 8075
rect 30205 8041 30239 8075
rect 40509 8041 40543 8075
rect 41613 8041 41647 8075
rect 45293 8041 45327 8075
rect 45661 8041 45695 8075
rect 46765 8041 46799 8075
rect 47133 8041 47167 8075
rect 5365 7973 5399 8007
rect 11069 7973 11103 8007
rect 13921 7973 13955 8007
rect 27077 7973 27111 8007
rect 34253 7973 34287 8007
rect 37013 7973 37047 8007
rect 46029 7973 46063 8007
rect 46397 7973 46431 8007
rect 18521 7905 18555 7939
rect 1777 7837 1811 7871
rect 2421 7837 2455 7871
rect 4169 7837 4203 7871
rect 5181 7837 5215 7871
rect 6745 7837 6779 7871
rect 9321 7837 9355 7871
rect 10793 7837 10827 7871
rect 10885 7837 10919 7871
rect 11161 7837 11195 7871
rect 11897 7837 11931 7871
rect 11989 7837 12023 7871
rect 12534 7837 12568 7871
rect 12817 7837 12851 7871
rect 12909 7837 12943 7871
rect 13553 7837 13587 7871
rect 13737 7837 13771 7871
rect 14197 7837 14231 7871
rect 14565 7837 14599 7871
rect 16773 7837 16807 7871
rect 17141 7837 17175 7871
rect 17969 7837 18003 7871
rect 18337 7837 18371 7871
rect 18705 7837 18739 7871
rect 19349 7837 19383 7871
rect 19625 7837 19659 7871
rect 20085 7837 20119 7871
rect 20361 7837 20395 7871
rect 21557 7837 21591 7871
rect 26249 7837 26283 7871
rect 27261 7837 27295 7871
rect 28457 7837 28491 7871
rect 29745 7837 29779 7871
rect 30021 7837 30055 7871
rect 30297 7837 30331 7871
rect 30389 7837 30423 7871
rect 30849 7837 30883 7871
rect 34437 7837 34471 7871
rect 36829 7837 36863 7871
rect 39681 7837 39715 7871
rect 40693 7837 40727 7871
rect 41705 7837 41739 7871
rect 41797 7837 41831 7871
rect 45109 7837 45143 7871
rect 45477 7837 45511 7871
rect 45845 7837 45879 7871
rect 46213 7837 46247 7871
rect 46581 7837 46615 7871
rect 46949 7837 46983 7871
rect 2237 7769 2271 7803
rect 12173 7701 12207 7735
rect 12817 7701 12851 7735
rect 18429 7701 18463 7735
rect 18797 7701 18831 7735
rect 21741 7701 21775 7735
rect 26065 7701 26099 7735
rect 28273 7701 28307 7735
rect 29561 7701 29595 7735
rect 30573 7701 30607 7735
rect 30665 7701 30699 7735
rect 39497 7701 39531 7735
rect 41981 7701 42015 7735
rect 14657 7497 14691 7531
rect 15669 7497 15703 7531
rect 15945 7497 15979 7531
rect 17141 7497 17175 7531
rect 22017 7497 22051 7531
rect 41981 7497 42015 7531
rect 44557 7497 44591 7531
rect 45293 7497 45327 7531
rect 46581 7497 46615 7531
rect 46949 7497 46983 7531
rect 47317 7497 47351 7531
rect 7757 7429 7791 7463
rect 7941 7429 7975 7463
rect 15117 7429 15151 7463
rect 14473 7361 14507 7395
rect 15301 7361 15335 7395
rect 15493 7361 15527 7395
rect 15761 7361 15795 7395
rect 17325 7361 17359 7395
rect 21833 7361 21867 7395
rect 26617 7361 26651 7395
rect 33517 7361 33551 7395
rect 41705 7361 41739 7395
rect 41797 7361 41831 7395
rect 42533 7361 42567 7395
rect 43361 7361 43395 7395
rect 44373 7361 44407 7395
rect 45109 7361 45143 7395
rect 45385 7361 45419 7395
rect 45661 7361 45695 7395
rect 46029 7361 46063 7395
rect 46397 7361 46431 7395
rect 46765 7361 46799 7395
rect 47133 7361 47167 7395
rect 26433 7225 26467 7259
rect 42717 7225 42751 7259
rect 43545 7225 43579 7259
rect 45569 7225 45603 7259
rect 33333 7157 33367 7191
rect 41613 7157 41647 7191
rect 45845 7157 45879 7191
rect 46213 7157 46247 7191
rect 15485 6749 15519 6783
rect 15577 6749 15611 6783
rect 16221 6749 16255 6783
rect 16313 6749 16347 6783
rect 23489 6749 23523 6783
rect 29377 6749 29411 6783
rect 32505 6749 32539 6783
rect 35541 6749 35575 6783
rect 45661 6749 45695 6783
rect 45845 6749 45879 6783
rect 46121 6749 46155 6783
rect 46489 6749 46523 6783
rect 46857 6749 46891 6783
rect 47225 6749 47259 6783
rect 15761 6613 15795 6647
rect 16497 6613 16531 6647
rect 23673 6613 23707 6647
rect 29193 6613 29227 6647
rect 32321 6613 32355 6647
rect 35357 6613 35391 6647
rect 46029 6613 46063 6647
rect 46305 6613 46339 6647
rect 46673 6613 46707 6647
rect 47041 6613 47075 6647
rect 47409 6613 47443 6647
rect 39681 6409 39715 6443
rect 46949 6409 46983 6443
rect 47317 6409 47351 6443
rect 36369 6341 36403 6375
rect 24685 6273 24719 6307
rect 25421 6273 25455 6307
rect 25513 6273 25547 6307
rect 25973 6273 26007 6307
rect 26433 6273 26467 6307
rect 32965 6273 32999 6307
rect 39865 6273 39899 6307
rect 46397 6273 46431 6307
rect 46765 6273 46799 6307
rect 47133 6273 47167 6307
rect 25697 6137 25731 6171
rect 36185 6137 36219 6171
rect 24501 6069 24535 6103
rect 25329 6069 25363 6103
rect 25789 6069 25823 6103
rect 26249 6069 26283 6103
rect 33149 6069 33183 6103
rect 46581 6069 46615 6103
rect 14473 5865 14507 5899
rect 17785 5865 17819 5899
rect 22477 5865 22511 5899
rect 47409 5865 47443 5899
rect 28825 5797 28859 5831
rect 30205 5797 30239 5831
rect 38945 5797 38979 5831
rect 14565 5661 14599 5695
rect 14749 5661 14783 5695
rect 14933 5661 14967 5695
rect 22661 5661 22695 5695
rect 29009 5661 29043 5695
rect 30389 5661 30423 5695
rect 31677 5661 31711 5695
rect 39129 5661 39163 5695
rect 46857 5661 46891 5695
rect 47225 5661 47259 5695
rect 17509 5593 17543 5627
rect 17693 5593 17727 5627
rect 17417 5525 17451 5559
rect 31493 5525 31527 5559
rect 47041 5525 47075 5559
rect 21833 5321 21867 5355
rect 23673 5321 23707 5355
rect 47317 5321 47351 5355
rect 9229 5253 9263 5287
rect 9413 5185 9447 5219
rect 21557 5185 21591 5219
rect 22017 5185 22051 5219
rect 23857 5185 23891 5219
rect 37749 5185 37783 5219
rect 46765 5185 46799 5219
rect 47133 5185 47167 5219
rect 37565 5117 37599 5151
rect 21373 4981 21407 5015
rect 46949 4981 46983 5015
rect 18061 4777 18095 4811
rect 20085 4777 20119 4811
rect 20453 4777 20487 4811
rect 20821 4709 20855 4743
rect 23213 4709 23247 4743
rect 47409 4709 47443 4743
rect 18245 4573 18279 4607
rect 20177 4573 20211 4607
rect 20269 4573 20303 4607
rect 21005 4573 21039 4607
rect 21465 4573 21499 4607
rect 23305 4573 23339 4607
rect 23397 4573 23431 4607
rect 24961 4573 24995 4607
rect 25053 4573 25087 4607
rect 46857 4573 46891 4607
rect 47225 4573 47259 4607
rect 21281 4437 21315 4471
rect 23581 4437 23615 4471
rect 24869 4437 24903 4471
rect 25237 4437 25271 4471
rect 47041 4437 47075 4471
rect 12725 4097 12759 4131
rect 15853 4097 15887 4131
rect 16865 4097 16899 4131
rect 18061 4097 18095 4131
rect 18245 4097 18279 4131
rect 22661 4097 22695 4131
rect 22753 4097 22787 4131
rect 46765 4097 46799 4131
rect 47133 4097 47167 4131
rect 16681 3961 16715 3995
rect 17969 3961 18003 3995
rect 18429 3961 18463 3995
rect 47317 3961 47351 3995
rect 12541 3893 12575 3927
rect 15669 3893 15703 3927
rect 22569 3893 22603 3927
rect 22937 3893 22971 3927
rect 46949 3893 46983 3927
rect 24777 3689 24811 3723
rect 47409 3621 47443 3655
rect 24961 3553 24995 3587
rect 14289 3485 14323 3519
rect 20177 3485 20211 3519
rect 24593 3485 24627 3519
rect 25145 3485 25179 3519
rect 46857 3485 46891 3519
rect 47225 3485 47259 3519
rect 25053 3417 25087 3451
rect 14105 3349 14139 3383
rect 19993 3349 20027 3383
rect 25329 3349 25363 3383
rect 47041 3349 47075 3383
rect 8861 3145 8895 3179
rect 12817 3145 12851 3179
rect 17693 3145 17727 3179
rect 22109 3145 22143 3179
rect 23121 3145 23155 3179
rect 38761 3145 38795 3179
rect 39681 3145 39715 3179
rect 40509 3145 40543 3179
rect 43269 3145 43303 3179
rect 44005 3145 44039 3179
rect 47317 3145 47351 3179
rect 8769 3077 8803 3111
rect 13093 3077 13127 3111
rect 17785 3077 17819 3111
rect 17969 3077 18003 3111
rect 18153 3077 18187 3111
rect 8217 3009 8251 3043
rect 8401 3009 8435 3043
rect 10885 3009 10919 3043
rect 12725 3009 12759 3043
rect 15761 3009 15795 3043
rect 16773 3009 16807 3043
rect 18705 3009 18739 3043
rect 20177 3009 20211 3043
rect 20269 3009 20303 3043
rect 20821 3009 20855 3043
rect 20913 3009 20947 3043
rect 21925 3009 21959 3043
rect 22753 3009 22787 3043
rect 22937 3009 22971 3043
rect 25329 3009 25363 3043
rect 27261 3009 27295 3043
rect 27537 3009 27571 3043
rect 29285 3009 29319 3043
rect 36553 3009 36587 3043
rect 36737 3009 36771 3043
rect 37289 3009 37323 3043
rect 37473 3009 37507 3043
rect 38577 3009 38611 3043
rect 39497 3009 39531 3043
rect 40325 3009 40359 3043
rect 43085 3009 43119 3043
rect 43821 3009 43855 3043
rect 46765 3009 46799 3043
rect 47133 3009 47167 3043
rect 11069 2941 11103 2975
rect 8585 2873 8619 2907
rect 13277 2873 13311 2907
rect 15945 2873 15979 2907
rect 18889 2873 18923 2907
rect 8125 2805 8159 2839
rect 16865 2805 16899 2839
rect 20085 2805 20119 2839
rect 20453 2805 20487 2839
rect 20729 2805 20763 2839
rect 21097 2805 21131 2839
rect 25513 2805 25547 2839
rect 27445 2805 27479 2839
rect 27721 2805 27755 2839
rect 29469 2805 29503 2839
rect 36921 2805 36955 2839
rect 37657 2805 37691 2839
rect 46949 2805 46983 2839
rect 45845 2601 45879 2635
rect 47317 2533 47351 2567
rect 45661 2397 45695 2431
rect 46029 2397 46063 2431
rect 46397 2397 46431 2431
rect 46765 2397 46799 2431
rect 47133 2397 47167 2431
rect 46213 2261 46247 2295
rect 46581 2261 46615 2295
rect 46949 2261 46983 2295
<< metal1 >>
rect 13538 11160 13544 11212
rect 13596 11200 13602 11212
rect 39482 11200 39488 11212
rect 13596 11172 39488 11200
rect 13596 11160 13602 11172
rect 39482 11160 39488 11172
rect 39540 11160 39546 11212
rect 14918 11092 14924 11144
rect 14976 11132 14982 11144
rect 38746 11132 38752 11144
rect 14976 11104 38752 11132
rect 14976 11092 14982 11104
rect 38746 11092 38752 11104
rect 38804 11092 38810 11144
rect 18230 11024 18236 11076
rect 18288 11064 18294 11076
rect 36538 11064 36544 11076
rect 18288 11036 36544 11064
rect 18288 11024 18294 11036
rect 36538 11024 36544 11036
rect 36596 11024 36602 11076
rect 11790 10956 11796 11008
rect 11848 10996 11854 11008
rect 29178 10996 29184 11008
rect 11848 10968 29184 10996
rect 11848 10956 11854 10968
rect 29178 10956 29184 10968
rect 29236 10956 29242 11008
rect 18322 10888 18328 10940
rect 18380 10928 18386 10940
rect 36170 10928 36176 10940
rect 18380 10900 36176 10928
rect 18380 10888 18386 10900
rect 36170 10888 36176 10900
rect 36228 10888 36234 10940
rect 21910 10684 21916 10736
rect 21968 10724 21974 10736
rect 24026 10724 24032 10736
rect 21968 10696 24032 10724
rect 21968 10684 21974 10696
rect 24026 10684 24032 10696
rect 24084 10684 24090 10736
rect 1302 9324 1308 9376
rect 1360 9364 1366 9376
rect 7650 9364 7656 9376
rect 1360 9336 7656 9364
rect 1360 9324 1366 9336
rect 7650 9324 7656 9336
rect 7708 9324 7714 9376
rect 8754 9324 8760 9376
rect 8812 9364 8818 9376
rect 16850 9364 16856 9376
rect 8812 9336 16856 9364
rect 8812 9324 8818 9336
rect 16850 9324 16856 9336
rect 16908 9324 16914 9376
rect 20254 9364 20260 9376
rect 17052 9336 20260 9364
rect 4338 9256 4344 9308
rect 4396 9296 4402 9308
rect 17052 9296 17080 9336
rect 20254 9324 20260 9336
rect 20312 9324 20318 9376
rect 25774 9296 25780 9308
rect 4396 9268 17080 9296
rect 17236 9268 25780 9296
rect 4396 9256 4402 9268
rect 6270 9188 6276 9240
rect 6328 9228 6334 9240
rect 17236 9228 17264 9268
rect 25774 9256 25780 9268
rect 25832 9256 25838 9308
rect 6328 9200 17264 9228
rect 6328 9188 6334 9200
rect 19150 9188 19156 9240
rect 19208 9228 19214 9240
rect 26786 9228 26792 9240
rect 19208 9200 26792 9228
rect 19208 9188 19214 9200
rect 26786 9188 26792 9200
rect 26844 9188 26850 9240
rect 23382 9160 23388 9172
rect 6748 9132 23388 9160
rect 3510 8984 3516 9036
rect 3568 9024 3574 9036
rect 6748 9024 6776 9132
rect 23382 9120 23388 9132
rect 23440 9120 23446 9172
rect 34422 9120 34428 9172
rect 34480 9160 34486 9172
rect 45554 9160 45560 9172
rect 34480 9132 45560 9160
rect 34480 9120 34486 9132
rect 45554 9120 45560 9132
rect 45612 9120 45618 9172
rect 7006 9052 7012 9104
rect 7064 9092 7070 9104
rect 15470 9092 15476 9104
rect 7064 9064 15476 9092
rect 7064 9052 7070 9064
rect 15470 9052 15476 9064
rect 15528 9052 15534 9104
rect 15654 9052 15660 9104
rect 15712 9092 15718 9104
rect 38378 9092 38384 9104
rect 15712 9064 38384 9092
rect 15712 9052 15718 9064
rect 38378 9052 38384 9064
rect 38436 9052 38442 9104
rect 8478 9024 8484 9036
rect 3568 8996 6776 9024
rect 7576 8996 8484 9024
rect 3568 8984 3574 8996
rect 4706 8916 4712 8968
rect 4764 8956 4770 8968
rect 7576 8956 7604 8996
rect 8478 8984 8484 8996
rect 8536 8984 8542 9036
rect 14550 8984 14556 9036
rect 14608 9024 14614 9036
rect 39114 9024 39120 9036
rect 14608 8996 39120 9024
rect 14608 8984 14614 8996
rect 39114 8984 39120 8996
rect 39172 8984 39178 9036
rect 4764 8928 7604 8956
rect 4764 8916 4770 8928
rect 7650 8916 7656 8968
rect 7708 8956 7714 8968
rect 7708 8928 22094 8956
rect 7708 8916 7714 8928
rect 6178 8848 6184 8900
rect 6236 8888 6242 8900
rect 14642 8888 14648 8900
rect 6236 8860 14648 8888
rect 6236 8848 6242 8860
rect 14642 8848 14648 8860
rect 14700 8848 14706 8900
rect 15470 8848 15476 8900
rect 15528 8888 15534 8900
rect 15746 8888 15752 8900
rect 15528 8860 15752 8888
rect 15528 8848 15534 8860
rect 15746 8848 15752 8860
rect 15804 8848 15810 8900
rect 22066 8888 22094 8928
rect 26786 8916 26792 8968
rect 26844 8956 26850 8968
rect 36906 8956 36912 8968
rect 26844 8928 36912 8956
rect 26844 8916 26850 8928
rect 36906 8916 36912 8928
rect 36964 8916 36970 8968
rect 42886 8916 42892 8968
rect 42944 8956 42950 8968
rect 46566 8956 46572 8968
rect 42944 8928 46572 8956
rect 42944 8916 42950 8928
rect 46566 8916 46572 8928
rect 46624 8916 46630 8968
rect 32398 8888 32404 8900
rect 22066 8860 32404 8888
rect 32398 8848 32404 8860
rect 32456 8848 32462 8900
rect 43254 8848 43260 8900
rect 43312 8888 43318 8900
rect 45462 8888 45468 8900
rect 43312 8860 45468 8888
rect 43312 8848 43318 8860
rect 45462 8848 45468 8860
rect 45520 8848 45526 8900
rect 5074 8780 5080 8832
rect 5132 8820 5138 8832
rect 8662 8820 8668 8832
rect 5132 8792 8668 8820
rect 5132 8780 5138 8792
rect 8662 8780 8668 8792
rect 8720 8780 8726 8832
rect 10226 8780 10232 8832
rect 10284 8820 10290 8832
rect 18966 8820 18972 8832
rect 10284 8792 18972 8820
rect 10284 8780 10290 8792
rect 18966 8780 18972 8792
rect 19024 8780 19030 8832
rect 19702 8780 19708 8832
rect 19760 8820 19766 8832
rect 40494 8820 40500 8832
rect 19760 8792 40500 8820
rect 19760 8780 19766 8792
rect 40494 8780 40500 8792
rect 40552 8780 40558 8832
rect 40770 8780 40776 8832
rect 40828 8820 40834 8832
rect 43714 8820 43720 8832
rect 40828 8792 43720 8820
rect 40828 8780 40834 8792
rect 43714 8780 43720 8792
rect 43772 8780 43778 8832
rect 45370 8780 45376 8832
rect 45428 8820 45434 8832
rect 46382 8820 46388 8832
rect 45428 8792 46388 8820
rect 45428 8780 45434 8792
rect 46382 8780 46388 8792
rect 46440 8780 46446 8832
rect 1104 8730 47840 8752
rect 1104 8678 3010 8730
rect 3062 8678 3074 8730
rect 3126 8678 3138 8730
rect 3190 8678 3202 8730
rect 3254 8678 3266 8730
rect 3318 8678 9010 8730
rect 9062 8678 9074 8730
rect 9126 8678 9138 8730
rect 9190 8678 9202 8730
rect 9254 8678 9266 8730
rect 9318 8678 15010 8730
rect 15062 8678 15074 8730
rect 15126 8678 15138 8730
rect 15190 8678 15202 8730
rect 15254 8678 15266 8730
rect 15318 8678 21010 8730
rect 21062 8678 21074 8730
rect 21126 8678 21138 8730
rect 21190 8678 21202 8730
rect 21254 8678 21266 8730
rect 21318 8678 27010 8730
rect 27062 8678 27074 8730
rect 27126 8678 27138 8730
rect 27190 8678 27202 8730
rect 27254 8678 27266 8730
rect 27318 8678 33010 8730
rect 33062 8678 33074 8730
rect 33126 8678 33138 8730
rect 33190 8678 33202 8730
rect 33254 8678 33266 8730
rect 33318 8678 39010 8730
rect 39062 8678 39074 8730
rect 39126 8678 39138 8730
rect 39190 8678 39202 8730
rect 39254 8678 39266 8730
rect 39318 8678 45010 8730
rect 45062 8678 45074 8730
rect 45126 8678 45138 8730
rect 45190 8678 45202 8730
rect 45254 8678 45266 8730
rect 45318 8678 47840 8730
rect 1104 8656 47840 8678
rect 1765 8619 1823 8625
rect 1765 8585 1777 8619
rect 1811 8616 1823 8619
rect 1946 8616 1952 8628
rect 1811 8588 1952 8616
rect 1811 8585 1823 8588
rect 1765 8579 1823 8585
rect 1946 8576 1952 8588
rect 2004 8576 2010 8628
rect 2133 8619 2191 8625
rect 2133 8585 2145 8619
rect 2179 8616 2191 8619
rect 2314 8616 2320 8628
rect 2179 8588 2320 8616
rect 2179 8585 2191 8588
rect 2133 8579 2191 8585
rect 2314 8576 2320 8588
rect 2372 8576 2378 8628
rect 2501 8619 2559 8625
rect 2501 8585 2513 8619
rect 2547 8616 2559 8619
rect 2682 8616 2688 8628
rect 2547 8588 2688 8616
rect 2547 8585 2559 8588
rect 2501 8579 2559 8585
rect 2682 8576 2688 8588
rect 2740 8576 2746 8628
rect 2866 8576 2872 8628
rect 2924 8616 2930 8628
rect 3053 8619 3111 8625
rect 3053 8616 3065 8619
rect 2924 8588 3065 8616
rect 2924 8576 2930 8588
rect 3053 8585 3065 8588
rect 3099 8585 3111 8619
rect 3053 8579 3111 8585
rect 3418 8576 3424 8628
rect 3476 8576 3482 8628
rect 4154 8576 4160 8628
rect 4212 8576 4218 8628
rect 4522 8576 4528 8628
rect 4580 8576 4586 8628
rect 4890 8576 4896 8628
rect 4948 8576 4954 8628
rect 5258 8576 5264 8628
rect 5316 8576 5322 8628
rect 5626 8576 5632 8628
rect 5684 8576 5690 8628
rect 5994 8576 6000 8628
rect 6052 8576 6058 8628
rect 6178 8616 6184 8628
rect 6104 8588 6184 8616
rect 1949 8483 2007 8489
rect 1949 8449 1961 8483
rect 1995 8449 2007 8483
rect 1949 8443 2007 8449
rect 1964 8276 1992 8443
rect 2314 8440 2320 8492
rect 2372 8440 2378 8492
rect 2590 8440 2596 8492
rect 2648 8480 2654 8492
rect 2685 8483 2743 8489
rect 2685 8480 2697 8483
rect 2648 8452 2697 8480
rect 2648 8440 2654 8452
rect 2685 8449 2697 8452
rect 2731 8449 2743 8483
rect 2685 8443 2743 8449
rect 2869 8483 2927 8489
rect 2869 8449 2881 8483
rect 2915 8480 2927 8483
rect 3237 8483 3295 8489
rect 3237 8480 3249 8483
rect 2915 8452 3249 8480
rect 2915 8449 2927 8452
rect 2869 8443 2927 8449
rect 3237 8449 3249 8452
rect 3283 8480 3295 8483
rect 3510 8480 3516 8492
rect 3283 8452 3516 8480
rect 3283 8449 3295 8452
rect 3237 8443 3295 8449
rect 3510 8440 3516 8452
rect 3568 8440 3574 8492
rect 3605 8483 3663 8489
rect 3605 8449 3617 8483
rect 3651 8449 3663 8483
rect 3605 8443 3663 8449
rect 3620 8344 3648 8443
rect 4338 8440 4344 8492
rect 4396 8440 4402 8492
rect 4706 8440 4712 8492
rect 4764 8440 4770 8492
rect 5074 8440 5080 8492
rect 5132 8440 5138 8492
rect 5445 8483 5503 8489
rect 5445 8449 5457 8483
rect 5491 8449 5503 8483
rect 5445 8443 5503 8449
rect 5813 8483 5871 8489
rect 5813 8449 5825 8483
rect 5859 8480 5871 8483
rect 6104 8480 6132 8588
rect 6178 8576 6184 8588
rect 6236 8576 6242 8628
rect 6730 8576 6736 8628
rect 6788 8576 6794 8628
rect 7098 8576 7104 8628
rect 7156 8576 7162 8628
rect 7466 8576 7472 8628
rect 7524 8576 7530 8628
rect 7834 8576 7840 8628
rect 7892 8576 7898 8628
rect 8202 8576 8208 8628
rect 8260 8576 8266 8628
rect 8570 8576 8576 8628
rect 8628 8576 8634 8628
rect 9309 8619 9367 8625
rect 9309 8585 9321 8619
rect 9355 8616 9367 8619
rect 9398 8616 9404 8628
rect 9355 8588 9404 8616
rect 9355 8585 9367 8588
rect 9309 8579 9367 8585
rect 9398 8576 9404 8588
rect 9456 8576 9462 8628
rect 9674 8576 9680 8628
rect 9732 8576 9738 8628
rect 10042 8576 10048 8628
rect 10100 8576 10106 8628
rect 10410 8576 10416 8628
rect 10468 8576 10474 8628
rect 10778 8576 10784 8628
rect 10836 8576 10842 8628
rect 11146 8576 11152 8628
rect 11204 8576 11210 8628
rect 11882 8576 11888 8628
rect 11940 8576 11946 8628
rect 12250 8576 12256 8628
rect 12308 8576 12314 8628
rect 12618 8576 12624 8628
rect 12676 8576 12682 8628
rect 12986 8576 12992 8628
rect 13044 8576 13050 8628
rect 13354 8576 13360 8628
rect 13412 8616 13418 8628
rect 13449 8619 13507 8625
rect 13449 8616 13461 8619
rect 13412 8588 13461 8616
rect 13412 8576 13418 8588
rect 13449 8585 13461 8588
rect 13495 8585 13507 8619
rect 13449 8579 13507 8585
rect 13722 8576 13728 8628
rect 13780 8616 13786 8628
rect 13817 8619 13875 8625
rect 13817 8616 13829 8619
rect 13780 8588 13829 8616
rect 13780 8576 13786 8588
rect 13817 8585 13829 8588
rect 13863 8585 13875 8619
rect 13817 8579 13875 8585
rect 14458 8576 14464 8628
rect 14516 8616 14522 8628
rect 14553 8619 14611 8625
rect 14553 8616 14565 8619
rect 14516 8588 14565 8616
rect 14516 8576 14522 8588
rect 14553 8585 14565 8588
rect 14599 8585 14611 8619
rect 14553 8579 14611 8585
rect 14826 8576 14832 8628
rect 14884 8616 14890 8628
rect 14921 8619 14979 8625
rect 14921 8616 14933 8619
rect 14884 8588 14933 8616
rect 14884 8576 14890 8588
rect 14921 8585 14933 8588
rect 14967 8585 14979 8619
rect 14921 8579 14979 8585
rect 15289 8619 15347 8625
rect 15289 8585 15301 8619
rect 15335 8616 15347 8619
rect 15378 8616 15384 8628
rect 15335 8588 15384 8616
rect 15335 8585 15347 8588
rect 15289 8579 15347 8585
rect 15378 8576 15384 8588
rect 15436 8576 15442 8628
rect 15562 8576 15568 8628
rect 15620 8616 15626 8628
rect 15657 8619 15715 8625
rect 15657 8616 15669 8619
rect 15620 8588 15669 8616
rect 15620 8576 15626 8588
rect 15657 8585 15669 8588
rect 15703 8585 15715 8619
rect 15657 8579 15715 8585
rect 15930 8576 15936 8628
rect 15988 8616 15994 8628
rect 16025 8619 16083 8625
rect 16025 8616 16037 8619
rect 15988 8588 16037 8616
rect 15988 8576 15994 8588
rect 16025 8585 16037 8588
rect 16071 8585 16083 8619
rect 16025 8579 16083 8585
rect 16298 8576 16304 8628
rect 16356 8616 16362 8628
rect 16393 8619 16451 8625
rect 16393 8616 16405 8619
rect 16356 8588 16405 8616
rect 16356 8576 16362 8588
rect 16393 8585 16405 8588
rect 16439 8585 16451 8619
rect 16393 8579 16451 8585
rect 17129 8619 17187 8625
rect 17129 8585 17141 8619
rect 17175 8616 17187 8619
rect 17402 8616 17408 8628
rect 17175 8588 17408 8616
rect 17175 8585 17187 8588
rect 17129 8579 17187 8585
rect 17402 8576 17408 8588
rect 17460 8576 17466 8628
rect 17773 8619 17831 8625
rect 17773 8585 17785 8619
rect 17819 8616 17831 8619
rect 18046 8616 18052 8628
rect 17819 8588 18052 8616
rect 17819 8585 17831 8588
rect 17773 8579 17831 8585
rect 18046 8576 18052 8588
rect 18104 8576 18110 8628
rect 18141 8619 18199 8625
rect 18141 8585 18153 8619
rect 18187 8616 18199 8619
rect 18506 8616 18512 8628
rect 18187 8588 18512 8616
rect 18187 8585 18199 8588
rect 18141 8579 18199 8585
rect 18506 8576 18512 8588
rect 18564 8576 18570 8628
rect 18877 8619 18935 8625
rect 18877 8585 18889 8619
rect 18923 8616 18935 8619
rect 19242 8616 19248 8628
rect 18923 8588 19248 8616
rect 18923 8585 18935 8588
rect 18877 8579 18935 8585
rect 19242 8576 19248 8588
rect 19300 8576 19306 8628
rect 19610 8576 19616 8628
rect 19668 8576 19674 8628
rect 19702 8576 19708 8628
rect 19760 8576 19766 8628
rect 19978 8576 19984 8628
rect 20036 8616 20042 8628
rect 20165 8619 20223 8625
rect 20165 8616 20177 8619
rect 20036 8588 20177 8616
rect 20036 8576 20042 8588
rect 20165 8585 20177 8588
rect 20211 8585 20223 8619
rect 20165 8579 20223 8585
rect 20346 8576 20352 8628
rect 20404 8616 20410 8628
rect 20533 8619 20591 8625
rect 20533 8616 20545 8619
rect 20404 8588 20545 8616
rect 20404 8576 20410 8588
rect 20533 8585 20545 8588
rect 20579 8585 20591 8619
rect 20533 8579 20591 8585
rect 39850 8576 39856 8628
rect 39908 8616 39914 8628
rect 39945 8619 40003 8625
rect 39945 8616 39957 8619
rect 39908 8588 39957 8616
rect 39908 8576 39914 8588
rect 39945 8585 39957 8588
rect 39991 8585 40003 8619
rect 39945 8579 40003 8585
rect 40218 8576 40224 8628
rect 40276 8616 40282 8628
rect 40497 8619 40555 8625
rect 40497 8616 40509 8619
rect 40276 8588 40509 8616
rect 40276 8576 40282 8588
rect 40497 8585 40509 8588
rect 40543 8585 40555 8619
rect 40497 8579 40555 8585
rect 40586 8576 40592 8628
rect 40644 8616 40650 8628
rect 40865 8619 40923 8625
rect 40865 8616 40877 8619
rect 40644 8588 40877 8616
rect 40644 8576 40650 8588
rect 40865 8585 40877 8588
rect 40911 8585 40923 8619
rect 40865 8579 40923 8585
rect 40954 8576 40960 8628
rect 41012 8616 41018 8628
rect 41233 8619 41291 8625
rect 41233 8616 41245 8619
rect 41012 8588 41245 8616
rect 41012 8576 41018 8588
rect 41233 8585 41245 8588
rect 41279 8585 41291 8619
rect 41233 8579 41291 8585
rect 41322 8576 41328 8628
rect 41380 8616 41386 8628
rect 41601 8619 41659 8625
rect 41601 8616 41613 8619
rect 41380 8588 41613 8616
rect 41380 8576 41386 8588
rect 41601 8585 41613 8588
rect 41647 8585 41659 8619
rect 41601 8579 41659 8585
rect 41690 8576 41696 8628
rect 41748 8616 41754 8628
rect 41969 8619 42027 8625
rect 41969 8616 41981 8619
rect 41748 8588 41981 8616
rect 41748 8576 41754 8588
rect 41969 8585 41981 8588
rect 42015 8585 42027 8619
rect 41969 8579 42027 8585
rect 42058 8576 42064 8628
rect 42116 8616 42122 8628
rect 42613 8619 42671 8625
rect 42613 8616 42625 8619
rect 42116 8588 42625 8616
rect 42116 8576 42122 8588
rect 42613 8585 42625 8588
rect 42659 8585 42671 8619
rect 42613 8579 42671 8585
rect 42794 8576 42800 8628
rect 42852 8616 42858 8628
rect 43349 8619 43407 8625
rect 43349 8616 43361 8619
rect 42852 8588 43361 8616
rect 42852 8576 42858 8588
rect 43349 8585 43361 8588
rect 43395 8585 43407 8619
rect 43349 8579 43407 8585
rect 43898 8576 43904 8628
rect 43956 8616 43962 8628
rect 44453 8619 44511 8625
rect 44453 8616 44465 8619
rect 43956 8588 44465 8616
rect 43956 8576 43962 8588
rect 44453 8585 44465 8588
rect 44499 8585 44511 8619
rect 44453 8579 44511 8585
rect 44634 8576 44640 8628
rect 44692 8616 44698 8628
rect 45557 8619 45615 8625
rect 45557 8616 45569 8619
rect 44692 8588 45569 8616
rect 44692 8576 44698 8588
rect 45557 8585 45569 8588
rect 45603 8585 45615 8619
rect 45557 8579 45615 8585
rect 45925 8619 45983 8625
rect 45925 8585 45937 8619
rect 45971 8585 45983 8619
rect 45925 8579 45983 8585
rect 6549 8551 6607 8557
rect 6549 8517 6561 8551
rect 6595 8548 6607 8551
rect 11238 8548 11244 8560
rect 6595 8520 7788 8548
rect 6595 8517 6607 8520
rect 6549 8511 6607 8517
rect 5859 8452 6132 8480
rect 6181 8483 6239 8489
rect 5859 8449 5871 8452
rect 5813 8443 5871 8449
rect 6181 8449 6193 8483
rect 6227 8480 6239 8483
rect 6270 8480 6276 8492
rect 6227 8452 6276 8480
rect 6227 8449 6239 8452
rect 6181 8443 6239 8449
rect 5460 8412 5488 8443
rect 6270 8440 6276 8452
rect 6328 8440 6334 8492
rect 6822 8480 6828 8492
rect 6472 8452 6828 8480
rect 6472 8412 6500 8452
rect 6822 8440 6828 8452
rect 6880 8440 6886 8492
rect 6932 8489 6960 8520
rect 6917 8483 6975 8489
rect 6917 8449 6929 8483
rect 6963 8449 6975 8483
rect 6917 8443 6975 8449
rect 7285 8483 7343 8489
rect 7285 8449 7297 8483
rect 7331 8480 7343 8483
rect 7331 8452 7512 8480
rect 7331 8449 7343 8452
rect 7285 8443 7343 8449
rect 5460 8384 6500 8412
rect 6822 8344 6828 8356
rect 3620 8316 6828 8344
rect 6822 8304 6828 8316
rect 6880 8304 6886 8356
rect 7484 8344 7512 8452
rect 7650 8440 7656 8492
rect 7708 8440 7714 8492
rect 7760 8412 7788 8520
rect 10612 8520 11244 8548
rect 7834 8440 7840 8492
rect 7892 8480 7898 8492
rect 8021 8483 8079 8489
rect 8021 8480 8033 8483
rect 7892 8452 8033 8480
rect 7892 8440 7898 8452
rect 8021 8449 8033 8452
rect 8067 8449 8079 8483
rect 8021 8443 8079 8449
rect 8386 8440 8392 8492
rect 8444 8440 8450 8492
rect 8754 8440 8760 8492
rect 8812 8440 8818 8492
rect 9490 8440 9496 8492
rect 9548 8440 9554 8492
rect 9858 8440 9864 8492
rect 9916 8440 9922 8492
rect 10226 8440 10232 8492
rect 10284 8440 10290 8492
rect 10612 8489 10640 8520
rect 11238 8508 11244 8520
rect 11296 8508 11302 8560
rect 11422 8508 11428 8560
rect 11480 8548 11486 8560
rect 11480 8520 13308 8548
rect 11480 8508 11486 8520
rect 10597 8483 10655 8489
rect 10597 8449 10609 8483
rect 10643 8449 10655 8483
rect 10597 8443 10655 8449
rect 10962 8440 10968 8492
rect 11020 8440 11026 8492
rect 11333 8483 11391 8489
rect 11333 8449 11345 8483
rect 11379 8449 11391 8483
rect 11333 8443 11391 8449
rect 12069 8483 12127 8489
rect 12069 8449 12081 8483
rect 12115 8449 12127 8483
rect 12069 8443 12127 8449
rect 12437 8483 12495 8489
rect 12437 8449 12449 8483
rect 12483 8480 12495 8483
rect 12710 8480 12716 8492
rect 12483 8452 12716 8480
rect 12483 8449 12495 8452
rect 12437 8443 12495 8449
rect 7760 8384 11284 8412
rect 11146 8344 11152 8356
rect 7484 8316 11152 8344
rect 11146 8304 11152 8316
rect 11204 8304 11210 8356
rect 7006 8276 7012 8288
rect 1964 8248 7012 8276
rect 7006 8236 7012 8248
rect 7064 8236 7070 8288
rect 11256 8276 11284 8384
rect 11348 8344 11376 8443
rect 12084 8412 12112 8443
rect 12710 8440 12716 8452
rect 12768 8440 12774 8492
rect 12805 8483 12863 8489
rect 12805 8449 12817 8483
rect 12851 8449 12863 8483
rect 12805 8443 12863 8449
rect 12618 8412 12624 8424
rect 12084 8384 12624 8412
rect 12618 8372 12624 8384
rect 12676 8372 12682 8424
rect 12820 8412 12848 8443
rect 13170 8440 13176 8492
rect 13228 8440 13234 8492
rect 13280 8489 13308 8520
rect 14642 8508 14648 8560
rect 14700 8548 14706 8560
rect 19426 8548 19432 8560
rect 14700 8520 18092 8548
rect 14700 8508 14706 8520
rect 13265 8483 13323 8489
rect 13265 8449 13277 8483
rect 13311 8449 13323 8483
rect 13265 8443 13323 8449
rect 13630 8440 13636 8492
rect 13688 8440 13694 8492
rect 13722 8440 13728 8492
rect 13780 8480 13786 8492
rect 14369 8483 14427 8489
rect 14369 8480 14381 8483
rect 13780 8452 14381 8480
rect 13780 8440 13786 8452
rect 14369 8449 14381 8452
rect 14415 8449 14427 8483
rect 14369 8443 14427 8449
rect 14458 8440 14464 8492
rect 14516 8480 14522 8492
rect 14737 8483 14795 8489
rect 14737 8480 14749 8483
rect 14516 8452 14749 8480
rect 14516 8440 14522 8452
rect 14737 8449 14749 8452
rect 14783 8449 14795 8483
rect 14737 8443 14795 8449
rect 15102 8440 15108 8492
rect 15160 8440 15166 8492
rect 15470 8440 15476 8492
rect 15528 8440 15534 8492
rect 15838 8440 15844 8492
rect 15896 8440 15902 8492
rect 16206 8440 16212 8492
rect 16264 8440 16270 8492
rect 16942 8440 16948 8492
rect 17000 8440 17006 8492
rect 17586 8440 17592 8492
rect 17644 8440 17650 8492
rect 17954 8440 17960 8492
rect 18012 8440 18018 8492
rect 18064 8480 18092 8520
rect 18340 8520 19432 8548
rect 18138 8480 18144 8492
rect 18064 8452 18144 8480
rect 18138 8440 18144 8452
rect 18196 8440 18202 8492
rect 18340 8489 18368 8520
rect 19426 8508 19432 8520
rect 19484 8508 19490 8560
rect 18325 8483 18383 8489
rect 18325 8449 18337 8483
rect 18371 8449 18383 8483
rect 18325 8443 18383 8449
rect 18693 8483 18751 8489
rect 18693 8449 18705 8483
rect 18739 8480 18751 8483
rect 19073 8483 19131 8489
rect 18739 8452 19012 8480
rect 18739 8449 18751 8452
rect 18693 8443 18751 8449
rect 16482 8412 16488 8424
rect 12820 8384 16488 8412
rect 16482 8372 16488 8384
rect 16540 8372 16546 8424
rect 17770 8412 17776 8424
rect 17420 8384 17776 8412
rect 12434 8344 12440 8356
rect 11348 8316 12440 8344
rect 12434 8304 12440 8316
rect 12492 8304 12498 8356
rect 17420 8353 17448 8384
rect 17770 8372 17776 8384
rect 17828 8372 17834 8424
rect 17405 8347 17463 8353
rect 12544 8316 17356 8344
rect 12544 8276 12572 8316
rect 11256 8248 12572 8276
rect 17328 8276 17356 8316
rect 17405 8313 17417 8347
rect 17451 8313 17463 8347
rect 18046 8344 18052 8356
rect 17405 8307 17463 8313
rect 17512 8316 18052 8344
rect 17512 8276 17540 8316
rect 18046 8304 18052 8316
rect 18104 8304 18110 8356
rect 18509 8347 18567 8353
rect 18509 8313 18521 8347
rect 18555 8344 18567 8347
rect 18874 8344 18880 8356
rect 18555 8316 18880 8344
rect 18555 8313 18567 8316
rect 18509 8307 18567 8313
rect 18874 8304 18880 8316
rect 18932 8304 18938 8356
rect 18984 8344 19012 8452
rect 19073 8449 19085 8483
rect 19119 8480 19131 8483
rect 19720 8480 19748 8576
rect 29086 8508 29092 8560
rect 29144 8548 29150 8560
rect 29144 8520 41092 8548
rect 29144 8508 29150 8520
rect 19119 8452 19748 8480
rect 19797 8483 19855 8489
rect 19119 8449 19131 8452
rect 19073 8443 19131 8449
rect 19797 8449 19809 8483
rect 19843 8449 19855 8483
rect 19797 8443 19855 8449
rect 19981 8483 20039 8489
rect 19981 8449 19993 8483
rect 20027 8480 20039 8483
rect 20349 8483 20407 8489
rect 20349 8480 20361 8483
rect 20027 8452 20361 8480
rect 20027 8449 20039 8452
rect 19981 8443 20039 8449
rect 20349 8449 20361 8452
rect 20395 8449 20407 8483
rect 20349 8443 20407 8449
rect 20717 8483 20775 8489
rect 20717 8449 20729 8483
rect 20763 8480 20775 8483
rect 20901 8483 20959 8489
rect 20901 8480 20913 8483
rect 20763 8452 20913 8480
rect 20763 8449 20775 8452
rect 20717 8443 20775 8449
rect 20901 8449 20913 8452
rect 20947 8480 20959 8483
rect 37182 8480 37188 8492
rect 20947 8452 37188 8480
rect 20947 8449 20959 8452
rect 20901 8443 20959 8449
rect 19812 8412 19840 8443
rect 37182 8440 37188 8452
rect 37240 8440 37246 8492
rect 38746 8440 38752 8492
rect 38804 8480 38810 8492
rect 40129 8483 40187 8489
rect 40129 8480 40141 8483
rect 38804 8452 40141 8480
rect 38804 8440 38810 8452
rect 40129 8449 40141 8452
rect 40175 8449 40187 8483
rect 40129 8443 40187 8449
rect 40313 8483 40371 8489
rect 40313 8449 40325 8483
rect 40359 8449 40371 8483
rect 40313 8443 40371 8449
rect 30742 8412 30748 8424
rect 19812 8384 30748 8412
rect 30742 8372 30748 8384
rect 30800 8372 30806 8424
rect 35802 8372 35808 8424
rect 35860 8412 35866 8424
rect 35860 8384 38700 8412
rect 35860 8372 35866 8384
rect 19702 8344 19708 8356
rect 18984 8316 19708 8344
rect 19702 8304 19708 8316
rect 19760 8304 19766 8356
rect 19981 8347 20039 8353
rect 19981 8313 19993 8347
rect 20027 8344 20039 8347
rect 38562 8344 38568 8356
rect 20027 8316 38568 8344
rect 20027 8313 20039 8316
rect 19981 8307 20039 8313
rect 38562 8304 38568 8316
rect 38620 8304 38626 8356
rect 38672 8344 38700 8384
rect 39666 8372 39672 8424
rect 39724 8412 39730 8424
rect 40328 8412 40356 8443
rect 40678 8440 40684 8492
rect 40736 8440 40742 8492
rect 41064 8489 41092 8520
rect 41156 8520 44312 8548
rect 41049 8483 41107 8489
rect 41049 8449 41061 8483
rect 41095 8449 41107 8483
rect 41049 8443 41107 8449
rect 39724 8384 40356 8412
rect 39724 8372 39730 8384
rect 41156 8344 41184 8520
rect 41414 8440 41420 8492
rect 41472 8440 41478 8492
rect 41782 8440 41788 8492
rect 41840 8440 41846 8492
rect 41874 8440 41880 8492
rect 41932 8480 41938 8492
rect 42429 8483 42487 8489
rect 42429 8480 42441 8483
rect 41932 8452 42441 8480
rect 41932 8440 41938 8452
rect 42429 8449 42441 8452
rect 42475 8449 42487 8483
rect 42429 8443 42487 8449
rect 42797 8483 42855 8489
rect 42797 8449 42809 8483
rect 42843 8480 42855 8483
rect 42978 8480 42984 8492
rect 42843 8452 42984 8480
rect 42843 8449 42855 8452
rect 42797 8443 42855 8449
rect 42978 8440 42984 8452
rect 43036 8440 43042 8492
rect 43165 8483 43223 8489
rect 43165 8449 43177 8483
rect 43211 8449 43223 8483
rect 43165 8443 43223 8449
rect 42242 8372 42248 8424
rect 42300 8412 42306 8424
rect 43180 8412 43208 8443
rect 43346 8440 43352 8492
rect 43404 8480 43410 8492
rect 43533 8483 43591 8489
rect 43533 8480 43545 8483
rect 43404 8452 43545 8480
rect 43404 8440 43410 8452
rect 43533 8449 43545 8452
rect 43579 8449 43591 8483
rect 43533 8443 43591 8449
rect 43714 8440 43720 8492
rect 43772 8480 43778 8492
rect 43901 8483 43959 8489
rect 43901 8480 43913 8483
rect 43772 8452 43913 8480
rect 43772 8440 43778 8452
rect 43901 8449 43913 8452
rect 43947 8449 43959 8483
rect 43901 8443 43959 8449
rect 43990 8440 43996 8492
rect 44048 8480 44054 8492
rect 44284 8489 44312 8520
rect 44910 8508 44916 8560
rect 44968 8548 44974 8560
rect 45940 8548 45968 8579
rect 46014 8576 46020 8628
rect 46072 8616 46078 8628
rect 46661 8619 46719 8625
rect 46661 8616 46673 8619
rect 46072 8588 46673 8616
rect 46072 8576 46078 8588
rect 46661 8585 46673 8588
rect 46707 8585 46719 8619
rect 46661 8579 46719 8585
rect 44968 8520 45968 8548
rect 46032 8520 46520 8548
rect 44968 8508 44974 8520
rect 46032 8492 46060 8520
rect 44269 8483 44327 8489
rect 44048 8452 44220 8480
rect 44048 8440 44054 8452
rect 42300 8384 43208 8412
rect 42300 8372 42306 8384
rect 43622 8372 43628 8424
rect 43680 8412 43686 8424
rect 44192 8412 44220 8452
rect 44269 8449 44281 8483
rect 44315 8449 44327 8483
rect 44269 8443 44327 8449
rect 44358 8440 44364 8492
rect 44416 8480 44422 8492
rect 45005 8483 45063 8489
rect 45005 8480 45017 8483
rect 44416 8452 45017 8480
rect 44416 8440 44422 8452
rect 45005 8449 45017 8452
rect 45051 8449 45063 8483
rect 45005 8443 45063 8449
rect 45373 8483 45431 8489
rect 45373 8449 45385 8483
rect 45419 8480 45431 8483
rect 45462 8480 45468 8492
rect 45419 8452 45468 8480
rect 45419 8449 45431 8452
rect 45373 8443 45431 8449
rect 45462 8440 45468 8452
rect 45520 8440 45526 8492
rect 45741 8483 45799 8489
rect 45741 8449 45753 8483
rect 45787 8449 45799 8483
rect 45741 8443 45799 8449
rect 45756 8412 45784 8443
rect 46014 8440 46020 8492
rect 46072 8440 46078 8492
rect 46492 8489 46520 8520
rect 46109 8483 46167 8489
rect 46109 8449 46121 8483
rect 46155 8449 46167 8483
rect 46109 8443 46167 8449
rect 46477 8483 46535 8489
rect 46477 8449 46489 8483
rect 46523 8449 46535 8483
rect 46477 8443 46535 8449
rect 46124 8412 46152 8443
rect 46566 8440 46572 8492
rect 46624 8480 46630 8492
rect 46845 8483 46903 8489
rect 46845 8480 46857 8483
rect 46624 8452 46857 8480
rect 46624 8440 46630 8452
rect 46845 8449 46857 8452
rect 46891 8449 46903 8483
rect 46845 8443 46903 8449
rect 43680 8384 44128 8412
rect 44192 8384 45784 8412
rect 45848 8384 46152 8412
rect 43680 8372 43686 8384
rect 38672 8316 41184 8344
rect 42426 8304 42432 8356
rect 42484 8344 42490 8356
rect 42981 8347 43039 8353
rect 42981 8344 42993 8347
rect 42484 8316 42993 8344
rect 42484 8304 42490 8316
rect 42981 8313 42993 8316
rect 43027 8313 43039 8347
rect 42981 8307 43039 8313
rect 43162 8304 43168 8356
rect 43220 8344 43226 8356
rect 44100 8353 44128 8384
rect 43717 8347 43775 8353
rect 43717 8344 43729 8347
rect 43220 8316 43729 8344
rect 43220 8304 43226 8316
rect 43717 8313 43729 8316
rect 43763 8313 43775 8347
rect 43717 8307 43775 8313
rect 44085 8347 44143 8353
rect 44085 8313 44097 8347
rect 44131 8313 44143 8347
rect 44085 8307 44143 8313
rect 44266 8304 44272 8356
rect 44324 8344 44330 8356
rect 45189 8347 45247 8353
rect 45189 8344 45201 8347
rect 44324 8316 45201 8344
rect 44324 8304 44330 8316
rect 45189 8313 45201 8316
rect 45235 8313 45247 8347
rect 45189 8307 45247 8313
rect 45462 8304 45468 8356
rect 45520 8344 45526 8356
rect 45848 8344 45876 8384
rect 46198 8372 46204 8424
rect 46256 8412 46262 8424
rect 46256 8384 47072 8412
rect 46256 8372 46262 8384
rect 45520 8316 45876 8344
rect 46293 8347 46351 8353
rect 45520 8304 45526 8316
rect 46293 8313 46305 8347
rect 46339 8344 46351 8347
rect 46382 8344 46388 8356
rect 46339 8316 46388 8344
rect 46339 8313 46351 8316
rect 46293 8307 46351 8313
rect 46382 8304 46388 8316
rect 46440 8304 46446 8356
rect 47044 8353 47072 8384
rect 47029 8347 47087 8353
rect 47029 8313 47041 8347
rect 47075 8313 47087 8347
rect 47029 8307 47087 8313
rect 17328 8248 17540 8276
rect 39942 8236 39948 8288
rect 40000 8276 40006 8288
rect 46014 8276 46020 8288
rect 40000 8248 46020 8276
rect 40000 8236 40006 8248
rect 46014 8236 46020 8248
rect 46072 8236 46078 8288
rect 1104 8186 47840 8208
rect 1104 8134 1950 8186
rect 2002 8134 2014 8186
rect 2066 8134 2078 8186
rect 2130 8134 2142 8186
rect 2194 8134 2206 8186
rect 2258 8134 7950 8186
rect 8002 8134 8014 8186
rect 8066 8134 8078 8186
rect 8130 8134 8142 8186
rect 8194 8134 8206 8186
rect 8258 8134 13950 8186
rect 14002 8134 14014 8186
rect 14066 8134 14078 8186
rect 14130 8134 14142 8186
rect 14194 8134 14206 8186
rect 14258 8134 19950 8186
rect 20002 8134 20014 8186
rect 20066 8134 20078 8186
rect 20130 8134 20142 8186
rect 20194 8134 20206 8186
rect 20258 8134 25950 8186
rect 26002 8134 26014 8186
rect 26066 8134 26078 8186
rect 26130 8134 26142 8186
rect 26194 8134 26206 8186
rect 26258 8134 31950 8186
rect 32002 8134 32014 8186
rect 32066 8134 32078 8186
rect 32130 8134 32142 8186
rect 32194 8134 32206 8186
rect 32258 8134 37950 8186
rect 38002 8134 38014 8186
rect 38066 8134 38078 8186
rect 38130 8134 38142 8186
rect 38194 8134 38206 8186
rect 38258 8134 43950 8186
rect 44002 8134 44014 8186
rect 44066 8134 44078 8186
rect 44130 8134 44142 8186
rect 44194 8134 44206 8186
rect 44258 8134 47840 8186
rect 1104 8112 47840 8134
rect 1578 8032 1584 8084
rect 1636 8032 1642 8084
rect 3786 8032 3792 8084
rect 3844 8072 3850 8084
rect 3973 8075 4031 8081
rect 3973 8072 3985 8075
rect 3844 8044 3985 8072
rect 3844 8032 3850 8044
rect 3973 8041 3985 8044
rect 4019 8041 4031 8075
rect 3973 8035 4031 8041
rect 6362 8032 6368 8084
rect 6420 8072 6426 8084
rect 6549 8075 6607 8081
rect 6549 8072 6561 8075
rect 6420 8044 6561 8072
rect 6420 8032 6426 8044
rect 6549 8041 6561 8044
rect 6595 8041 6607 8075
rect 6549 8035 6607 8041
rect 8846 8032 8852 8084
rect 8904 8072 8910 8084
rect 9125 8075 9183 8081
rect 9125 8072 9137 8075
rect 8904 8044 9137 8072
rect 8904 8032 8910 8044
rect 9125 8041 9137 8044
rect 9171 8041 9183 8075
rect 9125 8035 9183 8041
rect 10781 8075 10839 8081
rect 10781 8041 10793 8075
rect 10827 8072 10839 8075
rect 10870 8072 10876 8084
rect 10827 8044 10876 8072
rect 10827 8041 10839 8044
rect 10781 8035 10839 8041
rect 10870 8032 10876 8044
rect 10928 8032 10934 8084
rect 11333 8075 11391 8081
rect 11333 8041 11345 8075
rect 11379 8072 11391 8075
rect 11422 8072 11428 8084
rect 11379 8044 11428 8072
rect 11379 8041 11391 8044
rect 11333 8035 11391 8041
rect 11422 8032 11428 8044
rect 11480 8032 11486 8084
rect 11514 8032 11520 8084
rect 11572 8072 11578 8084
rect 12345 8075 12403 8081
rect 12345 8072 12357 8075
rect 11572 8044 12357 8072
rect 11572 8032 11578 8044
rect 12345 8041 12357 8044
rect 12391 8041 12403 8075
rect 12345 8035 12403 8041
rect 12434 8032 12440 8084
rect 12492 8072 12498 8084
rect 12986 8072 12992 8084
rect 12492 8044 12992 8072
rect 12492 8032 12498 8044
rect 12986 8032 12992 8044
rect 13044 8032 13050 8084
rect 13081 8075 13139 8081
rect 13081 8041 13093 8075
rect 13127 8072 13139 8075
rect 13722 8072 13728 8084
rect 13127 8044 13728 8072
rect 13127 8041 13139 8044
rect 13081 8035 13139 8041
rect 13722 8032 13728 8044
rect 13780 8032 13786 8084
rect 14274 8032 14280 8084
rect 14332 8072 14338 8084
rect 14369 8075 14427 8081
rect 14369 8072 14381 8075
rect 14332 8044 14381 8072
rect 14332 8032 14338 8044
rect 14369 8041 14381 8044
rect 14415 8041 14427 8075
rect 14369 8035 14427 8041
rect 14737 8075 14795 8081
rect 14737 8041 14749 8075
rect 14783 8072 14795 8075
rect 15102 8072 15108 8084
rect 14783 8044 15108 8072
rect 14783 8041 14795 8044
rect 14737 8035 14795 8041
rect 15102 8032 15108 8044
rect 15160 8032 15166 8084
rect 16666 8032 16672 8084
rect 16724 8072 16730 8084
rect 16945 8075 17003 8081
rect 16945 8072 16957 8075
rect 16724 8044 16957 8072
rect 16724 8032 16730 8044
rect 16945 8041 16957 8044
rect 16991 8041 17003 8075
rect 16945 8035 17003 8041
rect 17034 8032 17040 8084
rect 17092 8072 17098 8084
rect 17313 8075 17371 8081
rect 17313 8072 17325 8075
rect 17092 8044 17325 8072
rect 17092 8032 17098 8044
rect 17313 8041 17325 8044
rect 17359 8041 17371 8075
rect 17313 8035 17371 8041
rect 17586 8032 17592 8084
rect 17644 8072 17650 8084
rect 17773 8075 17831 8081
rect 17773 8072 17785 8075
rect 17644 8044 17785 8072
rect 17644 8032 17650 8044
rect 17773 8041 17785 8044
rect 17819 8041 17831 8075
rect 17773 8035 17831 8041
rect 17954 8032 17960 8084
rect 18012 8072 18018 8084
rect 18141 8075 18199 8081
rect 18141 8072 18153 8075
rect 18012 8044 18153 8072
rect 18012 8032 18018 8044
rect 18141 8041 18153 8044
rect 18187 8041 18199 8075
rect 18141 8035 18199 8041
rect 19426 8032 19432 8084
rect 19484 8032 19490 8084
rect 19702 8032 19708 8084
rect 19760 8072 19766 8084
rect 20165 8075 20223 8081
rect 20165 8072 20177 8075
rect 19760 8044 20177 8072
rect 19760 8032 19766 8044
rect 20165 8041 20177 8044
rect 20211 8041 20223 8075
rect 20165 8035 20223 8041
rect 21358 8032 21364 8084
rect 21416 8072 21422 8084
rect 22646 8072 22652 8084
rect 21416 8044 22652 8072
rect 21416 8032 21422 8044
rect 22646 8032 22652 8044
rect 22704 8032 22710 8084
rect 24118 8032 24124 8084
rect 24176 8072 24182 8084
rect 29825 8075 29883 8081
rect 29825 8072 29837 8075
rect 24176 8044 29837 8072
rect 24176 8032 24182 8044
rect 29825 8041 29837 8044
rect 29871 8041 29883 8075
rect 29825 8035 29883 8041
rect 30190 8032 30196 8084
rect 30248 8032 30254 8084
rect 35066 8032 35072 8084
rect 35124 8072 35130 8084
rect 35124 8044 40172 8072
rect 35124 8032 35130 8044
rect 5350 7964 5356 8016
rect 5408 7964 5414 8016
rect 11057 8007 11115 8013
rect 11057 7973 11069 8007
rect 11103 8004 11115 8007
rect 13630 8004 13636 8016
rect 11103 7976 13636 8004
rect 11103 7973 11115 7976
rect 11057 7967 11115 7973
rect 13630 7964 13636 7976
rect 13688 7964 13694 8016
rect 13909 8007 13967 8013
rect 13909 7973 13921 8007
rect 13955 8004 13967 8007
rect 14458 8004 14464 8016
rect 13955 7976 14464 8004
rect 13955 7973 13967 7976
rect 13909 7967 13967 7973
rect 14458 7964 14464 7976
rect 14516 7964 14522 8016
rect 18046 7964 18052 8016
rect 18104 8004 18110 8016
rect 27065 8007 27123 8013
rect 27065 8004 27077 8007
rect 18104 7976 25820 8004
rect 18104 7964 18110 7976
rect 12434 7936 12440 7948
rect 1780 7908 12440 7936
rect 1780 7877 1808 7908
rect 12434 7896 12440 7908
rect 12492 7896 12498 7948
rect 13170 7896 13176 7948
rect 13228 7936 13234 7948
rect 16298 7936 16304 7948
rect 13228 7908 16304 7936
rect 13228 7896 13234 7908
rect 16298 7896 16304 7908
rect 16356 7896 16362 7948
rect 18509 7939 18567 7945
rect 18509 7905 18521 7939
rect 18555 7936 18567 7939
rect 18555 7908 18736 7936
rect 18555 7905 18567 7908
rect 18509 7899 18567 7905
rect 1765 7871 1823 7877
rect 1765 7837 1777 7871
rect 1811 7837 1823 7871
rect 1765 7831 1823 7837
rect 2406 7828 2412 7880
rect 2464 7828 2470 7880
rect 4154 7828 4160 7880
rect 4212 7828 4218 7880
rect 5166 7828 5172 7880
rect 5224 7828 5230 7880
rect 6730 7828 6736 7880
rect 6788 7828 6794 7880
rect 9309 7871 9367 7877
rect 9309 7837 9321 7871
rect 9355 7868 9367 7871
rect 9582 7868 9588 7880
rect 9355 7840 9588 7868
rect 9355 7837 9367 7840
rect 9309 7831 9367 7837
rect 9582 7828 9588 7840
rect 9640 7828 9646 7880
rect 10781 7871 10839 7877
rect 10781 7837 10793 7871
rect 10827 7868 10839 7871
rect 10873 7871 10931 7877
rect 10873 7868 10885 7871
rect 10827 7840 10885 7868
rect 10827 7837 10839 7840
rect 10781 7831 10839 7837
rect 10873 7837 10885 7840
rect 10919 7837 10931 7871
rect 10873 7831 10931 7837
rect 11149 7871 11207 7877
rect 11149 7837 11161 7871
rect 11195 7868 11207 7871
rect 11790 7868 11796 7880
rect 11195 7840 11796 7868
rect 11195 7837 11207 7840
rect 11149 7831 11207 7837
rect 11790 7828 11796 7840
rect 11848 7828 11854 7880
rect 11885 7871 11943 7877
rect 11885 7837 11897 7871
rect 11931 7868 11943 7871
rect 11974 7868 11980 7880
rect 11931 7840 11980 7868
rect 11931 7837 11943 7840
rect 11885 7831 11943 7837
rect 11974 7828 11980 7840
rect 12032 7828 12038 7880
rect 12526 7877 12532 7880
rect 12522 7831 12532 7877
rect 12526 7828 12532 7831
rect 12584 7828 12590 7880
rect 12805 7871 12863 7877
rect 12805 7837 12817 7871
rect 12851 7868 12863 7871
rect 12897 7871 12955 7877
rect 12897 7868 12909 7871
rect 12851 7840 12909 7868
rect 12851 7837 12863 7840
rect 12805 7831 12863 7837
rect 12897 7837 12909 7840
rect 12943 7837 12955 7871
rect 12897 7831 12955 7837
rect 13538 7828 13544 7880
rect 13596 7868 13602 7880
rect 13725 7871 13783 7877
rect 13725 7868 13737 7871
rect 13596 7840 13737 7868
rect 13596 7828 13602 7840
rect 13725 7837 13737 7840
rect 13771 7837 13783 7871
rect 13725 7831 13783 7837
rect 14185 7871 14243 7877
rect 14185 7837 14197 7871
rect 14231 7837 14243 7871
rect 14185 7831 14243 7837
rect 198 7760 204 7812
rect 256 7800 262 7812
rect 2225 7803 2283 7809
rect 2225 7800 2237 7803
rect 256 7772 2237 7800
rect 256 7760 262 7772
rect 2225 7769 2237 7772
rect 2271 7769 2283 7803
rect 14200 7800 14228 7831
rect 14550 7828 14556 7880
rect 14608 7828 14614 7880
rect 16758 7828 16764 7880
rect 16816 7828 16822 7880
rect 17126 7828 17132 7880
rect 17184 7828 17190 7880
rect 17957 7871 18015 7877
rect 17957 7837 17969 7871
rect 18003 7868 18015 7871
rect 18230 7868 18236 7880
rect 18003 7840 18236 7868
rect 18003 7837 18015 7840
rect 17957 7831 18015 7837
rect 18230 7828 18236 7840
rect 18288 7828 18294 7880
rect 18322 7828 18328 7880
rect 18380 7828 18386 7880
rect 18708 7877 18736 7908
rect 18874 7896 18880 7948
rect 18932 7936 18938 7948
rect 24118 7936 24124 7948
rect 18932 7908 24124 7936
rect 18932 7896 18938 7908
rect 24118 7896 24124 7908
rect 24176 7896 24182 7948
rect 25792 7936 25820 7976
rect 25976 7976 27077 8004
rect 25976 7936 26004 7976
rect 27065 7973 27077 7976
rect 27111 7973 27123 8007
rect 34241 8007 34299 8013
rect 34241 8004 34253 8007
rect 27065 7967 27123 7973
rect 27172 7976 34253 8004
rect 27172 7936 27200 7976
rect 34241 7973 34253 7976
rect 34287 7973 34299 8007
rect 34241 7967 34299 7973
rect 37001 8007 37059 8013
rect 37001 7973 37013 8007
rect 37047 8004 37059 8007
rect 39942 8004 39948 8016
rect 37047 7976 39948 8004
rect 37047 7973 37059 7976
rect 37001 7967 37059 7973
rect 39942 7964 39948 7976
rect 40000 7964 40006 8016
rect 40144 8004 40172 8044
rect 40494 8032 40500 8084
rect 40552 8032 40558 8084
rect 41598 8032 41604 8084
rect 41656 8032 41662 8084
rect 44818 8032 44824 8084
rect 44876 8072 44882 8084
rect 45281 8075 45339 8081
rect 45281 8072 45293 8075
rect 44876 8044 45293 8072
rect 44876 8032 44882 8044
rect 45281 8041 45293 8044
rect 45327 8041 45339 8075
rect 45281 8035 45339 8041
rect 45646 8032 45652 8084
rect 45704 8032 45710 8084
rect 46474 8032 46480 8084
rect 46532 8072 46538 8084
rect 46753 8075 46811 8081
rect 46753 8072 46765 8075
rect 46532 8044 46765 8072
rect 46532 8032 46538 8044
rect 46753 8041 46765 8044
rect 46799 8041 46811 8075
rect 46753 8035 46811 8041
rect 46842 8032 46848 8084
rect 46900 8072 46906 8084
rect 47121 8075 47179 8081
rect 47121 8072 47133 8075
rect 46900 8044 47133 8072
rect 46900 8032 46906 8044
rect 47121 8041 47133 8044
rect 47167 8041 47179 8075
rect 47121 8035 47179 8041
rect 40144 7976 40724 8004
rect 25792 7908 26004 7936
rect 26068 7908 27200 7936
rect 18693 7871 18751 7877
rect 18693 7837 18705 7871
rect 18739 7837 18751 7871
rect 18693 7831 18751 7837
rect 19337 7871 19395 7877
rect 19337 7837 19349 7871
rect 19383 7868 19395 7871
rect 19613 7871 19671 7877
rect 19613 7868 19625 7871
rect 19383 7840 19625 7868
rect 19383 7837 19395 7840
rect 19337 7831 19395 7837
rect 19613 7837 19625 7840
rect 19659 7868 19671 7871
rect 19794 7868 19800 7880
rect 19659 7840 19800 7868
rect 19659 7837 19671 7840
rect 19613 7831 19671 7837
rect 19794 7828 19800 7840
rect 19852 7828 19858 7880
rect 20073 7871 20131 7877
rect 20073 7837 20085 7871
rect 20119 7868 20131 7871
rect 20349 7871 20407 7877
rect 20349 7868 20361 7871
rect 20119 7840 20361 7868
rect 20119 7837 20131 7840
rect 20073 7831 20131 7837
rect 20349 7837 20361 7840
rect 20395 7868 20407 7871
rect 20438 7868 20444 7880
rect 20395 7840 20444 7868
rect 20395 7837 20407 7840
rect 20349 7831 20407 7837
rect 20438 7828 20444 7840
rect 20496 7828 20502 7880
rect 20530 7828 20536 7880
rect 20588 7868 20594 7880
rect 21545 7871 21603 7877
rect 21545 7868 21557 7871
rect 20588 7840 21557 7868
rect 20588 7828 20594 7840
rect 21545 7837 21557 7840
rect 21591 7837 21603 7871
rect 21545 7831 21603 7837
rect 21634 7828 21640 7880
rect 21692 7868 21698 7880
rect 26068 7868 26096 7908
rect 27706 7896 27712 7948
rect 27764 7936 27770 7948
rect 27764 7908 28580 7936
rect 27764 7896 27770 7908
rect 21692 7840 26096 7868
rect 26237 7871 26295 7877
rect 21692 7828 21698 7840
rect 26237 7837 26249 7871
rect 26283 7868 26295 7871
rect 26602 7868 26608 7880
rect 26283 7840 26608 7868
rect 26283 7837 26295 7840
rect 26237 7831 26295 7837
rect 26602 7828 26608 7840
rect 26660 7828 26666 7880
rect 26878 7828 26884 7880
rect 26936 7868 26942 7880
rect 27249 7871 27307 7877
rect 27249 7868 27261 7871
rect 26936 7840 27261 7868
rect 26936 7828 26942 7840
rect 27249 7837 27261 7840
rect 27295 7837 27307 7871
rect 27249 7831 27307 7837
rect 27338 7828 27344 7880
rect 27396 7868 27402 7880
rect 28445 7871 28503 7877
rect 28445 7868 28457 7871
rect 27396 7840 28457 7868
rect 27396 7828 27402 7840
rect 28445 7837 28457 7840
rect 28491 7837 28503 7871
rect 28552 7868 28580 7908
rect 29546 7896 29552 7948
rect 29604 7936 29610 7948
rect 29604 7908 30880 7936
rect 29604 7896 29610 7908
rect 29733 7871 29791 7877
rect 29733 7868 29745 7871
rect 28552 7840 29745 7868
rect 28445 7831 28503 7837
rect 29733 7837 29745 7840
rect 29779 7837 29791 7871
rect 29733 7831 29791 7837
rect 29914 7828 29920 7880
rect 29972 7868 29978 7880
rect 30852 7877 30880 7908
rect 34698 7896 34704 7948
rect 34756 7936 34762 7948
rect 34756 7908 38424 7936
rect 34756 7896 34762 7908
rect 30009 7871 30067 7877
rect 30009 7868 30021 7871
rect 29972 7840 30021 7868
rect 29972 7828 29978 7840
rect 30009 7837 30021 7840
rect 30055 7837 30067 7871
rect 30009 7831 30067 7837
rect 30285 7871 30343 7877
rect 30285 7837 30297 7871
rect 30331 7868 30343 7871
rect 30377 7871 30435 7877
rect 30377 7868 30389 7871
rect 30331 7840 30389 7868
rect 30331 7837 30343 7840
rect 30285 7831 30343 7837
rect 30377 7837 30389 7840
rect 30423 7837 30435 7871
rect 30377 7831 30435 7837
rect 30837 7871 30895 7877
rect 30837 7837 30849 7871
rect 30883 7837 30895 7871
rect 30837 7831 30895 7837
rect 32490 7828 32496 7880
rect 32548 7868 32554 7880
rect 34425 7871 34483 7877
rect 34425 7868 34437 7871
rect 32548 7840 34437 7868
rect 32548 7828 32554 7840
rect 34425 7837 34437 7840
rect 34471 7837 34483 7871
rect 34425 7831 34483 7837
rect 36817 7871 36875 7877
rect 36817 7837 36829 7871
rect 36863 7868 36875 7871
rect 38286 7868 38292 7880
rect 36863 7840 38292 7868
rect 36863 7837 36875 7840
rect 36817 7831 36875 7837
rect 38286 7828 38292 7840
rect 38344 7828 38350 7880
rect 38396 7868 38424 7908
rect 40696 7877 40724 7976
rect 46014 7964 46020 8016
rect 46072 7964 46078 8016
rect 46385 8007 46443 8013
rect 46385 7973 46397 8007
rect 46431 8004 46443 8007
rect 47210 8004 47216 8016
rect 46431 7976 47216 8004
rect 46431 7973 46443 7976
rect 46385 7967 46443 7973
rect 47210 7964 47216 7976
rect 47268 7964 47274 8016
rect 44542 7896 44548 7948
rect 44600 7936 44606 7948
rect 44600 7908 46612 7936
rect 44600 7896 44606 7908
rect 39669 7871 39727 7877
rect 39669 7868 39681 7871
rect 38396 7840 39681 7868
rect 39669 7837 39681 7840
rect 39715 7837 39727 7871
rect 39669 7831 39727 7837
rect 40681 7871 40739 7877
rect 40681 7837 40693 7871
rect 40727 7837 40739 7871
rect 40681 7831 40739 7837
rect 41693 7871 41751 7877
rect 41693 7837 41705 7871
rect 41739 7868 41751 7871
rect 41785 7871 41843 7877
rect 41785 7868 41797 7871
rect 41739 7840 41797 7868
rect 41739 7837 41751 7840
rect 41693 7831 41751 7837
rect 41785 7837 41797 7840
rect 41831 7837 41843 7871
rect 41785 7831 41843 7837
rect 45094 7828 45100 7880
rect 45152 7828 45158 7880
rect 45465 7871 45523 7877
rect 45465 7837 45477 7871
rect 45511 7837 45523 7871
rect 45465 7831 45523 7837
rect 2225 7763 2283 7769
rect 12728 7772 14228 7800
rect 12161 7735 12219 7741
rect 12161 7701 12173 7735
rect 12207 7732 12219 7735
rect 12728 7732 12756 7772
rect 14274 7760 14280 7812
rect 14332 7800 14338 7812
rect 21358 7800 21364 7812
rect 14332 7772 21364 7800
rect 14332 7760 14338 7772
rect 21358 7760 21364 7772
rect 21416 7760 21422 7812
rect 25774 7760 25780 7812
rect 25832 7800 25838 7812
rect 25832 7772 28396 7800
rect 25832 7760 25838 7772
rect 12207 7704 12756 7732
rect 12805 7735 12863 7741
rect 12207 7701 12219 7704
rect 12161 7695 12219 7701
rect 12805 7701 12817 7735
rect 12851 7732 12863 7735
rect 15562 7732 15568 7744
rect 12851 7704 15568 7732
rect 12851 7701 12863 7704
rect 12805 7695 12863 7701
rect 15562 7692 15568 7704
rect 15620 7692 15626 7744
rect 17862 7692 17868 7744
rect 17920 7732 17926 7744
rect 18417 7735 18475 7741
rect 18417 7732 18429 7735
rect 17920 7704 18429 7732
rect 17920 7692 17926 7704
rect 18417 7701 18429 7704
rect 18463 7701 18475 7735
rect 18417 7695 18475 7701
rect 18782 7692 18788 7744
rect 18840 7692 18846 7744
rect 18966 7692 18972 7744
rect 19024 7732 19030 7744
rect 21634 7732 21640 7744
rect 19024 7704 21640 7732
rect 19024 7692 19030 7704
rect 21634 7692 21640 7704
rect 21692 7692 21698 7744
rect 21726 7692 21732 7744
rect 21784 7692 21790 7744
rect 22646 7692 22652 7744
rect 22704 7732 22710 7744
rect 26053 7735 26111 7741
rect 26053 7732 26065 7735
rect 22704 7704 26065 7732
rect 22704 7692 22710 7704
rect 26053 7701 26065 7704
rect 26099 7701 26111 7735
rect 26053 7695 26111 7701
rect 28258 7692 28264 7744
rect 28316 7692 28322 7744
rect 28368 7732 28396 7772
rect 29822 7760 29828 7812
rect 29880 7800 29886 7812
rect 29880 7772 30696 7800
rect 29880 7760 29886 7772
rect 29549 7735 29607 7741
rect 29549 7732 29561 7735
rect 28368 7704 29561 7732
rect 29549 7701 29561 7704
rect 29595 7701 29607 7735
rect 29549 7695 29607 7701
rect 30558 7692 30564 7744
rect 30616 7692 30622 7744
rect 30668 7741 30696 7772
rect 30742 7760 30748 7812
rect 30800 7800 30806 7812
rect 30800 7772 39528 7800
rect 30800 7760 30806 7772
rect 39500 7741 39528 7772
rect 39574 7760 39580 7812
rect 39632 7800 39638 7812
rect 45480 7800 45508 7831
rect 45830 7828 45836 7880
rect 45888 7828 45894 7880
rect 46198 7828 46204 7880
rect 46256 7828 46262 7880
rect 46584 7877 46612 7908
rect 46569 7871 46627 7877
rect 46569 7837 46581 7871
rect 46615 7837 46627 7871
rect 46569 7831 46627 7837
rect 46658 7828 46664 7880
rect 46716 7868 46722 7880
rect 46937 7871 46995 7877
rect 46937 7868 46949 7871
rect 46716 7840 46949 7868
rect 46716 7828 46722 7840
rect 46937 7837 46949 7840
rect 46983 7837 46995 7871
rect 46937 7831 46995 7837
rect 39632 7772 45508 7800
rect 39632 7760 39638 7772
rect 30653 7735 30711 7741
rect 30653 7701 30665 7735
rect 30699 7701 30711 7735
rect 30653 7695 30711 7701
rect 39485 7735 39543 7741
rect 39485 7701 39497 7735
rect 39531 7701 39543 7735
rect 39485 7695 39543 7701
rect 41969 7735 42027 7741
rect 41969 7701 41981 7735
rect 42015 7732 42027 7735
rect 43714 7732 43720 7744
rect 42015 7704 43720 7732
rect 42015 7701 42027 7704
rect 41969 7695 42027 7701
rect 43714 7692 43720 7704
rect 43772 7692 43778 7744
rect 1104 7642 47840 7664
rect 1104 7590 3010 7642
rect 3062 7590 3074 7642
rect 3126 7590 3138 7642
rect 3190 7590 3202 7642
rect 3254 7590 3266 7642
rect 3318 7590 9010 7642
rect 9062 7590 9074 7642
rect 9126 7590 9138 7642
rect 9190 7590 9202 7642
rect 9254 7590 9266 7642
rect 9318 7590 15010 7642
rect 15062 7590 15074 7642
rect 15126 7590 15138 7642
rect 15190 7590 15202 7642
rect 15254 7590 15266 7642
rect 15318 7590 21010 7642
rect 21062 7590 21074 7642
rect 21126 7590 21138 7642
rect 21190 7590 21202 7642
rect 21254 7590 21266 7642
rect 21318 7590 27010 7642
rect 27062 7590 27074 7642
rect 27126 7590 27138 7642
rect 27190 7590 27202 7642
rect 27254 7590 27266 7642
rect 27318 7590 33010 7642
rect 33062 7590 33074 7642
rect 33126 7590 33138 7642
rect 33190 7590 33202 7642
rect 33254 7590 33266 7642
rect 33318 7590 39010 7642
rect 39062 7590 39074 7642
rect 39126 7590 39138 7642
rect 39190 7590 39202 7642
rect 39254 7590 39266 7642
rect 39318 7590 45010 7642
rect 45062 7590 45074 7642
rect 45126 7590 45138 7642
rect 45190 7590 45202 7642
rect 45254 7590 45266 7642
rect 45318 7590 47840 7642
rect 1104 7568 47840 7590
rect 4154 7488 4160 7540
rect 4212 7528 4218 7540
rect 13722 7528 13728 7540
rect 4212 7500 13728 7528
rect 4212 7488 4218 7500
rect 13722 7488 13728 7500
rect 13780 7488 13786 7540
rect 14645 7531 14703 7537
rect 14645 7497 14657 7531
rect 14691 7528 14703 7531
rect 15470 7528 15476 7540
rect 14691 7500 15476 7528
rect 14691 7497 14703 7500
rect 14645 7491 14703 7497
rect 15470 7488 15476 7500
rect 15528 7488 15534 7540
rect 15657 7531 15715 7537
rect 15657 7497 15669 7531
rect 15703 7528 15715 7531
rect 15838 7528 15844 7540
rect 15703 7500 15844 7528
rect 15703 7497 15715 7500
rect 15657 7491 15715 7497
rect 15838 7488 15844 7500
rect 15896 7488 15902 7540
rect 15933 7531 15991 7537
rect 15933 7497 15945 7531
rect 15979 7528 15991 7531
rect 16206 7528 16212 7540
rect 15979 7500 16212 7528
rect 15979 7497 15991 7500
rect 15933 7491 15991 7497
rect 16206 7488 16212 7500
rect 16264 7488 16270 7540
rect 16942 7488 16948 7540
rect 17000 7528 17006 7540
rect 17129 7531 17187 7537
rect 17129 7528 17141 7531
rect 17000 7500 17141 7528
rect 17000 7488 17006 7500
rect 17129 7497 17141 7500
rect 17175 7497 17187 7531
rect 17129 7491 17187 7497
rect 22005 7531 22063 7537
rect 22005 7497 22017 7531
rect 22051 7497 22063 7531
rect 22005 7491 22063 7497
rect 7742 7420 7748 7472
rect 7800 7420 7806 7472
rect 7929 7463 7987 7469
rect 7929 7429 7941 7463
rect 7975 7460 7987 7463
rect 8294 7460 8300 7472
rect 7975 7432 8300 7460
rect 7975 7429 7987 7432
rect 7929 7423 7987 7429
rect 8294 7420 8300 7432
rect 8352 7420 8358 7472
rect 15105 7463 15163 7469
rect 15105 7429 15117 7463
rect 15151 7460 15163 7463
rect 15151 7432 15792 7460
rect 15151 7429 15163 7432
rect 15105 7423 15163 7429
rect 14461 7395 14519 7401
rect 14461 7361 14473 7395
rect 14507 7392 14519 7395
rect 14918 7392 14924 7404
rect 14507 7364 14924 7392
rect 14507 7361 14519 7364
rect 14461 7355 14519 7361
rect 14918 7352 14924 7364
rect 14976 7352 14982 7404
rect 15289 7395 15347 7401
rect 15470 7396 15476 7404
rect 15289 7361 15301 7395
rect 15335 7392 15347 7395
rect 15396 7392 15476 7396
rect 15528 7401 15534 7404
rect 15764 7401 15792 7432
rect 16482 7420 16488 7472
rect 16540 7460 16546 7472
rect 18874 7460 18880 7472
rect 16540 7432 18880 7460
rect 16540 7420 16546 7432
rect 18874 7420 18880 7432
rect 18932 7420 18938 7472
rect 22020 7460 22048 7491
rect 30558 7488 30564 7540
rect 30616 7528 30622 7540
rect 39574 7528 39580 7540
rect 30616 7500 39580 7528
rect 30616 7488 30622 7500
rect 39574 7488 39580 7500
rect 39632 7488 39638 7540
rect 41969 7531 42027 7537
rect 41969 7497 41981 7531
rect 42015 7528 42027 7531
rect 44082 7528 44088 7540
rect 42015 7500 44088 7528
rect 42015 7497 42027 7500
rect 41969 7491 42027 7497
rect 44082 7488 44088 7500
rect 44140 7488 44146 7540
rect 44542 7488 44548 7540
rect 44600 7488 44606 7540
rect 45281 7531 45339 7537
rect 45281 7497 45293 7531
rect 45327 7528 45339 7531
rect 46198 7528 46204 7540
rect 45327 7500 46204 7528
rect 45327 7497 45339 7500
rect 45281 7491 45339 7497
rect 46198 7488 46204 7500
rect 46256 7488 46262 7540
rect 46566 7488 46572 7540
rect 46624 7488 46630 7540
rect 46934 7488 46940 7540
rect 46992 7488 46998 7540
rect 47302 7488 47308 7540
rect 47360 7488 47366 7540
rect 25498 7460 25504 7472
rect 22020 7432 25504 7460
rect 25498 7420 25504 7432
rect 25556 7420 25562 7472
rect 35894 7420 35900 7472
rect 35952 7460 35958 7472
rect 35952 7432 43392 7460
rect 35952 7420 35958 7432
rect 15335 7368 15476 7392
rect 15335 7364 15424 7368
rect 15335 7361 15347 7364
rect 15289 7355 15347 7361
rect 15470 7352 15476 7368
rect 15528 7392 15539 7401
rect 15749 7395 15807 7401
rect 15528 7364 15621 7392
rect 15528 7355 15539 7364
rect 15749 7361 15761 7395
rect 15795 7392 15807 7395
rect 16574 7392 16580 7404
rect 15795 7364 16580 7392
rect 15795 7361 15807 7364
rect 15749 7355 15807 7361
rect 15528 7352 15534 7355
rect 16574 7352 16580 7364
rect 16632 7352 16638 7404
rect 17313 7395 17371 7401
rect 17313 7361 17325 7395
rect 17359 7392 17371 7395
rect 19150 7392 19156 7404
rect 17359 7364 19156 7392
rect 17359 7361 17371 7364
rect 17313 7355 17371 7361
rect 19150 7352 19156 7364
rect 19208 7352 19214 7404
rect 20714 7352 20720 7404
rect 20772 7392 20778 7404
rect 21821 7395 21879 7401
rect 21821 7392 21833 7395
rect 20772 7364 21833 7392
rect 20772 7352 20778 7364
rect 21821 7361 21833 7364
rect 21867 7361 21879 7395
rect 21821 7355 21879 7361
rect 26326 7352 26332 7404
rect 26384 7392 26390 7404
rect 26605 7395 26663 7401
rect 26605 7392 26617 7395
rect 26384 7364 26617 7392
rect 26384 7352 26390 7364
rect 26605 7361 26617 7364
rect 26651 7361 26663 7395
rect 26605 7355 26663 7361
rect 32306 7352 32312 7404
rect 32364 7392 32370 7404
rect 43364 7401 43392 7432
rect 43622 7420 43628 7472
rect 43680 7460 43686 7472
rect 43680 7432 46428 7460
rect 43680 7420 43686 7432
rect 33505 7395 33563 7401
rect 33505 7392 33517 7395
rect 32364 7364 33517 7392
rect 32364 7352 32370 7364
rect 33505 7361 33517 7364
rect 33551 7361 33563 7395
rect 33505 7355 33563 7361
rect 41693 7395 41751 7401
rect 41693 7361 41705 7395
rect 41739 7392 41751 7395
rect 41785 7395 41843 7401
rect 41785 7392 41797 7395
rect 41739 7364 41797 7392
rect 41739 7361 41751 7364
rect 41693 7355 41751 7361
rect 41785 7361 41797 7364
rect 41831 7361 41843 7395
rect 41785 7355 41843 7361
rect 42521 7395 42579 7401
rect 42521 7361 42533 7395
rect 42567 7361 42579 7395
rect 42521 7355 42579 7361
rect 43349 7395 43407 7401
rect 43349 7361 43361 7395
rect 43395 7361 43407 7395
rect 43349 7355 43407 7361
rect 44361 7395 44419 7401
rect 44361 7361 44373 7395
rect 44407 7361 44419 7395
rect 44361 7355 44419 7361
rect 45097 7395 45155 7401
rect 45097 7361 45109 7395
rect 45143 7361 45155 7395
rect 45097 7355 45155 7361
rect 6730 7284 6736 7336
rect 6788 7324 6794 7336
rect 15378 7324 15384 7336
rect 6788 7296 15384 7324
rect 6788 7284 6794 7296
rect 15378 7284 15384 7296
rect 15436 7284 15442 7336
rect 15654 7284 15660 7336
rect 15712 7324 15718 7336
rect 28258 7324 28264 7336
rect 15712 7296 28264 7324
rect 15712 7284 15718 7296
rect 28258 7284 28264 7296
rect 28316 7284 28322 7336
rect 40494 7284 40500 7336
rect 40552 7324 40558 7336
rect 42536 7324 42564 7355
rect 40552 7296 42564 7324
rect 40552 7284 40558 7296
rect 42794 7284 42800 7336
rect 42852 7324 42858 7336
rect 44376 7324 44404 7355
rect 42852 7296 44404 7324
rect 45112 7324 45140 7355
rect 45370 7352 45376 7404
rect 45428 7352 45434 7404
rect 45646 7352 45652 7404
rect 45704 7352 45710 7404
rect 45738 7352 45744 7404
rect 45796 7392 45802 7404
rect 46400 7401 46428 7432
rect 46017 7395 46075 7401
rect 46017 7392 46029 7395
rect 45796 7364 46029 7392
rect 45796 7352 45802 7364
rect 46017 7361 46029 7364
rect 46063 7361 46075 7395
rect 46017 7355 46075 7361
rect 46385 7395 46443 7401
rect 46385 7361 46397 7395
rect 46431 7361 46443 7395
rect 46385 7355 46443 7361
rect 46750 7352 46756 7404
rect 46808 7352 46814 7404
rect 47118 7352 47124 7404
rect 47176 7352 47182 7404
rect 47210 7324 47216 7336
rect 45112 7296 47216 7324
rect 42852 7284 42858 7296
rect 47210 7284 47216 7296
rect 47268 7284 47274 7336
rect 7650 7216 7656 7268
rect 7708 7256 7714 7268
rect 26421 7259 26479 7265
rect 26421 7256 26433 7259
rect 7708 7228 14964 7256
rect 7708 7216 7714 7228
rect 11238 7148 11244 7200
rect 11296 7188 11302 7200
rect 14826 7188 14832 7200
rect 11296 7160 14832 7188
rect 11296 7148 11302 7160
rect 14826 7148 14832 7160
rect 14884 7148 14890 7200
rect 14936 7188 14964 7228
rect 15580 7228 26433 7256
rect 15580 7188 15608 7228
rect 26421 7225 26433 7228
rect 26467 7225 26479 7259
rect 26421 7219 26479 7225
rect 42705 7259 42763 7265
rect 42705 7225 42717 7259
rect 42751 7256 42763 7259
rect 42886 7256 42892 7268
rect 42751 7228 42892 7256
rect 42751 7225 42763 7228
rect 42705 7219 42763 7225
rect 42886 7216 42892 7228
rect 42944 7216 42950 7268
rect 43533 7259 43591 7265
rect 43533 7225 43545 7259
rect 43579 7256 43591 7259
rect 45462 7256 45468 7268
rect 43579 7228 45468 7256
rect 43579 7225 43591 7228
rect 43533 7219 43591 7225
rect 45462 7216 45468 7228
rect 45520 7216 45526 7268
rect 45557 7259 45615 7265
rect 45557 7225 45569 7259
rect 45603 7256 45615 7259
rect 46658 7256 46664 7268
rect 45603 7228 46664 7256
rect 45603 7225 45615 7228
rect 45557 7219 45615 7225
rect 46658 7216 46664 7228
rect 46716 7216 46722 7268
rect 14936 7160 15608 7188
rect 16298 7148 16304 7200
rect 16356 7188 16362 7200
rect 29822 7188 29828 7200
rect 16356 7160 29828 7188
rect 16356 7148 16362 7160
rect 29822 7148 29828 7160
rect 29880 7148 29886 7200
rect 33318 7148 33324 7200
rect 33376 7148 33382 7200
rect 41598 7148 41604 7200
rect 41656 7148 41662 7200
rect 45833 7191 45891 7197
rect 45833 7157 45845 7191
rect 45879 7188 45891 7191
rect 45922 7188 45928 7200
rect 45879 7160 45928 7188
rect 45879 7157 45891 7160
rect 45833 7151 45891 7157
rect 45922 7148 45928 7160
rect 45980 7148 45986 7200
rect 46201 7191 46259 7197
rect 46201 7157 46213 7191
rect 46247 7188 46259 7191
rect 46290 7188 46296 7200
rect 46247 7160 46296 7188
rect 46247 7157 46259 7160
rect 46201 7151 46259 7157
rect 46290 7148 46296 7160
rect 46348 7148 46354 7200
rect 1104 7098 47840 7120
rect 1104 7046 1950 7098
rect 2002 7046 2014 7098
rect 2066 7046 2078 7098
rect 2130 7046 2142 7098
rect 2194 7046 2206 7098
rect 2258 7046 7950 7098
rect 8002 7046 8014 7098
rect 8066 7046 8078 7098
rect 8130 7046 8142 7098
rect 8194 7046 8206 7098
rect 8258 7046 13950 7098
rect 14002 7046 14014 7098
rect 14066 7046 14078 7098
rect 14130 7046 14142 7098
rect 14194 7046 14206 7098
rect 14258 7046 19950 7098
rect 20002 7046 20014 7098
rect 20066 7046 20078 7098
rect 20130 7046 20142 7098
rect 20194 7046 20206 7098
rect 20258 7046 25950 7098
rect 26002 7046 26014 7098
rect 26066 7046 26078 7098
rect 26130 7046 26142 7098
rect 26194 7046 26206 7098
rect 26258 7046 31950 7098
rect 32002 7046 32014 7098
rect 32066 7046 32078 7098
rect 32130 7046 32142 7098
rect 32194 7046 32206 7098
rect 32258 7046 37950 7098
rect 38002 7046 38014 7098
rect 38066 7046 38078 7098
rect 38130 7046 38142 7098
rect 38194 7046 38206 7098
rect 38258 7046 43950 7098
rect 44002 7046 44014 7098
rect 44066 7046 44078 7098
rect 44130 7046 44142 7098
rect 44194 7046 44206 7098
rect 44258 7046 47840 7098
rect 1104 7024 47840 7046
rect 12526 6944 12532 6996
rect 12584 6984 12590 6996
rect 19334 6984 19340 6996
rect 12584 6956 19340 6984
rect 12584 6944 12590 6956
rect 19334 6944 19340 6956
rect 19392 6944 19398 6996
rect 36906 6944 36912 6996
rect 36964 6984 36970 6996
rect 45830 6984 45836 6996
rect 36964 6956 45836 6984
rect 36964 6944 36970 6956
rect 45830 6944 45836 6956
rect 45888 6944 45894 6996
rect 14826 6876 14832 6928
rect 14884 6916 14890 6928
rect 33318 6916 33324 6928
rect 14884 6888 33324 6916
rect 14884 6876 14890 6888
rect 33318 6876 33324 6888
rect 33376 6876 33382 6928
rect 13630 6808 13636 6860
rect 13688 6848 13694 6860
rect 13688 6820 16528 6848
rect 13688 6808 13694 6820
rect 15473 6783 15531 6789
rect 15473 6749 15485 6783
rect 15519 6780 15531 6783
rect 15565 6783 15623 6789
rect 15565 6780 15577 6783
rect 15519 6752 15577 6780
rect 15519 6749 15531 6752
rect 15473 6743 15531 6749
rect 15565 6749 15577 6752
rect 15611 6780 15623 6783
rect 16022 6780 16028 6792
rect 15611 6752 16028 6780
rect 15611 6749 15623 6752
rect 15565 6743 15623 6749
rect 16022 6740 16028 6752
rect 16080 6740 16086 6792
rect 16209 6783 16267 6789
rect 16209 6749 16221 6783
rect 16255 6780 16267 6783
rect 16301 6783 16359 6789
rect 16301 6780 16313 6783
rect 16255 6752 16313 6780
rect 16255 6749 16267 6752
rect 16209 6743 16267 6749
rect 16301 6749 16313 6752
rect 16347 6780 16359 6783
rect 16390 6780 16396 6792
rect 16347 6752 16396 6780
rect 16347 6749 16359 6752
rect 16301 6743 16359 6749
rect 16390 6740 16396 6752
rect 16448 6740 16454 6792
rect 16500 6780 16528 6820
rect 17770 6808 17776 6860
rect 17828 6848 17834 6860
rect 39390 6848 39396 6860
rect 17828 6820 39396 6848
rect 17828 6808 17834 6820
rect 39390 6808 39396 6820
rect 39448 6808 39454 6860
rect 43714 6808 43720 6860
rect 43772 6848 43778 6860
rect 43772 6820 46888 6848
rect 43772 6808 43778 6820
rect 23477 6783 23535 6789
rect 23477 6780 23489 6783
rect 16500 6752 23489 6780
rect 23477 6749 23489 6752
rect 23523 6749 23535 6783
rect 23477 6743 23535 6749
rect 29365 6783 29423 6789
rect 29365 6749 29377 6783
rect 29411 6780 29423 6783
rect 30282 6780 30288 6792
rect 29411 6752 30288 6780
rect 29411 6749 29423 6752
rect 29365 6743 29423 6749
rect 30282 6740 30288 6752
rect 30340 6740 30346 6792
rect 31754 6740 31760 6792
rect 31812 6780 31818 6792
rect 32493 6783 32551 6789
rect 32493 6780 32505 6783
rect 31812 6752 32505 6780
rect 31812 6740 31818 6752
rect 32493 6749 32505 6752
rect 32539 6749 32551 6783
rect 32493 6743 32551 6749
rect 32858 6740 32864 6792
rect 32916 6780 32922 6792
rect 35529 6783 35587 6789
rect 35529 6780 35541 6783
rect 32916 6752 35541 6780
rect 32916 6740 32922 6752
rect 35529 6749 35541 6752
rect 35575 6749 35587 6783
rect 35529 6743 35587 6749
rect 45554 6740 45560 6792
rect 45612 6780 45618 6792
rect 45649 6783 45707 6789
rect 45649 6780 45661 6783
rect 45612 6752 45661 6780
rect 45612 6740 45618 6752
rect 45649 6749 45661 6752
rect 45695 6780 45707 6783
rect 45833 6783 45891 6789
rect 45833 6780 45845 6783
rect 45695 6752 45845 6780
rect 45695 6749 45707 6752
rect 45649 6743 45707 6749
rect 45833 6749 45845 6752
rect 45879 6749 45891 6783
rect 45833 6743 45891 6749
rect 46106 6740 46112 6792
rect 46164 6740 46170 6792
rect 46198 6740 46204 6792
rect 46256 6780 46262 6792
rect 46860 6789 46888 6820
rect 46477 6783 46535 6789
rect 46477 6780 46489 6783
rect 46256 6752 46489 6780
rect 46256 6740 46262 6752
rect 46477 6749 46489 6752
rect 46523 6749 46535 6783
rect 46477 6743 46535 6749
rect 46845 6783 46903 6789
rect 46845 6749 46857 6783
rect 46891 6749 46903 6783
rect 46845 6743 46903 6749
rect 47213 6783 47271 6789
rect 47213 6749 47225 6783
rect 47259 6749 47271 6783
rect 47213 6743 47271 6749
rect 16758 6712 16764 6724
rect 15764 6684 16764 6712
rect 15764 6653 15792 6684
rect 16758 6672 16764 6684
rect 16816 6672 16822 6724
rect 17218 6672 17224 6724
rect 17276 6712 17282 6724
rect 17276 6684 29224 6712
rect 17276 6672 17282 6684
rect 15749 6647 15807 6653
rect 15749 6613 15761 6647
rect 15795 6613 15807 6647
rect 15749 6607 15807 6613
rect 16485 6647 16543 6653
rect 16485 6613 16497 6647
rect 16531 6644 16543 6647
rect 17126 6644 17132 6656
rect 16531 6616 17132 6644
rect 16531 6613 16543 6616
rect 16485 6607 16543 6613
rect 17126 6604 17132 6616
rect 17184 6604 17190 6656
rect 23658 6604 23664 6656
rect 23716 6604 23722 6656
rect 29196 6653 29224 6684
rect 32766 6672 32772 6724
rect 32824 6712 32830 6724
rect 47228 6712 47256 6743
rect 32824 6684 47256 6712
rect 32824 6672 32830 6684
rect 29181 6647 29239 6653
rect 29181 6613 29193 6647
rect 29227 6613 29239 6647
rect 29181 6607 29239 6613
rect 29270 6604 29276 6656
rect 29328 6644 29334 6656
rect 32309 6647 32367 6653
rect 32309 6644 32321 6647
rect 29328 6616 32321 6644
rect 29328 6604 29334 6616
rect 32309 6613 32321 6616
rect 32355 6613 32367 6647
rect 32309 6607 32367 6613
rect 35342 6604 35348 6656
rect 35400 6604 35406 6656
rect 46014 6604 46020 6656
rect 46072 6604 46078 6656
rect 46290 6604 46296 6656
rect 46348 6604 46354 6656
rect 46658 6604 46664 6656
rect 46716 6604 46722 6656
rect 47026 6604 47032 6656
rect 47084 6604 47090 6656
rect 47394 6604 47400 6656
rect 47452 6604 47458 6656
rect 1104 6554 47840 6576
rect 1104 6502 3010 6554
rect 3062 6502 3074 6554
rect 3126 6502 3138 6554
rect 3190 6502 3202 6554
rect 3254 6502 3266 6554
rect 3318 6502 9010 6554
rect 9062 6502 9074 6554
rect 9126 6502 9138 6554
rect 9190 6502 9202 6554
rect 9254 6502 9266 6554
rect 9318 6502 15010 6554
rect 15062 6502 15074 6554
rect 15126 6502 15138 6554
rect 15190 6502 15202 6554
rect 15254 6502 15266 6554
rect 15318 6502 21010 6554
rect 21062 6502 21074 6554
rect 21126 6502 21138 6554
rect 21190 6502 21202 6554
rect 21254 6502 21266 6554
rect 21318 6502 27010 6554
rect 27062 6502 27074 6554
rect 27126 6502 27138 6554
rect 27190 6502 27202 6554
rect 27254 6502 27266 6554
rect 27318 6502 33010 6554
rect 33062 6502 33074 6554
rect 33126 6502 33138 6554
rect 33190 6502 33202 6554
rect 33254 6502 33266 6554
rect 33318 6502 39010 6554
rect 39062 6502 39074 6554
rect 39126 6502 39138 6554
rect 39190 6502 39202 6554
rect 39254 6502 39266 6554
rect 39318 6502 45010 6554
rect 45062 6502 45074 6554
rect 45126 6502 45138 6554
rect 45190 6502 45202 6554
rect 45254 6502 45266 6554
rect 45318 6502 47840 6554
rect 1104 6480 47840 6502
rect 12710 6400 12716 6452
rect 12768 6440 12774 6452
rect 17218 6440 17224 6452
rect 12768 6412 17224 6440
rect 12768 6400 12774 6412
rect 17218 6400 17224 6412
rect 17276 6400 17282 6452
rect 23658 6400 23664 6452
rect 23716 6440 23722 6452
rect 23716 6412 36492 6440
rect 23716 6400 23722 6412
rect 10962 6332 10968 6384
rect 11020 6372 11026 6384
rect 29270 6372 29276 6384
rect 11020 6344 29276 6372
rect 11020 6332 11026 6344
rect 29270 6332 29276 6344
rect 29328 6332 29334 6384
rect 33410 6332 33416 6384
rect 33468 6372 33474 6384
rect 36357 6375 36415 6381
rect 36357 6372 36369 6375
rect 33468 6344 36369 6372
rect 33468 6332 33474 6344
rect 36357 6341 36369 6344
rect 36403 6341 36415 6375
rect 36464 6372 36492 6412
rect 38562 6400 38568 6452
rect 38620 6440 38626 6452
rect 39669 6443 39727 6449
rect 39669 6440 39681 6443
rect 38620 6412 39681 6440
rect 38620 6400 38626 6412
rect 39669 6409 39681 6412
rect 39715 6409 39727 6443
rect 39669 6403 39727 6409
rect 41386 6412 46796 6440
rect 40034 6372 40040 6384
rect 36464 6344 40040 6372
rect 36357 6335 36415 6341
rect 40034 6332 40040 6344
rect 40092 6332 40098 6384
rect 16850 6264 16856 6316
rect 16908 6304 16914 6316
rect 24486 6304 24492 6316
rect 16908 6276 24492 6304
rect 16908 6264 16914 6276
rect 24486 6264 24492 6276
rect 24544 6264 24550 6316
rect 24673 6307 24731 6313
rect 24673 6273 24685 6307
rect 24719 6304 24731 6307
rect 25130 6304 25136 6316
rect 24719 6276 25136 6304
rect 24719 6273 24731 6276
rect 24673 6267 24731 6273
rect 25130 6264 25136 6276
rect 25188 6264 25194 6316
rect 25409 6307 25467 6313
rect 25409 6273 25421 6307
rect 25455 6304 25467 6307
rect 25501 6307 25559 6313
rect 25501 6304 25513 6307
rect 25455 6276 25513 6304
rect 25455 6273 25467 6276
rect 25409 6267 25467 6273
rect 25501 6273 25513 6276
rect 25547 6273 25559 6307
rect 25501 6267 25559 6273
rect 25590 6264 25596 6316
rect 25648 6304 25654 6316
rect 25961 6307 26019 6313
rect 25961 6304 25973 6307
rect 25648 6276 25973 6304
rect 25648 6264 25654 6276
rect 25961 6273 25973 6276
rect 26007 6273 26019 6307
rect 25961 6267 26019 6273
rect 26421 6307 26479 6313
rect 26421 6273 26433 6307
rect 26467 6273 26479 6307
rect 26421 6267 26479 6273
rect 7834 6196 7840 6248
rect 7892 6236 7898 6248
rect 25774 6236 25780 6248
rect 7892 6208 25780 6236
rect 7892 6196 7898 6208
rect 25774 6196 25780 6208
rect 25832 6196 25838 6248
rect 25866 6196 25872 6248
rect 25924 6236 25930 6248
rect 26436 6236 26464 6267
rect 32398 6264 32404 6316
rect 32456 6304 32462 6316
rect 32953 6307 33011 6313
rect 32953 6304 32965 6307
rect 32456 6276 32965 6304
rect 32456 6264 32462 6276
rect 32953 6273 32965 6276
rect 32999 6273 33011 6307
rect 32953 6267 33011 6273
rect 34330 6264 34336 6316
rect 34388 6304 34394 6316
rect 39853 6307 39911 6313
rect 39853 6304 39865 6307
rect 34388 6276 39865 6304
rect 34388 6264 34394 6276
rect 39853 6273 39865 6276
rect 39899 6273 39911 6307
rect 39853 6267 39911 6273
rect 25924 6208 26464 6236
rect 25924 6196 25930 6208
rect 26510 6196 26516 6248
rect 26568 6236 26574 6248
rect 41386 6236 41414 6412
rect 46014 6332 46020 6384
rect 46072 6372 46078 6384
rect 46072 6344 46704 6372
rect 46072 6332 46078 6344
rect 46382 6264 46388 6316
rect 46440 6264 46446 6316
rect 26568 6208 41414 6236
rect 46676 6236 46704 6344
rect 46768 6313 46796 6412
rect 46934 6400 46940 6452
rect 46992 6400 46998 6452
rect 47305 6443 47363 6449
rect 47305 6409 47317 6443
rect 47351 6440 47363 6443
rect 47486 6440 47492 6452
rect 47351 6412 47492 6440
rect 47351 6409 47363 6412
rect 47305 6403 47363 6409
rect 47486 6400 47492 6412
rect 47544 6400 47550 6452
rect 46753 6307 46811 6313
rect 46753 6273 46765 6307
rect 46799 6273 46811 6307
rect 46753 6267 46811 6273
rect 47121 6307 47179 6313
rect 47121 6273 47133 6307
rect 47167 6273 47179 6307
rect 47121 6267 47179 6273
rect 47136 6236 47164 6267
rect 46676 6208 47164 6236
rect 26568 6196 26574 6208
rect 8386 6128 8392 6180
rect 8444 6168 8450 6180
rect 25685 6171 25743 6177
rect 8444 6140 25452 6168
rect 8444 6128 8450 6140
rect 6822 6060 6828 6112
rect 6880 6100 6886 6112
rect 22462 6100 22468 6112
rect 6880 6072 22468 6100
rect 6880 6060 6886 6072
rect 22462 6060 22468 6072
rect 22520 6060 22526 6112
rect 24486 6060 24492 6112
rect 24544 6060 24550 6112
rect 24670 6060 24676 6112
rect 24728 6100 24734 6112
rect 25317 6103 25375 6109
rect 25317 6100 25329 6103
rect 24728 6072 25329 6100
rect 24728 6060 24734 6072
rect 25317 6069 25329 6072
rect 25363 6069 25375 6103
rect 25424 6100 25452 6140
rect 25685 6137 25697 6171
rect 25731 6168 25743 6171
rect 34422 6168 34428 6180
rect 25731 6140 34428 6168
rect 25731 6137 25743 6140
rect 25685 6131 25743 6137
rect 34422 6128 34428 6140
rect 34480 6128 34486 6180
rect 36170 6128 36176 6180
rect 36228 6128 36234 6180
rect 36262 6128 36268 6180
rect 36320 6168 36326 6180
rect 46198 6168 46204 6180
rect 36320 6140 46204 6168
rect 36320 6128 36326 6140
rect 46198 6128 46204 6140
rect 46256 6128 46262 6180
rect 25777 6103 25835 6109
rect 25777 6100 25789 6103
rect 25424 6072 25789 6100
rect 25317 6063 25375 6069
rect 25777 6069 25789 6072
rect 25823 6069 25835 6103
rect 25777 6063 25835 6069
rect 25866 6060 25872 6112
rect 25924 6100 25930 6112
rect 26237 6103 26295 6109
rect 26237 6100 26249 6103
rect 25924 6072 26249 6100
rect 25924 6060 25930 6072
rect 26237 6069 26249 6072
rect 26283 6069 26295 6103
rect 26237 6063 26295 6069
rect 33134 6060 33140 6112
rect 33192 6060 33198 6112
rect 46566 6060 46572 6112
rect 46624 6060 46630 6112
rect 1104 6010 47840 6032
rect 1104 5958 1950 6010
rect 2002 5958 2014 6010
rect 2066 5958 2078 6010
rect 2130 5958 2142 6010
rect 2194 5958 2206 6010
rect 2258 5958 7950 6010
rect 8002 5958 8014 6010
rect 8066 5958 8078 6010
rect 8130 5958 8142 6010
rect 8194 5958 8206 6010
rect 8258 5958 13950 6010
rect 14002 5958 14014 6010
rect 14066 5958 14078 6010
rect 14130 5958 14142 6010
rect 14194 5958 14206 6010
rect 14258 5958 19950 6010
rect 20002 5958 20014 6010
rect 20066 5958 20078 6010
rect 20130 5958 20142 6010
rect 20194 5958 20206 6010
rect 20258 5958 25950 6010
rect 26002 5958 26014 6010
rect 26066 5958 26078 6010
rect 26130 5958 26142 6010
rect 26194 5958 26206 6010
rect 26258 5958 31950 6010
rect 32002 5958 32014 6010
rect 32066 5958 32078 6010
rect 32130 5958 32142 6010
rect 32194 5958 32206 6010
rect 32258 5958 37950 6010
rect 38002 5958 38014 6010
rect 38066 5958 38078 6010
rect 38130 5958 38142 6010
rect 38194 5958 38206 6010
rect 38258 5958 43950 6010
rect 44002 5958 44014 6010
rect 44066 5958 44078 6010
rect 44130 5958 44142 6010
rect 44194 5958 44206 6010
rect 44258 5958 47840 6010
rect 1104 5936 47840 5958
rect 11054 5856 11060 5908
rect 11112 5896 11118 5908
rect 14461 5899 14519 5905
rect 14461 5896 14473 5899
rect 11112 5868 14473 5896
rect 11112 5856 11118 5868
rect 14461 5865 14473 5868
rect 14507 5865 14519 5899
rect 14461 5859 14519 5865
rect 17770 5856 17776 5908
rect 17828 5856 17834 5908
rect 22462 5856 22468 5908
rect 22520 5856 22526 5908
rect 27614 5856 27620 5908
rect 27672 5896 27678 5908
rect 27672 5868 31156 5896
rect 27672 5856 27678 5868
rect 12618 5788 12624 5840
rect 12676 5828 12682 5840
rect 28813 5831 28871 5837
rect 28813 5828 28825 5831
rect 12676 5800 28825 5828
rect 12676 5788 12682 5800
rect 28813 5797 28825 5800
rect 28859 5797 28871 5831
rect 28813 5791 28871 5797
rect 30193 5831 30251 5837
rect 30193 5797 30205 5831
rect 30239 5797 30251 5831
rect 31128 5828 31156 5868
rect 31202 5856 31208 5908
rect 31260 5896 31266 5908
rect 46382 5896 46388 5908
rect 31260 5868 46388 5896
rect 31260 5856 31266 5868
rect 46382 5856 46388 5868
rect 46440 5856 46446 5908
rect 47394 5856 47400 5908
rect 47452 5856 47458 5908
rect 36262 5828 36268 5840
rect 31128 5800 36268 5828
rect 30193 5791 30251 5797
rect 12802 5720 12808 5772
rect 12860 5760 12866 5772
rect 12860 5732 15056 5760
rect 12860 5720 12866 5732
rect 14553 5695 14611 5701
rect 14553 5661 14565 5695
rect 14599 5692 14611 5695
rect 14737 5695 14795 5701
rect 14737 5692 14749 5695
rect 14599 5664 14749 5692
rect 14599 5661 14611 5664
rect 14553 5655 14611 5661
rect 14737 5661 14749 5664
rect 14783 5661 14795 5695
rect 14737 5655 14795 5661
rect 14918 5652 14924 5704
rect 14976 5652 14982 5704
rect 15028 5692 15056 5732
rect 19334 5720 19340 5772
rect 19392 5760 19398 5772
rect 30208 5760 30236 5791
rect 36262 5788 36268 5800
rect 36320 5788 36326 5840
rect 37182 5788 37188 5840
rect 37240 5828 37246 5840
rect 38933 5831 38991 5837
rect 38933 5828 38945 5831
rect 37240 5800 38945 5828
rect 37240 5788 37246 5800
rect 38933 5797 38945 5800
rect 38979 5797 38991 5831
rect 38933 5791 38991 5797
rect 30650 5760 30656 5772
rect 19392 5732 30236 5760
rect 30300 5732 30656 5760
rect 19392 5720 19398 5732
rect 22649 5695 22707 5701
rect 15028 5664 22094 5692
rect 17497 5627 17555 5633
rect 17497 5593 17509 5627
rect 17543 5624 17555 5627
rect 17681 5627 17739 5633
rect 17681 5624 17693 5627
rect 17543 5596 17693 5624
rect 17543 5593 17555 5596
rect 17497 5587 17555 5593
rect 17681 5593 17693 5596
rect 17727 5593 17739 5627
rect 17681 5587 17739 5593
rect 17402 5516 17408 5568
rect 17460 5516 17466 5568
rect 22066 5556 22094 5664
rect 22649 5661 22661 5695
rect 22695 5692 22707 5695
rect 24394 5692 24400 5704
rect 22695 5664 24400 5692
rect 22695 5661 22707 5664
rect 22649 5655 22707 5661
rect 24394 5652 24400 5664
rect 24452 5652 24458 5704
rect 28997 5695 29055 5701
rect 28997 5661 29009 5695
rect 29043 5692 29055 5695
rect 30300 5692 30328 5732
rect 30650 5720 30656 5732
rect 30708 5720 30714 5772
rect 33134 5720 33140 5772
rect 33192 5760 33198 5772
rect 43622 5760 43628 5772
rect 33192 5732 43628 5760
rect 33192 5720 33198 5732
rect 43622 5720 43628 5732
rect 43680 5720 43686 5772
rect 29043 5664 30328 5692
rect 30377 5695 30435 5701
rect 29043 5661 29055 5664
rect 28997 5655 29055 5661
rect 30377 5661 30389 5695
rect 30423 5692 30435 5695
rect 31018 5692 31024 5704
rect 30423 5664 31024 5692
rect 30423 5661 30435 5664
rect 30377 5655 30435 5661
rect 31018 5652 31024 5664
rect 31076 5652 31082 5704
rect 31386 5652 31392 5704
rect 31444 5692 31450 5704
rect 31665 5695 31723 5701
rect 31665 5692 31677 5695
rect 31444 5664 31677 5692
rect 31444 5652 31450 5664
rect 31665 5661 31677 5664
rect 31711 5661 31723 5695
rect 31665 5655 31723 5661
rect 33962 5652 33968 5704
rect 34020 5692 34026 5704
rect 39117 5695 39175 5701
rect 39117 5692 39129 5695
rect 34020 5664 39129 5692
rect 34020 5652 34026 5664
rect 39117 5661 39129 5664
rect 39163 5661 39175 5695
rect 39117 5655 39175 5661
rect 39390 5652 39396 5704
rect 39448 5692 39454 5704
rect 46845 5695 46903 5701
rect 46845 5692 46857 5695
rect 39448 5664 46857 5692
rect 39448 5652 39454 5664
rect 46845 5661 46857 5664
rect 46891 5661 46903 5695
rect 46845 5655 46903 5661
rect 47213 5695 47271 5701
rect 47213 5661 47225 5695
rect 47259 5661 47271 5695
rect 47213 5655 47271 5661
rect 24946 5584 24952 5636
rect 25004 5624 25010 5636
rect 31202 5624 31208 5636
rect 25004 5596 31208 5624
rect 25004 5584 25010 5596
rect 31202 5584 31208 5596
rect 31260 5584 31266 5636
rect 44450 5584 44456 5636
rect 44508 5624 44514 5636
rect 47228 5624 47256 5655
rect 44508 5596 47256 5624
rect 44508 5584 44514 5596
rect 31481 5559 31539 5565
rect 31481 5556 31493 5559
rect 22066 5528 31493 5556
rect 31481 5525 31493 5528
rect 31527 5525 31539 5559
rect 31481 5519 31539 5525
rect 47026 5516 47032 5568
rect 47084 5516 47090 5568
rect 1104 5466 47840 5488
rect 1104 5414 3010 5466
rect 3062 5414 3074 5466
rect 3126 5414 3138 5466
rect 3190 5414 3202 5466
rect 3254 5414 3266 5466
rect 3318 5414 9010 5466
rect 9062 5414 9074 5466
rect 9126 5414 9138 5466
rect 9190 5414 9202 5466
rect 9254 5414 9266 5466
rect 9318 5414 15010 5466
rect 15062 5414 15074 5466
rect 15126 5414 15138 5466
rect 15190 5414 15202 5466
rect 15254 5414 15266 5466
rect 15318 5414 21010 5466
rect 21062 5414 21074 5466
rect 21126 5414 21138 5466
rect 21190 5414 21202 5466
rect 21254 5414 21266 5466
rect 21318 5414 27010 5466
rect 27062 5414 27074 5466
rect 27126 5414 27138 5466
rect 27190 5414 27202 5466
rect 27254 5414 27266 5466
rect 27318 5414 33010 5466
rect 33062 5414 33074 5466
rect 33126 5414 33138 5466
rect 33190 5414 33202 5466
rect 33254 5414 33266 5466
rect 33318 5414 39010 5466
rect 39062 5414 39074 5466
rect 39126 5414 39138 5466
rect 39190 5414 39202 5466
rect 39254 5414 39266 5466
rect 39318 5414 45010 5466
rect 45062 5414 45074 5466
rect 45126 5414 45138 5466
rect 45190 5414 45202 5466
rect 45254 5414 45266 5466
rect 45318 5414 47840 5466
rect 1104 5392 47840 5414
rect 13722 5312 13728 5364
rect 13780 5352 13786 5364
rect 21821 5355 21879 5361
rect 21821 5352 21833 5355
rect 13780 5324 21833 5352
rect 13780 5312 13786 5324
rect 21821 5321 21833 5324
rect 21867 5321 21879 5355
rect 21821 5315 21879 5321
rect 23382 5312 23388 5364
rect 23440 5352 23446 5364
rect 23661 5355 23719 5361
rect 23661 5352 23673 5355
rect 23440 5324 23673 5352
rect 23440 5312 23446 5324
rect 23661 5321 23673 5324
rect 23707 5321 23719 5355
rect 23661 5315 23719 5321
rect 26896 5324 47164 5352
rect 5994 5244 6000 5296
rect 6052 5284 6058 5296
rect 9217 5287 9275 5293
rect 9217 5284 9229 5287
rect 6052 5256 9229 5284
rect 6052 5244 6058 5256
rect 9217 5253 9229 5256
rect 9263 5253 9275 5287
rect 23566 5284 23572 5296
rect 9217 5247 9275 5253
rect 21560 5256 23572 5284
rect 9401 5219 9459 5225
rect 9401 5185 9413 5219
rect 9447 5216 9459 5219
rect 9582 5216 9588 5228
rect 9447 5188 9588 5216
rect 9447 5185 9459 5188
rect 9401 5179 9459 5185
rect 9582 5176 9588 5188
rect 9640 5176 9646 5228
rect 21560 5225 21588 5256
rect 23566 5244 23572 5256
rect 23624 5244 23630 5296
rect 21545 5219 21603 5225
rect 21545 5185 21557 5219
rect 21591 5185 21603 5219
rect 21545 5179 21603 5185
rect 21910 5176 21916 5228
rect 21968 5216 21974 5228
rect 22005 5219 22063 5225
rect 22005 5216 22017 5219
rect 21968 5188 22017 5216
rect 21968 5176 21974 5188
rect 22005 5185 22017 5188
rect 22051 5185 22063 5219
rect 22005 5179 22063 5185
rect 23845 5219 23903 5225
rect 23845 5185 23857 5219
rect 23891 5216 23903 5219
rect 24762 5216 24768 5228
rect 23891 5188 24768 5216
rect 23891 5185 23903 5188
rect 23845 5179 23903 5185
rect 24762 5176 24768 5188
rect 24820 5176 24826 5228
rect 18782 5108 18788 5160
rect 18840 5148 18846 5160
rect 26896 5148 26924 5324
rect 18840 5120 26924 5148
rect 31726 5256 41414 5284
rect 18840 5108 18846 5120
rect 18138 5040 18144 5092
rect 18196 5080 18202 5092
rect 18196 5052 21496 5080
rect 18196 5040 18202 5052
rect 20346 4972 20352 5024
rect 20404 5012 20410 5024
rect 21361 5015 21419 5021
rect 21361 5012 21373 5015
rect 20404 4984 21373 5012
rect 20404 4972 20410 4984
rect 21361 4981 21373 4984
rect 21407 4981 21419 5015
rect 21468 5012 21496 5052
rect 21726 5040 21732 5092
rect 21784 5080 21790 5092
rect 31726 5080 31754 5256
rect 33594 5176 33600 5228
rect 33652 5216 33658 5228
rect 37737 5219 37795 5225
rect 37737 5216 37749 5219
rect 33652 5188 37749 5216
rect 33652 5176 33658 5188
rect 37737 5185 37749 5188
rect 37783 5185 37795 5219
rect 41386 5216 41414 5256
rect 47136 5225 47164 5324
rect 47302 5312 47308 5364
rect 47360 5312 47366 5364
rect 46753 5219 46811 5225
rect 46753 5216 46765 5219
rect 41386 5188 46765 5216
rect 37737 5179 37795 5185
rect 46753 5185 46765 5188
rect 46799 5185 46811 5219
rect 46753 5179 46811 5185
rect 47121 5219 47179 5225
rect 47121 5185 47133 5219
rect 47167 5185 47179 5219
rect 47121 5179 47179 5185
rect 37550 5108 37556 5160
rect 37608 5108 37614 5160
rect 21784 5052 31754 5080
rect 21784 5040 21790 5052
rect 34422 5040 34428 5092
rect 34480 5080 34486 5092
rect 44358 5080 44364 5092
rect 34480 5052 44364 5080
rect 34480 5040 34486 5052
rect 44358 5040 44364 5052
rect 44416 5040 44422 5092
rect 27614 5012 27620 5024
rect 21468 4984 27620 5012
rect 21361 4975 21419 4981
rect 27614 4972 27620 4984
rect 27672 4972 27678 5024
rect 46934 4972 46940 5024
rect 46992 4972 46998 5024
rect 1104 4922 47840 4944
rect 1104 4870 1950 4922
rect 2002 4870 2014 4922
rect 2066 4870 2078 4922
rect 2130 4870 2142 4922
rect 2194 4870 2206 4922
rect 2258 4870 7950 4922
rect 8002 4870 8014 4922
rect 8066 4870 8078 4922
rect 8130 4870 8142 4922
rect 8194 4870 8206 4922
rect 8258 4870 13950 4922
rect 14002 4870 14014 4922
rect 14066 4870 14078 4922
rect 14130 4870 14142 4922
rect 14194 4870 14206 4922
rect 14258 4870 19950 4922
rect 20002 4870 20014 4922
rect 20066 4870 20078 4922
rect 20130 4870 20142 4922
rect 20194 4870 20206 4922
rect 20258 4870 25950 4922
rect 26002 4870 26014 4922
rect 26066 4870 26078 4922
rect 26130 4870 26142 4922
rect 26194 4870 26206 4922
rect 26258 4870 31950 4922
rect 32002 4870 32014 4922
rect 32066 4870 32078 4922
rect 32130 4870 32142 4922
rect 32194 4870 32206 4922
rect 32258 4870 37950 4922
rect 38002 4870 38014 4922
rect 38066 4870 38078 4922
rect 38130 4870 38142 4922
rect 38194 4870 38206 4922
rect 38258 4870 43950 4922
rect 44002 4870 44014 4922
rect 44066 4870 44078 4922
rect 44130 4870 44142 4922
rect 44194 4870 44206 4922
rect 44258 4870 47840 4922
rect 1104 4848 47840 4870
rect 18046 4768 18052 4820
rect 18104 4768 18110 4820
rect 19794 4768 19800 4820
rect 19852 4808 19858 4820
rect 20073 4811 20131 4817
rect 20073 4808 20085 4811
rect 19852 4780 20085 4808
rect 19852 4768 19858 4780
rect 20073 4777 20085 4780
rect 20119 4777 20131 4811
rect 20073 4771 20131 4777
rect 20441 4811 20499 4817
rect 20441 4777 20453 4811
rect 20487 4808 20499 4811
rect 24946 4808 24952 4820
rect 20487 4780 24952 4808
rect 20487 4777 20499 4780
rect 20441 4771 20499 4777
rect 24946 4768 24952 4780
rect 25004 4768 25010 4820
rect 47118 4808 47124 4820
rect 31726 4780 47124 4808
rect 8662 4700 8668 4752
rect 8720 4740 8726 4752
rect 20809 4743 20867 4749
rect 20809 4740 20821 4743
rect 8720 4712 20821 4740
rect 8720 4700 8726 4712
rect 20809 4709 20821 4712
rect 20855 4709 20867 4743
rect 23201 4743 23259 4749
rect 23201 4740 23213 4743
rect 20809 4703 20867 4709
rect 20916 4712 23213 4740
rect 17218 4632 17224 4684
rect 17276 4672 17282 4684
rect 20916 4672 20944 4712
rect 23201 4709 23213 4712
rect 23247 4709 23259 4743
rect 31726 4740 31754 4780
rect 47118 4768 47124 4780
rect 47176 4768 47182 4820
rect 23201 4703 23259 4709
rect 23308 4712 31754 4740
rect 22922 4672 22928 4684
rect 17276 4644 20944 4672
rect 21008 4644 22928 4672
rect 17276 4632 17282 4644
rect 18230 4564 18236 4616
rect 18288 4564 18294 4616
rect 21008 4613 21036 4644
rect 22922 4632 22928 4644
rect 22980 4632 22986 4684
rect 23106 4632 23112 4684
rect 23164 4672 23170 4684
rect 23308 4672 23336 4712
rect 47394 4700 47400 4752
rect 47452 4700 47458 4752
rect 23164 4644 23336 4672
rect 23164 4632 23170 4644
rect 25498 4632 25504 4684
rect 25556 4672 25562 4684
rect 25556 4644 47256 4672
rect 25556 4632 25562 4644
rect 20165 4607 20223 4613
rect 20165 4573 20177 4607
rect 20211 4604 20223 4607
rect 20257 4607 20315 4613
rect 20257 4604 20269 4607
rect 20211 4576 20269 4604
rect 20211 4573 20223 4576
rect 20165 4567 20223 4573
rect 20257 4573 20269 4576
rect 20303 4573 20315 4607
rect 20257 4567 20315 4573
rect 20993 4607 21051 4613
rect 20993 4573 21005 4607
rect 21039 4573 21051 4607
rect 20993 4567 21051 4573
rect 21453 4607 21511 4613
rect 21453 4573 21465 4607
rect 21499 4604 21511 4607
rect 23198 4604 23204 4616
rect 21499 4576 23204 4604
rect 21499 4573 21511 4576
rect 21453 4567 21511 4573
rect 23198 4564 23204 4576
rect 23256 4564 23262 4616
rect 23293 4607 23351 4613
rect 23293 4573 23305 4607
rect 23339 4604 23351 4607
rect 23385 4607 23443 4613
rect 23385 4604 23397 4607
rect 23339 4576 23397 4604
rect 23339 4573 23351 4576
rect 23293 4567 23351 4573
rect 23385 4573 23397 4576
rect 23431 4573 23443 4607
rect 23385 4567 23443 4573
rect 24949 4607 25007 4613
rect 24949 4573 24961 4607
rect 24995 4604 25007 4607
rect 25041 4607 25099 4613
rect 25041 4604 25053 4607
rect 24995 4576 25053 4604
rect 24995 4573 25007 4576
rect 24949 4567 25007 4573
rect 25041 4573 25053 4576
rect 25087 4573 25099 4607
rect 25041 4567 25099 4573
rect 40034 4564 40040 4616
rect 40092 4604 40098 4616
rect 47228 4613 47256 4644
rect 46845 4607 46903 4613
rect 46845 4604 46857 4607
rect 40092 4576 46857 4604
rect 40092 4564 40098 4576
rect 46845 4573 46857 4576
rect 46891 4573 46903 4607
rect 46845 4567 46903 4573
rect 47213 4607 47271 4613
rect 47213 4573 47225 4607
rect 47259 4573 47271 4607
rect 47213 4567 47271 4573
rect 8478 4496 8484 4548
rect 8536 4536 8542 4548
rect 47118 4536 47124 4548
rect 8536 4508 21312 4536
rect 8536 4496 8542 4508
rect 21284 4477 21312 4508
rect 23584 4508 47124 4536
rect 23584 4477 23612 4508
rect 47118 4496 47124 4508
rect 47176 4496 47182 4548
rect 21269 4471 21327 4477
rect 21269 4437 21281 4471
rect 21315 4437 21327 4471
rect 21269 4431 21327 4437
rect 23569 4471 23627 4477
rect 23569 4437 23581 4471
rect 23615 4437 23627 4471
rect 23569 4431 23627 4437
rect 24854 4428 24860 4480
rect 24912 4428 24918 4480
rect 25222 4428 25228 4480
rect 25280 4428 25286 4480
rect 47026 4428 47032 4480
rect 47084 4428 47090 4480
rect 1104 4378 47840 4400
rect 1104 4326 3010 4378
rect 3062 4326 3074 4378
rect 3126 4326 3138 4378
rect 3190 4326 3202 4378
rect 3254 4326 3266 4378
rect 3318 4326 9010 4378
rect 9062 4326 9074 4378
rect 9126 4326 9138 4378
rect 9190 4326 9202 4378
rect 9254 4326 9266 4378
rect 9318 4326 15010 4378
rect 15062 4326 15074 4378
rect 15126 4326 15138 4378
rect 15190 4326 15202 4378
rect 15254 4326 15266 4378
rect 15318 4326 21010 4378
rect 21062 4326 21074 4378
rect 21126 4326 21138 4378
rect 21190 4326 21202 4378
rect 21254 4326 21266 4378
rect 21318 4326 27010 4378
rect 27062 4326 27074 4378
rect 27126 4326 27138 4378
rect 27190 4326 27202 4378
rect 27254 4326 27266 4378
rect 27318 4326 33010 4378
rect 33062 4326 33074 4378
rect 33126 4326 33138 4378
rect 33190 4326 33202 4378
rect 33254 4326 33266 4378
rect 33318 4326 39010 4378
rect 39062 4326 39074 4378
rect 39126 4326 39138 4378
rect 39190 4326 39202 4378
rect 39254 4326 39266 4378
rect 39318 4326 45010 4378
rect 45062 4326 45074 4378
rect 45126 4326 45138 4378
rect 45190 4326 45202 4378
rect 45254 4326 45266 4378
rect 45318 4326 47840 4378
rect 1104 4304 47840 4326
rect 25222 4224 25228 4276
rect 25280 4264 25286 4276
rect 42702 4264 42708 4276
rect 25280 4236 42708 4264
rect 25280 4224 25286 4236
rect 42702 4224 42708 4236
rect 42760 4224 42766 4276
rect 16776 4168 16988 4196
rect 12713 4131 12771 4137
rect 12713 4097 12725 4131
rect 12759 4097 12771 4131
rect 12713 4091 12771 4097
rect 15841 4131 15899 4137
rect 15841 4097 15853 4131
rect 15887 4128 15899 4131
rect 16776 4128 16804 4168
rect 15887 4100 16804 4128
rect 16853 4131 16911 4137
rect 15887 4097 15899 4100
rect 15841 4091 15899 4097
rect 16853 4097 16865 4131
rect 16899 4097 16911 4131
rect 16960 4128 16988 4168
rect 17972 4168 18368 4196
rect 17972 4128 18000 4168
rect 16960 4100 18000 4128
rect 18049 4131 18107 4137
rect 16853 4091 16911 4097
rect 18049 4097 18061 4131
rect 18095 4128 18107 4131
rect 18233 4131 18291 4137
rect 18233 4128 18245 4131
rect 18095 4100 18245 4128
rect 18095 4097 18107 4100
rect 18049 4091 18107 4097
rect 18233 4097 18245 4100
rect 18279 4097 18291 4131
rect 18340 4128 18368 4168
rect 21450 4128 21456 4140
rect 18340 4100 21456 4128
rect 18233 4091 18291 4097
rect 12728 4060 12756 4091
rect 16868 4060 16896 4091
rect 21450 4088 21456 4100
rect 21508 4088 21514 4140
rect 22649 4131 22707 4137
rect 22649 4097 22661 4131
rect 22695 4128 22707 4131
rect 22741 4131 22799 4137
rect 22741 4128 22753 4131
rect 22695 4100 22753 4128
rect 22695 4097 22707 4100
rect 22649 4091 22707 4097
rect 22741 4097 22753 4100
rect 22787 4097 22799 4131
rect 46753 4131 46811 4137
rect 46753 4128 46765 4131
rect 22741 4091 22799 4097
rect 31726 4100 46765 4128
rect 21818 4060 21824 4072
rect 12728 4032 16804 4060
rect 16868 4032 21824 4060
rect 12986 3952 12992 4004
rect 13044 3992 13050 4004
rect 16669 3995 16727 4001
rect 16669 3992 16681 3995
rect 13044 3964 16681 3992
rect 13044 3952 13050 3964
rect 16669 3961 16681 3964
rect 16715 3961 16727 3995
rect 16669 3955 16727 3961
rect 2590 3884 2596 3936
rect 2648 3924 2654 3936
rect 12529 3927 12587 3933
rect 12529 3924 12541 3927
rect 2648 3896 12541 3924
rect 2648 3884 2654 3896
rect 12529 3893 12541 3896
rect 12575 3893 12587 3927
rect 12529 3887 12587 3893
rect 15657 3927 15715 3933
rect 15657 3893 15669 3927
rect 15703 3924 15715 3927
rect 15746 3924 15752 3936
rect 15703 3896 15752 3924
rect 15703 3893 15715 3896
rect 15657 3887 15715 3893
rect 15746 3884 15752 3896
rect 15804 3884 15810 3936
rect 16776 3924 16804 4032
rect 21818 4020 21824 4032
rect 21876 4020 21882 4072
rect 17954 3952 17960 4004
rect 18012 3952 18018 4004
rect 18417 3995 18475 4001
rect 18417 3961 18429 3995
rect 18463 3992 18475 3995
rect 31726 3992 31754 4100
rect 46753 4097 46765 4100
rect 46799 4097 46811 4131
rect 46753 4091 46811 4097
rect 47121 4131 47179 4137
rect 47121 4097 47133 4131
rect 47167 4097 47179 4131
rect 47121 4091 47179 4097
rect 44358 4020 44364 4072
rect 44416 4060 44422 4072
rect 47136 4060 47164 4091
rect 44416 4032 47164 4060
rect 44416 4020 44422 4032
rect 18463 3964 31754 3992
rect 18463 3961 18475 3964
rect 18417 3955 18475 3961
rect 47302 3952 47308 4004
rect 47360 3952 47366 4004
rect 19518 3924 19524 3936
rect 16776 3896 19524 3924
rect 19518 3884 19524 3896
rect 19576 3884 19582 3936
rect 20714 3884 20720 3936
rect 20772 3924 20778 3936
rect 22557 3927 22615 3933
rect 22557 3924 22569 3927
rect 20772 3896 22569 3924
rect 20772 3884 20778 3896
rect 22557 3893 22569 3896
rect 22603 3893 22615 3927
rect 22557 3887 22615 3893
rect 22925 3927 22983 3933
rect 22925 3893 22937 3927
rect 22971 3924 22983 3927
rect 25866 3924 25872 3936
rect 22971 3896 25872 3924
rect 22971 3893 22983 3896
rect 22925 3887 22983 3893
rect 25866 3884 25872 3896
rect 25924 3884 25930 3936
rect 37642 3884 37648 3936
rect 37700 3924 37706 3936
rect 46750 3924 46756 3936
rect 37700 3896 46756 3924
rect 37700 3884 37706 3896
rect 46750 3884 46756 3896
rect 46808 3884 46814 3936
rect 46934 3884 46940 3936
rect 46992 3884 46998 3936
rect 1104 3834 47840 3856
rect 1104 3782 1950 3834
rect 2002 3782 2014 3834
rect 2066 3782 2078 3834
rect 2130 3782 2142 3834
rect 2194 3782 2206 3834
rect 2258 3782 7950 3834
rect 8002 3782 8014 3834
rect 8066 3782 8078 3834
rect 8130 3782 8142 3834
rect 8194 3782 8206 3834
rect 8258 3782 13950 3834
rect 14002 3782 14014 3834
rect 14066 3782 14078 3834
rect 14130 3782 14142 3834
rect 14194 3782 14206 3834
rect 14258 3782 19950 3834
rect 20002 3782 20014 3834
rect 20066 3782 20078 3834
rect 20130 3782 20142 3834
rect 20194 3782 20206 3834
rect 20258 3782 25950 3834
rect 26002 3782 26014 3834
rect 26066 3782 26078 3834
rect 26130 3782 26142 3834
rect 26194 3782 26206 3834
rect 26258 3782 31950 3834
rect 32002 3782 32014 3834
rect 32066 3782 32078 3834
rect 32130 3782 32142 3834
rect 32194 3782 32206 3834
rect 32258 3782 37950 3834
rect 38002 3782 38014 3834
rect 38066 3782 38078 3834
rect 38130 3782 38142 3834
rect 38194 3782 38206 3834
rect 38258 3782 43950 3834
rect 44002 3782 44014 3834
rect 44066 3782 44078 3834
rect 44130 3782 44142 3834
rect 44194 3782 44206 3834
rect 44258 3782 47840 3834
rect 1104 3760 47840 3782
rect 24765 3723 24823 3729
rect 24765 3689 24777 3723
rect 24811 3720 24823 3723
rect 43346 3720 43352 3732
rect 24811 3692 43352 3720
rect 24811 3689 24823 3692
rect 24765 3683 24823 3689
rect 43346 3680 43352 3692
rect 43404 3680 43410 3732
rect 12802 3612 12808 3664
rect 12860 3652 12866 3664
rect 41782 3652 41788 3664
rect 12860 3624 41788 3652
rect 12860 3612 12866 3624
rect 41782 3612 41788 3624
rect 41840 3612 41846 3664
rect 47394 3612 47400 3664
rect 47452 3612 47458 3664
rect 8846 3544 8852 3596
rect 8904 3584 8910 3596
rect 8904 3556 24716 3584
rect 8904 3544 8910 3556
rect 14277 3519 14335 3525
rect 14277 3485 14289 3519
rect 14323 3516 14335 3519
rect 20165 3519 20223 3525
rect 14323 3488 20116 3516
rect 14323 3485 14335 3488
rect 14277 3479 14335 3485
rect 2314 3408 2320 3460
rect 2372 3448 2378 3460
rect 2372 3420 2774 3448
rect 2372 3408 2378 3420
rect 2746 3380 2774 3420
rect 6914 3408 6920 3460
rect 6972 3448 6978 3460
rect 6972 3420 20024 3448
rect 6972 3408 6978 3420
rect 19996 3389 20024 3420
rect 14093 3383 14151 3389
rect 14093 3380 14105 3383
rect 2746 3352 14105 3380
rect 14093 3349 14105 3352
rect 14139 3349 14151 3383
rect 14093 3343 14151 3349
rect 19981 3383 20039 3389
rect 19981 3349 19993 3383
rect 20027 3349 20039 3383
rect 20088 3380 20116 3488
rect 20165 3485 20177 3519
rect 20211 3485 20223 3519
rect 20165 3479 20223 3485
rect 20180 3448 20208 3479
rect 22094 3476 22100 3528
rect 22152 3516 22158 3528
rect 24581 3519 24639 3525
rect 24581 3516 24593 3519
rect 22152 3488 24593 3516
rect 22152 3476 22158 3488
rect 24581 3485 24593 3488
rect 24627 3485 24639 3519
rect 24688 3516 24716 3556
rect 24762 3544 24768 3596
rect 24820 3584 24826 3596
rect 24949 3587 25007 3593
rect 24949 3584 24961 3587
rect 24820 3556 24961 3584
rect 24820 3544 24826 3556
rect 24949 3553 24961 3556
rect 24995 3553 25007 3587
rect 29086 3584 29092 3596
rect 24949 3547 25007 3553
rect 25056 3556 29092 3584
rect 25056 3516 25084 3556
rect 29086 3544 29092 3556
rect 29144 3544 29150 3596
rect 42702 3544 42708 3596
rect 42760 3584 42766 3596
rect 42760 3556 47256 3584
rect 42760 3544 42766 3556
rect 24688 3488 25084 3516
rect 25133 3519 25191 3525
rect 24581 3479 24639 3485
rect 25133 3485 25145 3519
rect 25179 3485 25191 3519
rect 29454 3516 29460 3528
rect 25133 3479 25191 3485
rect 27356 3488 29460 3516
rect 22554 3448 22560 3460
rect 20180 3420 22560 3448
rect 22554 3408 22560 3420
rect 22612 3408 22618 3460
rect 25041 3451 25099 3457
rect 25041 3417 25053 3451
rect 25087 3448 25099 3451
rect 25148 3448 25176 3479
rect 27356 3448 27384 3488
rect 29454 3476 29460 3488
rect 29512 3476 29518 3528
rect 44174 3476 44180 3528
rect 44232 3516 44238 3528
rect 47228 3525 47256 3556
rect 46845 3519 46903 3525
rect 46845 3516 46857 3519
rect 44232 3488 46857 3516
rect 44232 3476 44238 3488
rect 46845 3485 46857 3488
rect 46891 3485 46903 3519
rect 46845 3479 46903 3485
rect 47213 3519 47271 3525
rect 47213 3485 47225 3519
rect 47259 3485 47271 3519
rect 47213 3479 47271 3485
rect 25087 3420 25176 3448
rect 25240 3420 27384 3448
rect 25087 3417 25099 3420
rect 25041 3411 25099 3417
rect 20898 3380 20904 3392
rect 20088 3352 20904 3380
rect 19981 3343 20039 3349
rect 20898 3340 20904 3352
rect 20956 3340 20962 3392
rect 23014 3340 23020 3392
rect 23072 3380 23078 3392
rect 25240 3380 25268 3420
rect 27430 3408 27436 3460
rect 27488 3448 27494 3460
rect 40770 3448 40776 3460
rect 27488 3420 40776 3448
rect 27488 3408 27494 3420
rect 40770 3408 40776 3420
rect 40828 3408 40834 3460
rect 23072 3352 25268 3380
rect 25317 3383 25375 3389
rect 23072 3340 23078 3352
rect 25317 3349 25329 3383
rect 25363 3380 25375 3383
rect 28534 3380 28540 3392
rect 25363 3352 28540 3380
rect 25363 3349 25375 3352
rect 25317 3343 25375 3349
rect 28534 3340 28540 3352
rect 28592 3340 28598 3392
rect 33594 3340 33600 3392
rect 33652 3380 33658 3392
rect 43806 3380 43812 3392
rect 33652 3352 43812 3380
rect 33652 3340 33658 3352
rect 43806 3340 43812 3352
rect 43864 3340 43870 3392
rect 47026 3340 47032 3392
rect 47084 3340 47090 3392
rect 1104 3290 47840 3312
rect 1104 3238 3010 3290
rect 3062 3238 3074 3290
rect 3126 3238 3138 3290
rect 3190 3238 3202 3290
rect 3254 3238 3266 3290
rect 3318 3238 9010 3290
rect 9062 3238 9074 3290
rect 9126 3238 9138 3290
rect 9190 3238 9202 3290
rect 9254 3238 9266 3290
rect 9318 3238 15010 3290
rect 15062 3238 15074 3290
rect 15126 3238 15138 3290
rect 15190 3238 15202 3290
rect 15254 3238 15266 3290
rect 15318 3238 21010 3290
rect 21062 3238 21074 3290
rect 21126 3238 21138 3290
rect 21190 3238 21202 3290
rect 21254 3238 21266 3290
rect 21318 3238 27010 3290
rect 27062 3238 27074 3290
rect 27126 3238 27138 3290
rect 27190 3238 27202 3290
rect 27254 3238 27266 3290
rect 27318 3238 33010 3290
rect 33062 3238 33074 3290
rect 33126 3238 33138 3290
rect 33190 3238 33202 3290
rect 33254 3238 33266 3290
rect 33318 3238 39010 3290
rect 39062 3238 39074 3290
rect 39126 3238 39138 3290
rect 39190 3238 39202 3290
rect 39254 3238 39266 3290
rect 39318 3238 45010 3290
rect 45062 3238 45074 3290
rect 45126 3238 45138 3290
rect 45190 3238 45202 3290
rect 45254 3238 45266 3290
rect 45318 3238 47840 3290
rect 1104 3216 47840 3238
rect 8846 3136 8852 3188
rect 8904 3136 8910 3188
rect 12802 3136 12808 3188
rect 12860 3136 12866 3188
rect 13538 3136 13544 3188
rect 13596 3176 13602 3188
rect 17681 3179 17739 3185
rect 17681 3176 17693 3179
rect 13596 3148 17693 3176
rect 13596 3136 13602 3148
rect 17681 3145 17693 3148
rect 17727 3145 17739 3179
rect 17681 3139 17739 3145
rect 22097 3179 22155 3185
rect 22097 3145 22109 3179
rect 22143 3176 22155 3179
rect 23014 3176 23020 3188
rect 22143 3148 23020 3176
rect 22143 3145 22155 3148
rect 22097 3139 22155 3145
rect 23014 3136 23020 3148
rect 23072 3136 23078 3188
rect 23106 3136 23112 3188
rect 23164 3136 23170 3188
rect 26694 3136 26700 3188
rect 26752 3176 26758 3188
rect 26752 3148 29316 3176
rect 26752 3136 26758 3148
rect 8294 3068 8300 3120
rect 8352 3108 8358 3120
rect 8757 3111 8815 3117
rect 8757 3108 8769 3111
rect 8352 3080 8769 3108
rect 8352 3068 8358 3080
rect 8757 3077 8769 3080
rect 8803 3077 8815 3111
rect 8757 3071 8815 3077
rect 9582 3068 9588 3120
rect 9640 3108 9646 3120
rect 13081 3111 13139 3117
rect 13081 3108 13093 3111
rect 9640 3080 13093 3108
rect 9640 3068 9646 3080
rect 13081 3077 13093 3080
rect 13127 3077 13139 3111
rect 13081 3071 13139 3077
rect 17773 3111 17831 3117
rect 17773 3077 17785 3111
rect 17819 3108 17831 3111
rect 17957 3111 18015 3117
rect 17957 3108 17969 3111
rect 17819 3080 17969 3108
rect 17819 3077 17831 3080
rect 17773 3071 17831 3077
rect 17957 3077 17969 3080
rect 18003 3077 18015 3111
rect 17957 3071 18015 3077
rect 18138 3068 18144 3120
rect 18196 3068 18202 3120
rect 19794 3068 19800 3120
rect 19852 3108 19858 3120
rect 19852 3080 21956 3108
rect 19852 3068 19858 3080
rect 8205 3043 8263 3049
rect 8205 3009 8217 3043
rect 8251 3040 8263 3043
rect 8389 3043 8447 3049
rect 8389 3040 8401 3043
rect 8251 3012 8401 3040
rect 8251 3009 8263 3012
rect 8205 3003 8263 3009
rect 8389 3009 8401 3012
rect 8435 3009 8447 3043
rect 8389 3003 8447 3009
rect 10594 3000 10600 3052
rect 10652 3040 10658 3052
rect 10873 3043 10931 3049
rect 10873 3040 10885 3043
rect 10652 3012 10885 3040
rect 10652 3000 10658 3012
rect 10873 3009 10885 3012
rect 10919 3009 10931 3043
rect 10873 3003 10931 3009
rect 12713 3043 12771 3049
rect 12713 3009 12725 3043
rect 12759 3040 12771 3043
rect 12894 3040 12900 3052
rect 12759 3012 12900 3040
rect 12759 3009 12771 3012
rect 12713 3003 12771 3009
rect 12894 3000 12900 3012
rect 12952 3000 12958 3052
rect 15378 3000 15384 3052
rect 15436 3040 15442 3052
rect 21928 3049 21956 3080
rect 22066 3080 23796 3108
rect 15749 3043 15807 3049
rect 15749 3040 15761 3043
rect 15436 3012 15761 3040
rect 15436 3000 15442 3012
rect 15749 3009 15761 3012
rect 15795 3009 15807 3043
rect 15749 3003 15807 3009
rect 16761 3043 16819 3049
rect 16761 3009 16773 3043
rect 16807 3009 16819 3043
rect 16761 3003 16819 3009
rect 18693 3043 18751 3049
rect 18693 3009 18705 3043
rect 18739 3009 18751 3043
rect 18693 3003 18751 3009
rect 20165 3043 20223 3049
rect 20165 3009 20177 3043
rect 20211 3040 20223 3043
rect 20257 3043 20315 3049
rect 20257 3040 20269 3043
rect 20211 3012 20269 3040
rect 20211 3009 20223 3012
rect 20165 3003 20223 3009
rect 20257 3009 20269 3012
rect 20303 3009 20315 3043
rect 20257 3003 20315 3009
rect 20809 3043 20867 3049
rect 20809 3009 20821 3043
rect 20855 3040 20867 3043
rect 20901 3043 20959 3049
rect 20901 3040 20913 3043
rect 20855 3012 20913 3040
rect 20855 3009 20867 3012
rect 20809 3003 20867 3009
rect 20901 3009 20913 3012
rect 20947 3009 20959 3043
rect 20901 3003 20959 3009
rect 21913 3043 21971 3049
rect 21913 3009 21925 3043
rect 21959 3009 21971 3043
rect 21913 3003 21971 3009
rect 11054 2932 11060 2984
rect 11112 2932 11118 2984
rect 16776 2972 16804 3003
rect 12406 2944 16804 2972
rect 8570 2864 8576 2916
rect 8628 2864 8634 2916
rect 9490 2864 9496 2916
rect 9548 2904 9554 2916
rect 12406 2904 12434 2944
rect 17494 2932 17500 2984
rect 17552 2972 17558 2984
rect 18708 2972 18736 3003
rect 22066 2972 22094 3080
rect 22738 3000 22744 3052
rect 22796 3040 22802 3052
rect 22925 3043 22983 3049
rect 22925 3040 22937 3043
rect 22796 3012 22937 3040
rect 22796 3000 22802 3012
rect 22925 3009 22937 3012
rect 22971 3009 22983 3043
rect 22925 3003 22983 3009
rect 23768 2972 23796 3080
rect 24394 3068 24400 3120
rect 24452 3108 24458 3120
rect 24452 3080 27292 3108
rect 24452 3068 24458 3080
rect 25314 3000 25320 3052
rect 25372 3000 25378 3052
rect 27264 3049 27292 3080
rect 27249 3043 27307 3049
rect 27249 3009 27261 3043
rect 27295 3009 27307 3043
rect 27249 3003 27307 3009
rect 27522 3000 27528 3052
rect 27580 3000 27586 3052
rect 29288 3049 29316 3148
rect 29362 3136 29368 3188
rect 29420 3176 29426 3188
rect 29420 3148 31984 3176
rect 29420 3136 29426 3148
rect 29273 3043 29331 3049
rect 29273 3009 29285 3043
rect 29319 3009 29331 3043
rect 29273 3003 29331 3009
rect 29454 3000 29460 3052
rect 29512 3040 29518 3052
rect 31956 3040 31984 3148
rect 32030 3136 32036 3188
rect 32088 3176 32094 3188
rect 37734 3176 37740 3188
rect 32088 3148 37740 3176
rect 32088 3136 32094 3148
rect 37734 3136 37740 3148
rect 37792 3136 37798 3188
rect 38746 3136 38752 3188
rect 38804 3136 38810 3188
rect 39666 3136 39672 3188
rect 39724 3136 39730 3188
rect 40497 3179 40555 3185
rect 40497 3145 40509 3179
rect 40543 3176 40555 3179
rect 40678 3176 40684 3188
rect 40543 3148 40684 3176
rect 40543 3145 40555 3148
rect 40497 3139 40555 3145
rect 40678 3136 40684 3148
rect 40736 3136 40742 3188
rect 43254 3136 43260 3188
rect 43312 3136 43318 3188
rect 43898 3136 43904 3188
rect 43956 3176 43962 3188
rect 43993 3179 44051 3185
rect 43993 3176 44005 3179
rect 43956 3148 44005 3176
rect 43956 3136 43962 3148
rect 43993 3145 44005 3148
rect 44039 3145 44051 3179
rect 43993 3139 44051 3145
rect 47302 3136 47308 3188
rect 47360 3136 47366 3188
rect 44450 3108 44456 3120
rect 32140 3080 44456 3108
rect 32140 3040 32168 3080
rect 44450 3068 44456 3080
rect 44508 3068 44514 3120
rect 29512 3012 31892 3040
rect 31956 3012 32168 3040
rect 29512 3000 29518 3012
rect 31754 2972 31760 2984
rect 17552 2944 18736 2972
rect 18892 2944 22094 2972
rect 23032 2944 23244 2972
rect 23768 2944 31760 2972
rect 17552 2932 17558 2944
rect 9548 2876 12434 2904
rect 9548 2864 9554 2876
rect 13262 2864 13268 2916
rect 13320 2864 13326 2916
rect 18892 2913 18920 2944
rect 15933 2907 15991 2913
rect 15933 2873 15945 2907
rect 15979 2904 15991 2907
rect 18877 2907 18935 2913
rect 15979 2876 18828 2904
rect 15979 2873 15991 2876
rect 15933 2867 15991 2873
rect 1302 2796 1308 2848
rect 1360 2836 1366 2848
rect 8113 2839 8171 2845
rect 8113 2836 8125 2839
rect 1360 2808 8125 2836
rect 1360 2796 1366 2808
rect 8113 2805 8125 2808
rect 8159 2805 8171 2839
rect 8113 2799 8171 2805
rect 16850 2796 16856 2848
rect 16908 2796 16914 2848
rect 18800 2836 18828 2876
rect 18877 2873 18889 2907
rect 18923 2873 18935 2907
rect 23032 2904 23060 2944
rect 18877 2867 18935 2873
rect 18984 2876 23060 2904
rect 23216 2904 23244 2944
rect 31754 2932 31760 2944
rect 31812 2932 31818 2984
rect 31864 2972 31892 3012
rect 36446 3000 36452 3052
rect 36504 3040 36510 3052
rect 36541 3043 36599 3049
rect 36541 3040 36553 3043
rect 36504 3012 36553 3040
rect 36504 3000 36510 3012
rect 36541 3009 36553 3012
rect 36587 3040 36599 3043
rect 36725 3043 36783 3049
rect 36725 3040 36737 3043
rect 36587 3012 36737 3040
rect 36587 3009 36599 3012
rect 36541 3003 36599 3009
rect 36725 3009 36737 3012
rect 36771 3009 36783 3043
rect 36725 3003 36783 3009
rect 37274 3000 37280 3052
rect 37332 3040 37338 3052
rect 37461 3043 37519 3049
rect 37461 3040 37473 3043
rect 37332 3012 37473 3040
rect 37332 3000 37338 3012
rect 37461 3009 37473 3012
rect 37507 3009 37519 3043
rect 37461 3003 37519 3009
rect 38562 3000 38568 3052
rect 38620 3000 38626 3052
rect 39482 3000 39488 3052
rect 39540 3000 39546 3052
rect 40310 3000 40316 3052
rect 40368 3000 40374 3052
rect 43070 3000 43076 3052
rect 43128 3000 43134 3052
rect 43806 3000 43812 3052
rect 43864 3000 43870 3052
rect 46750 3000 46756 3052
rect 46808 3000 46814 3052
rect 47118 3000 47124 3052
rect 47176 3000 47182 3052
rect 42242 2972 42248 2984
rect 31864 2944 42248 2972
rect 42242 2932 42248 2944
rect 42300 2932 42306 2984
rect 41874 2904 41880 2916
rect 23216 2876 41880 2904
rect 18984 2836 19012 2876
rect 41874 2864 41880 2876
rect 41932 2864 41938 2916
rect 18800 2808 19012 2836
rect 19702 2796 19708 2848
rect 19760 2836 19766 2848
rect 20073 2839 20131 2845
rect 20073 2836 20085 2839
rect 19760 2808 20085 2836
rect 19760 2796 19766 2808
rect 20073 2805 20085 2808
rect 20119 2805 20131 2839
rect 20073 2799 20131 2805
rect 20438 2796 20444 2848
rect 20496 2796 20502 2848
rect 20714 2796 20720 2848
rect 20772 2796 20778 2848
rect 21082 2796 21088 2848
rect 21140 2796 21146 2848
rect 25501 2839 25559 2845
rect 25501 2805 25513 2839
rect 25547 2836 25559 2839
rect 26510 2836 26516 2848
rect 25547 2808 26516 2836
rect 25547 2805 25559 2808
rect 25501 2799 25559 2805
rect 26510 2796 26516 2808
rect 26568 2796 26574 2848
rect 27430 2796 27436 2848
rect 27488 2796 27494 2848
rect 27709 2839 27767 2845
rect 27709 2805 27721 2839
rect 27755 2836 27767 2839
rect 29362 2836 29368 2848
rect 27755 2808 29368 2836
rect 27755 2805 27767 2808
rect 27709 2799 27767 2805
rect 29362 2796 29368 2808
rect 29420 2796 29426 2848
rect 29457 2839 29515 2845
rect 29457 2805 29469 2839
rect 29503 2836 29515 2839
rect 35802 2836 35808 2848
rect 29503 2808 35808 2836
rect 29503 2805 29515 2808
rect 29457 2799 29515 2805
rect 35802 2796 35808 2808
rect 35860 2796 35866 2848
rect 36906 2796 36912 2848
rect 36964 2796 36970 2848
rect 37642 2796 37648 2848
rect 37700 2796 37706 2848
rect 37734 2796 37740 2848
rect 37792 2836 37798 2848
rect 42978 2836 42984 2848
rect 37792 2808 42984 2836
rect 37792 2796 37798 2808
rect 42978 2796 42984 2808
rect 43036 2796 43042 2848
rect 46934 2796 46940 2848
rect 46992 2796 46998 2848
rect 1104 2746 47840 2768
rect 1104 2694 1950 2746
rect 2002 2694 2014 2746
rect 2066 2694 2078 2746
rect 2130 2694 2142 2746
rect 2194 2694 2206 2746
rect 2258 2694 7950 2746
rect 8002 2694 8014 2746
rect 8066 2694 8078 2746
rect 8130 2694 8142 2746
rect 8194 2694 8206 2746
rect 8258 2694 13950 2746
rect 14002 2694 14014 2746
rect 14066 2694 14078 2746
rect 14130 2694 14142 2746
rect 14194 2694 14206 2746
rect 14258 2694 19950 2746
rect 20002 2694 20014 2746
rect 20066 2694 20078 2746
rect 20130 2694 20142 2746
rect 20194 2694 20206 2746
rect 20258 2694 25950 2746
rect 26002 2694 26014 2746
rect 26066 2694 26078 2746
rect 26130 2694 26142 2746
rect 26194 2694 26206 2746
rect 26258 2694 31950 2746
rect 32002 2694 32014 2746
rect 32066 2694 32078 2746
rect 32130 2694 32142 2746
rect 32194 2694 32206 2746
rect 32258 2694 37950 2746
rect 38002 2694 38014 2746
rect 38066 2694 38078 2746
rect 38130 2694 38142 2746
rect 38194 2694 38206 2746
rect 38258 2694 43950 2746
rect 44002 2694 44014 2746
rect 44066 2694 44078 2746
rect 44130 2694 44142 2746
rect 44194 2694 44206 2746
rect 44258 2694 47840 2746
rect 1104 2672 47840 2694
rect 20438 2592 20444 2644
rect 20496 2632 20502 2644
rect 42150 2632 42156 2644
rect 20496 2604 42156 2632
rect 20496 2592 20502 2604
rect 42150 2592 42156 2604
rect 42208 2592 42214 2644
rect 42904 2604 43208 2632
rect 16850 2524 16856 2576
rect 16908 2564 16914 2576
rect 42904 2564 42932 2604
rect 16908 2536 42932 2564
rect 43180 2564 43208 2604
rect 45830 2592 45836 2644
rect 45888 2592 45894 2644
rect 43180 2536 47164 2564
rect 16908 2524 16914 2536
rect 13262 2456 13268 2508
rect 13320 2496 13326 2508
rect 33134 2496 33140 2508
rect 13320 2468 33140 2496
rect 13320 2456 13326 2468
rect 33134 2456 33140 2468
rect 33192 2456 33198 2508
rect 43180 2468 46428 2496
rect 8570 2388 8576 2440
rect 8628 2428 8634 2440
rect 36262 2428 36268 2440
rect 8628 2400 36268 2428
rect 8628 2388 8634 2400
rect 36262 2388 36268 2400
rect 36320 2388 36326 2440
rect 36446 2388 36452 2440
rect 36504 2428 36510 2440
rect 43180 2428 43208 2468
rect 36504 2400 43208 2428
rect 36504 2388 36510 2400
rect 45646 2388 45652 2440
rect 45704 2388 45710 2440
rect 46400 2437 46428 2468
rect 47136 2437 47164 2536
rect 47302 2524 47308 2576
rect 47360 2524 47366 2576
rect 46017 2431 46075 2437
rect 46017 2397 46029 2431
rect 46063 2397 46075 2431
rect 46017 2391 46075 2397
rect 46385 2431 46443 2437
rect 46385 2397 46397 2431
rect 46431 2397 46443 2431
rect 46385 2391 46443 2397
rect 46753 2431 46811 2437
rect 46753 2397 46765 2431
rect 46799 2397 46811 2431
rect 46753 2391 46811 2397
rect 47121 2431 47179 2437
rect 47121 2397 47133 2431
rect 47167 2397 47179 2431
rect 47121 2391 47179 2397
rect 21082 2320 21088 2372
rect 21140 2360 21146 2372
rect 21140 2332 31754 2360
rect 21140 2320 21146 2332
rect 5626 2252 5632 2304
rect 5684 2292 5690 2304
rect 27522 2292 27528 2304
rect 5684 2264 27528 2292
rect 5684 2252 5690 2264
rect 27522 2252 27528 2264
rect 27580 2252 27586 2304
rect 31726 2292 31754 2332
rect 33134 2320 33140 2372
rect 33192 2360 33198 2372
rect 46032 2360 46060 2391
rect 46768 2360 46796 2391
rect 33192 2332 46060 2360
rect 46124 2332 46796 2360
rect 33192 2320 33198 2332
rect 46124 2292 46152 2332
rect 31726 2264 46152 2292
rect 46198 2252 46204 2304
rect 46256 2252 46262 2304
rect 46566 2252 46572 2304
rect 46624 2252 46630 2304
rect 46934 2252 46940 2304
rect 46992 2252 46998 2304
rect 1104 2202 47840 2224
rect 1104 2150 3010 2202
rect 3062 2150 3074 2202
rect 3126 2150 3138 2202
rect 3190 2150 3202 2202
rect 3254 2150 3266 2202
rect 3318 2150 9010 2202
rect 9062 2150 9074 2202
rect 9126 2150 9138 2202
rect 9190 2150 9202 2202
rect 9254 2150 9266 2202
rect 9318 2150 15010 2202
rect 15062 2150 15074 2202
rect 15126 2150 15138 2202
rect 15190 2150 15202 2202
rect 15254 2150 15266 2202
rect 15318 2150 21010 2202
rect 21062 2150 21074 2202
rect 21126 2150 21138 2202
rect 21190 2150 21202 2202
rect 21254 2150 21266 2202
rect 21318 2150 27010 2202
rect 27062 2150 27074 2202
rect 27126 2150 27138 2202
rect 27190 2150 27202 2202
rect 27254 2150 27266 2202
rect 27318 2150 33010 2202
rect 33062 2150 33074 2202
rect 33126 2150 33138 2202
rect 33190 2150 33202 2202
rect 33254 2150 33266 2202
rect 33318 2150 39010 2202
rect 39062 2150 39074 2202
rect 39126 2150 39138 2202
rect 39190 2150 39202 2202
rect 39254 2150 39266 2202
rect 39318 2150 45010 2202
rect 45062 2150 45074 2202
rect 45126 2150 45138 2202
rect 45190 2150 45202 2202
rect 45254 2150 45266 2202
rect 45318 2150 47840 2202
rect 1104 2128 47840 2150
rect 2866 2048 2872 2100
rect 2924 2088 2930 2100
rect 25314 2088 25320 2100
rect 2924 2060 25320 2088
rect 2924 2048 2930 2060
rect 25314 2048 25320 2060
rect 25372 2048 25378 2100
rect 31294 2048 31300 2100
rect 31352 2088 31358 2100
rect 43070 2088 43076 2100
rect 31352 2060 43076 2088
rect 31352 2048 31358 2060
rect 43070 2048 43076 2060
rect 43128 2048 43134 2100
rect 3694 144 3700 196
rect 3752 144 3758 196
rect 5994 144 6000 196
rect 6052 184 6058 196
rect 40310 184 40316 196
rect 6052 156 40316 184
rect 6052 144 6058 156
rect 40310 144 40316 156
rect 40368 144 40374 196
rect 3712 116 3740 144
rect 39482 116 39488 128
rect 3712 88 39488 116
rect 39482 76 39488 88
rect 39540 76 39546 128
rect 1486 8 1492 60
rect 1544 48 1550 60
rect 38562 48 38568 60
rect 1544 20 38568 48
rect 1544 8 1550 20
rect 38562 8 38568 20
rect 38620 8 38626 60
<< via1 >>
rect 13544 11160 13596 11212
rect 39488 11160 39540 11212
rect 14924 11092 14976 11144
rect 38752 11092 38804 11144
rect 18236 11024 18288 11076
rect 36544 11024 36596 11076
rect 11796 10956 11848 11008
rect 29184 10956 29236 11008
rect 18328 10888 18380 10940
rect 36176 10888 36228 10940
rect 21916 10684 21968 10736
rect 24032 10684 24084 10736
rect 1308 9324 1360 9376
rect 7656 9324 7708 9376
rect 8760 9324 8812 9376
rect 16856 9324 16908 9376
rect 4344 9256 4396 9308
rect 20260 9324 20312 9376
rect 6276 9188 6328 9240
rect 25780 9256 25832 9308
rect 19156 9188 19208 9240
rect 26792 9188 26844 9240
rect 3516 8984 3568 9036
rect 23388 9120 23440 9172
rect 34428 9120 34480 9172
rect 45560 9120 45612 9172
rect 7012 9052 7064 9104
rect 15476 9052 15528 9104
rect 15660 9052 15712 9104
rect 38384 9052 38436 9104
rect 4712 8916 4764 8968
rect 8484 8984 8536 9036
rect 14556 8984 14608 9036
rect 39120 8984 39172 9036
rect 7656 8916 7708 8968
rect 6184 8848 6236 8900
rect 14648 8848 14700 8900
rect 15476 8848 15528 8900
rect 15752 8848 15804 8900
rect 26792 8916 26844 8968
rect 36912 8916 36964 8968
rect 42892 8916 42944 8968
rect 46572 8916 46624 8968
rect 32404 8848 32456 8900
rect 43260 8848 43312 8900
rect 45468 8848 45520 8900
rect 5080 8780 5132 8832
rect 8668 8780 8720 8832
rect 10232 8780 10284 8832
rect 18972 8780 19024 8832
rect 19708 8780 19760 8832
rect 40500 8780 40552 8832
rect 40776 8780 40828 8832
rect 43720 8780 43772 8832
rect 45376 8780 45428 8832
rect 46388 8780 46440 8832
rect 3010 8678 3062 8730
rect 3074 8678 3126 8730
rect 3138 8678 3190 8730
rect 3202 8678 3254 8730
rect 3266 8678 3318 8730
rect 9010 8678 9062 8730
rect 9074 8678 9126 8730
rect 9138 8678 9190 8730
rect 9202 8678 9254 8730
rect 9266 8678 9318 8730
rect 15010 8678 15062 8730
rect 15074 8678 15126 8730
rect 15138 8678 15190 8730
rect 15202 8678 15254 8730
rect 15266 8678 15318 8730
rect 21010 8678 21062 8730
rect 21074 8678 21126 8730
rect 21138 8678 21190 8730
rect 21202 8678 21254 8730
rect 21266 8678 21318 8730
rect 27010 8678 27062 8730
rect 27074 8678 27126 8730
rect 27138 8678 27190 8730
rect 27202 8678 27254 8730
rect 27266 8678 27318 8730
rect 33010 8678 33062 8730
rect 33074 8678 33126 8730
rect 33138 8678 33190 8730
rect 33202 8678 33254 8730
rect 33266 8678 33318 8730
rect 39010 8678 39062 8730
rect 39074 8678 39126 8730
rect 39138 8678 39190 8730
rect 39202 8678 39254 8730
rect 39266 8678 39318 8730
rect 45010 8678 45062 8730
rect 45074 8678 45126 8730
rect 45138 8678 45190 8730
rect 45202 8678 45254 8730
rect 45266 8678 45318 8730
rect 1952 8576 2004 8628
rect 2320 8576 2372 8628
rect 2688 8576 2740 8628
rect 2872 8576 2924 8628
rect 3424 8619 3476 8628
rect 3424 8585 3433 8619
rect 3433 8585 3467 8619
rect 3467 8585 3476 8619
rect 3424 8576 3476 8585
rect 4160 8619 4212 8628
rect 4160 8585 4169 8619
rect 4169 8585 4203 8619
rect 4203 8585 4212 8619
rect 4160 8576 4212 8585
rect 4528 8619 4580 8628
rect 4528 8585 4537 8619
rect 4537 8585 4571 8619
rect 4571 8585 4580 8619
rect 4528 8576 4580 8585
rect 4896 8619 4948 8628
rect 4896 8585 4905 8619
rect 4905 8585 4939 8619
rect 4939 8585 4948 8619
rect 4896 8576 4948 8585
rect 5264 8619 5316 8628
rect 5264 8585 5273 8619
rect 5273 8585 5307 8619
rect 5307 8585 5316 8619
rect 5264 8576 5316 8585
rect 5632 8619 5684 8628
rect 5632 8585 5641 8619
rect 5641 8585 5675 8619
rect 5675 8585 5684 8619
rect 5632 8576 5684 8585
rect 6000 8619 6052 8628
rect 6000 8585 6009 8619
rect 6009 8585 6043 8619
rect 6043 8585 6052 8619
rect 6000 8576 6052 8585
rect 2320 8483 2372 8492
rect 2320 8449 2329 8483
rect 2329 8449 2363 8483
rect 2363 8449 2372 8483
rect 2320 8440 2372 8449
rect 2596 8440 2648 8492
rect 3516 8440 3568 8492
rect 4344 8483 4396 8492
rect 4344 8449 4353 8483
rect 4353 8449 4387 8483
rect 4387 8449 4396 8483
rect 4344 8440 4396 8449
rect 4712 8483 4764 8492
rect 4712 8449 4721 8483
rect 4721 8449 4755 8483
rect 4755 8449 4764 8483
rect 4712 8440 4764 8449
rect 5080 8483 5132 8492
rect 5080 8449 5089 8483
rect 5089 8449 5123 8483
rect 5123 8449 5132 8483
rect 5080 8440 5132 8449
rect 6184 8576 6236 8628
rect 6736 8619 6788 8628
rect 6736 8585 6745 8619
rect 6745 8585 6779 8619
rect 6779 8585 6788 8619
rect 6736 8576 6788 8585
rect 7104 8619 7156 8628
rect 7104 8585 7113 8619
rect 7113 8585 7147 8619
rect 7147 8585 7156 8619
rect 7104 8576 7156 8585
rect 7472 8619 7524 8628
rect 7472 8585 7481 8619
rect 7481 8585 7515 8619
rect 7515 8585 7524 8619
rect 7472 8576 7524 8585
rect 7840 8619 7892 8628
rect 7840 8585 7849 8619
rect 7849 8585 7883 8619
rect 7883 8585 7892 8619
rect 7840 8576 7892 8585
rect 8208 8619 8260 8628
rect 8208 8585 8217 8619
rect 8217 8585 8251 8619
rect 8251 8585 8260 8619
rect 8208 8576 8260 8585
rect 8576 8619 8628 8628
rect 8576 8585 8585 8619
rect 8585 8585 8619 8619
rect 8619 8585 8628 8619
rect 8576 8576 8628 8585
rect 9404 8576 9456 8628
rect 9680 8619 9732 8628
rect 9680 8585 9689 8619
rect 9689 8585 9723 8619
rect 9723 8585 9732 8619
rect 9680 8576 9732 8585
rect 10048 8619 10100 8628
rect 10048 8585 10057 8619
rect 10057 8585 10091 8619
rect 10091 8585 10100 8619
rect 10048 8576 10100 8585
rect 10416 8619 10468 8628
rect 10416 8585 10425 8619
rect 10425 8585 10459 8619
rect 10459 8585 10468 8619
rect 10416 8576 10468 8585
rect 10784 8619 10836 8628
rect 10784 8585 10793 8619
rect 10793 8585 10827 8619
rect 10827 8585 10836 8619
rect 10784 8576 10836 8585
rect 11152 8619 11204 8628
rect 11152 8585 11161 8619
rect 11161 8585 11195 8619
rect 11195 8585 11204 8619
rect 11152 8576 11204 8585
rect 11888 8619 11940 8628
rect 11888 8585 11897 8619
rect 11897 8585 11931 8619
rect 11931 8585 11940 8619
rect 11888 8576 11940 8585
rect 12256 8619 12308 8628
rect 12256 8585 12265 8619
rect 12265 8585 12299 8619
rect 12299 8585 12308 8619
rect 12256 8576 12308 8585
rect 12624 8619 12676 8628
rect 12624 8585 12633 8619
rect 12633 8585 12667 8619
rect 12667 8585 12676 8619
rect 12624 8576 12676 8585
rect 12992 8619 13044 8628
rect 12992 8585 13001 8619
rect 13001 8585 13035 8619
rect 13035 8585 13044 8619
rect 12992 8576 13044 8585
rect 13360 8576 13412 8628
rect 13728 8576 13780 8628
rect 14464 8576 14516 8628
rect 14832 8576 14884 8628
rect 15384 8576 15436 8628
rect 15568 8576 15620 8628
rect 15936 8576 15988 8628
rect 16304 8576 16356 8628
rect 17408 8576 17460 8628
rect 18052 8576 18104 8628
rect 18512 8576 18564 8628
rect 19248 8576 19300 8628
rect 19616 8619 19668 8628
rect 19616 8585 19625 8619
rect 19625 8585 19659 8619
rect 19659 8585 19668 8619
rect 19616 8576 19668 8585
rect 19708 8576 19760 8628
rect 19984 8576 20036 8628
rect 20352 8576 20404 8628
rect 39856 8576 39908 8628
rect 40224 8576 40276 8628
rect 40592 8576 40644 8628
rect 40960 8576 41012 8628
rect 41328 8576 41380 8628
rect 41696 8576 41748 8628
rect 42064 8576 42116 8628
rect 42800 8576 42852 8628
rect 43904 8576 43956 8628
rect 44640 8576 44692 8628
rect 6276 8440 6328 8492
rect 6828 8440 6880 8492
rect 6828 8304 6880 8356
rect 7656 8483 7708 8492
rect 7656 8449 7665 8483
rect 7665 8449 7699 8483
rect 7699 8449 7708 8483
rect 7656 8440 7708 8449
rect 7840 8440 7892 8492
rect 8392 8483 8444 8492
rect 8392 8449 8401 8483
rect 8401 8449 8435 8483
rect 8435 8449 8444 8483
rect 8392 8440 8444 8449
rect 8760 8483 8812 8492
rect 8760 8449 8769 8483
rect 8769 8449 8803 8483
rect 8803 8449 8812 8483
rect 8760 8440 8812 8449
rect 9496 8483 9548 8492
rect 9496 8449 9505 8483
rect 9505 8449 9539 8483
rect 9539 8449 9548 8483
rect 9496 8440 9548 8449
rect 9864 8483 9916 8492
rect 9864 8449 9873 8483
rect 9873 8449 9907 8483
rect 9907 8449 9916 8483
rect 9864 8440 9916 8449
rect 10232 8483 10284 8492
rect 10232 8449 10241 8483
rect 10241 8449 10275 8483
rect 10275 8449 10284 8483
rect 10232 8440 10284 8449
rect 11244 8508 11296 8560
rect 11428 8508 11480 8560
rect 10968 8483 11020 8492
rect 10968 8449 10977 8483
rect 10977 8449 11011 8483
rect 11011 8449 11020 8483
rect 10968 8440 11020 8449
rect 11152 8304 11204 8356
rect 7012 8236 7064 8288
rect 12716 8440 12768 8492
rect 12624 8372 12676 8424
rect 13176 8483 13228 8492
rect 13176 8449 13185 8483
rect 13185 8449 13219 8483
rect 13219 8449 13228 8483
rect 13176 8440 13228 8449
rect 14648 8508 14700 8560
rect 13636 8483 13688 8492
rect 13636 8449 13645 8483
rect 13645 8449 13679 8483
rect 13679 8449 13688 8483
rect 13636 8440 13688 8449
rect 13728 8440 13780 8492
rect 14464 8440 14516 8492
rect 15108 8483 15160 8492
rect 15108 8449 15117 8483
rect 15117 8449 15151 8483
rect 15151 8449 15160 8483
rect 15108 8440 15160 8449
rect 15476 8483 15528 8492
rect 15476 8449 15485 8483
rect 15485 8449 15519 8483
rect 15519 8449 15528 8483
rect 15476 8440 15528 8449
rect 15844 8483 15896 8492
rect 15844 8449 15853 8483
rect 15853 8449 15887 8483
rect 15887 8449 15896 8483
rect 15844 8440 15896 8449
rect 16212 8483 16264 8492
rect 16212 8449 16221 8483
rect 16221 8449 16255 8483
rect 16255 8449 16264 8483
rect 16212 8440 16264 8449
rect 16948 8483 17000 8492
rect 16948 8449 16957 8483
rect 16957 8449 16991 8483
rect 16991 8449 17000 8483
rect 16948 8440 17000 8449
rect 17592 8483 17644 8492
rect 17592 8449 17601 8483
rect 17601 8449 17635 8483
rect 17635 8449 17644 8483
rect 17592 8440 17644 8449
rect 17960 8483 18012 8492
rect 17960 8449 17969 8483
rect 17969 8449 18003 8483
rect 18003 8449 18012 8483
rect 17960 8440 18012 8449
rect 18144 8440 18196 8492
rect 19432 8508 19484 8560
rect 16488 8372 16540 8424
rect 12440 8304 12492 8356
rect 17776 8372 17828 8424
rect 18052 8304 18104 8356
rect 18880 8304 18932 8356
rect 29092 8508 29144 8560
rect 37188 8440 37240 8492
rect 38752 8440 38804 8492
rect 30748 8372 30800 8424
rect 35808 8372 35860 8424
rect 19708 8304 19760 8356
rect 38568 8304 38620 8356
rect 39672 8372 39724 8424
rect 40684 8483 40736 8492
rect 40684 8449 40693 8483
rect 40693 8449 40727 8483
rect 40727 8449 40736 8483
rect 40684 8440 40736 8449
rect 41420 8483 41472 8492
rect 41420 8449 41429 8483
rect 41429 8449 41463 8483
rect 41463 8449 41472 8483
rect 41420 8440 41472 8449
rect 41788 8483 41840 8492
rect 41788 8449 41797 8483
rect 41797 8449 41831 8483
rect 41831 8449 41840 8483
rect 41788 8440 41840 8449
rect 41880 8440 41932 8492
rect 42984 8440 43036 8492
rect 42248 8372 42300 8424
rect 43352 8440 43404 8492
rect 43720 8440 43772 8492
rect 43996 8440 44048 8492
rect 44916 8508 44968 8560
rect 46020 8576 46072 8628
rect 43628 8372 43680 8424
rect 44364 8440 44416 8492
rect 45468 8440 45520 8492
rect 46020 8440 46072 8492
rect 46572 8440 46624 8492
rect 42432 8304 42484 8356
rect 43168 8304 43220 8356
rect 44272 8304 44324 8356
rect 45468 8304 45520 8356
rect 46204 8372 46256 8424
rect 46388 8304 46440 8356
rect 39948 8236 40000 8288
rect 46020 8236 46072 8288
rect 1950 8134 2002 8186
rect 2014 8134 2066 8186
rect 2078 8134 2130 8186
rect 2142 8134 2194 8186
rect 2206 8134 2258 8186
rect 7950 8134 8002 8186
rect 8014 8134 8066 8186
rect 8078 8134 8130 8186
rect 8142 8134 8194 8186
rect 8206 8134 8258 8186
rect 13950 8134 14002 8186
rect 14014 8134 14066 8186
rect 14078 8134 14130 8186
rect 14142 8134 14194 8186
rect 14206 8134 14258 8186
rect 19950 8134 20002 8186
rect 20014 8134 20066 8186
rect 20078 8134 20130 8186
rect 20142 8134 20194 8186
rect 20206 8134 20258 8186
rect 25950 8134 26002 8186
rect 26014 8134 26066 8186
rect 26078 8134 26130 8186
rect 26142 8134 26194 8186
rect 26206 8134 26258 8186
rect 31950 8134 32002 8186
rect 32014 8134 32066 8186
rect 32078 8134 32130 8186
rect 32142 8134 32194 8186
rect 32206 8134 32258 8186
rect 37950 8134 38002 8186
rect 38014 8134 38066 8186
rect 38078 8134 38130 8186
rect 38142 8134 38194 8186
rect 38206 8134 38258 8186
rect 43950 8134 44002 8186
rect 44014 8134 44066 8186
rect 44078 8134 44130 8186
rect 44142 8134 44194 8186
rect 44206 8134 44258 8186
rect 1584 8075 1636 8084
rect 1584 8041 1593 8075
rect 1593 8041 1627 8075
rect 1627 8041 1636 8075
rect 1584 8032 1636 8041
rect 3792 8032 3844 8084
rect 6368 8032 6420 8084
rect 8852 8032 8904 8084
rect 10876 8032 10928 8084
rect 11428 8032 11480 8084
rect 11520 8032 11572 8084
rect 12440 8032 12492 8084
rect 12992 8032 13044 8084
rect 13728 8032 13780 8084
rect 14280 8032 14332 8084
rect 15108 8032 15160 8084
rect 16672 8032 16724 8084
rect 17040 8032 17092 8084
rect 17592 8032 17644 8084
rect 17960 8032 18012 8084
rect 19432 8075 19484 8084
rect 19432 8041 19441 8075
rect 19441 8041 19475 8075
rect 19475 8041 19484 8075
rect 19432 8032 19484 8041
rect 19708 8032 19760 8084
rect 21364 8032 21416 8084
rect 22652 8032 22704 8084
rect 24124 8032 24176 8084
rect 30196 8075 30248 8084
rect 30196 8041 30205 8075
rect 30205 8041 30239 8075
rect 30239 8041 30248 8075
rect 30196 8032 30248 8041
rect 35072 8032 35124 8084
rect 5356 8007 5408 8016
rect 5356 7973 5365 8007
rect 5365 7973 5399 8007
rect 5399 7973 5408 8007
rect 5356 7964 5408 7973
rect 13636 7964 13688 8016
rect 14464 7964 14516 8016
rect 18052 7964 18104 8016
rect 12440 7896 12492 7948
rect 13176 7896 13228 7948
rect 16304 7896 16356 7948
rect 2412 7871 2464 7880
rect 2412 7837 2421 7871
rect 2421 7837 2455 7871
rect 2455 7837 2464 7871
rect 2412 7828 2464 7837
rect 4160 7871 4212 7880
rect 4160 7837 4169 7871
rect 4169 7837 4203 7871
rect 4203 7837 4212 7871
rect 4160 7828 4212 7837
rect 5172 7871 5224 7880
rect 5172 7837 5181 7871
rect 5181 7837 5215 7871
rect 5215 7837 5224 7871
rect 5172 7828 5224 7837
rect 6736 7871 6788 7880
rect 6736 7837 6745 7871
rect 6745 7837 6779 7871
rect 6779 7837 6788 7871
rect 6736 7828 6788 7837
rect 9588 7828 9640 7880
rect 11796 7828 11848 7880
rect 11980 7871 12032 7880
rect 11980 7837 11989 7871
rect 11989 7837 12023 7871
rect 12023 7837 12032 7871
rect 11980 7828 12032 7837
rect 12532 7871 12584 7880
rect 12532 7837 12534 7871
rect 12534 7837 12568 7871
rect 12568 7837 12584 7871
rect 12532 7828 12584 7837
rect 13544 7871 13596 7880
rect 13544 7837 13553 7871
rect 13553 7837 13587 7871
rect 13587 7837 13596 7871
rect 13544 7828 13596 7837
rect 204 7760 256 7812
rect 14556 7871 14608 7880
rect 14556 7837 14565 7871
rect 14565 7837 14599 7871
rect 14599 7837 14608 7871
rect 14556 7828 14608 7837
rect 16764 7871 16816 7880
rect 16764 7837 16773 7871
rect 16773 7837 16807 7871
rect 16807 7837 16816 7871
rect 16764 7828 16816 7837
rect 17132 7871 17184 7880
rect 17132 7837 17141 7871
rect 17141 7837 17175 7871
rect 17175 7837 17184 7871
rect 17132 7828 17184 7837
rect 18236 7828 18288 7880
rect 18328 7871 18380 7880
rect 18328 7837 18337 7871
rect 18337 7837 18371 7871
rect 18371 7837 18380 7871
rect 18328 7828 18380 7837
rect 18880 7896 18932 7948
rect 24124 7896 24176 7948
rect 39948 7964 40000 8016
rect 40500 8075 40552 8084
rect 40500 8041 40509 8075
rect 40509 8041 40543 8075
rect 40543 8041 40552 8075
rect 40500 8032 40552 8041
rect 41604 8075 41656 8084
rect 41604 8041 41613 8075
rect 41613 8041 41647 8075
rect 41647 8041 41656 8075
rect 41604 8032 41656 8041
rect 44824 8032 44876 8084
rect 45652 8075 45704 8084
rect 45652 8041 45661 8075
rect 45661 8041 45695 8075
rect 45695 8041 45704 8075
rect 45652 8032 45704 8041
rect 46480 8032 46532 8084
rect 46848 8032 46900 8084
rect 19800 7828 19852 7880
rect 20444 7828 20496 7880
rect 20536 7828 20588 7880
rect 21640 7828 21692 7880
rect 27712 7896 27764 7948
rect 26608 7828 26660 7880
rect 26884 7828 26936 7880
rect 27344 7828 27396 7880
rect 29552 7896 29604 7948
rect 29920 7828 29972 7880
rect 34704 7896 34756 7948
rect 32496 7828 32548 7880
rect 38292 7828 38344 7880
rect 46020 8007 46072 8016
rect 46020 7973 46029 8007
rect 46029 7973 46063 8007
rect 46063 7973 46072 8007
rect 46020 7964 46072 7973
rect 47216 7964 47268 8016
rect 44548 7896 44600 7948
rect 45100 7871 45152 7880
rect 45100 7837 45109 7871
rect 45109 7837 45143 7871
rect 45143 7837 45152 7871
rect 45100 7828 45152 7837
rect 14280 7760 14332 7812
rect 21364 7760 21416 7812
rect 25780 7760 25832 7812
rect 15568 7692 15620 7744
rect 17868 7692 17920 7744
rect 18788 7735 18840 7744
rect 18788 7701 18797 7735
rect 18797 7701 18831 7735
rect 18831 7701 18840 7735
rect 18788 7692 18840 7701
rect 18972 7692 19024 7744
rect 21640 7692 21692 7744
rect 21732 7735 21784 7744
rect 21732 7701 21741 7735
rect 21741 7701 21775 7735
rect 21775 7701 21784 7735
rect 21732 7692 21784 7701
rect 22652 7692 22704 7744
rect 28264 7735 28316 7744
rect 28264 7701 28273 7735
rect 28273 7701 28307 7735
rect 28307 7701 28316 7735
rect 28264 7692 28316 7701
rect 29828 7760 29880 7812
rect 30564 7735 30616 7744
rect 30564 7701 30573 7735
rect 30573 7701 30607 7735
rect 30607 7701 30616 7735
rect 30564 7692 30616 7701
rect 30748 7760 30800 7812
rect 39580 7760 39632 7812
rect 45836 7871 45888 7880
rect 45836 7837 45845 7871
rect 45845 7837 45879 7871
rect 45879 7837 45888 7871
rect 45836 7828 45888 7837
rect 46204 7871 46256 7880
rect 46204 7837 46213 7871
rect 46213 7837 46247 7871
rect 46247 7837 46256 7871
rect 46204 7828 46256 7837
rect 46664 7828 46716 7880
rect 43720 7692 43772 7744
rect 3010 7590 3062 7642
rect 3074 7590 3126 7642
rect 3138 7590 3190 7642
rect 3202 7590 3254 7642
rect 3266 7590 3318 7642
rect 9010 7590 9062 7642
rect 9074 7590 9126 7642
rect 9138 7590 9190 7642
rect 9202 7590 9254 7642
rect 9266 7590 9318 7642
rect 15010 7590 15062 7642
rect 15074 7590 15126 7642
rect 15138 7590 15190 7642
rect 15202 7590 15254 7642
rect 15266 7590 15318 7642
rect 21010 7590 21062 7642
rect 21074 7590 21126 7642
rect 21138 7590 21190 7642
rect 21202 7590 21254 7642
rect 21266 7590 21318 7642
rect 27010 7590 27062 7642
rect 27074 7590 27126 7642
rect 27138 7590 27190 7642
rect 27202 7590 27254 7642
rect 27266 7590 27318 7642
rect 33010 7590 33062 7642
rect 33074 7590 33126 7642
rect 33138 7590 33190 7642
rect 33202 7590 33254 7642
rect 33266 7590 33318 7642
rect 39010 7590 39062 7642
rect 39074 7590 39126 7642
rect 39138 7590 39190 7642
rect 39202 7590 39254 7642
rect 39266 7590 39318 7642
rect 45010 7590 45062 7642
rect 45074 7590 45126 7642
rect 45138 7590 45190 7642
rect 45202 7590 45254 7642
rect 45266 7590 45318 7642
rect 4160 7488 4212 7540
rect 13728 7488 13780 7540
rect 15476 7488 15528 7540
rect 15844 7488 15896 7540
rect 16212 7488 16264 7540
rect 16948 7488 17000 7540
rect 7748 7463 7800 7472
rect 7748 7429 7757 7463
rect 7757 7429 7791 7463
rect 7791 7429 7800 7463
rect 7748 7420 7800 7429
rect 8300 7420 8352 7472
rect 14924 7352 14976 7404
rect 15476 7395 15528 7404
rect 16488 7420 16540 7472
rect 18880 7420 18932 7472
rect 30564 7488 30616 7540
rect 39580 7488 39632 7540
rect 44088 7488 44140 7540
rect 44548 7531 44600 7540
rect 44548 7497 44557 7531
rect 44557 7497 44591 7531
rect 44591 7497 44600 7531
rect 44548 7488 44600 7497
rect 46204 7488 46256 7540
rect 46572 7531 46624 7540
rect 46572 7497 46581 7531
rect 46581 7497 46615 7531
rect 46615 7497 46624 7531
rect 46572 7488 46624 7497
rect 46940 7531 46992 7540
rect 46940 7497 46949 7531
rect 46949 7497 46983 7531
rect 46983 7497 46992 7531
rect 46940 7488 46992 7497
rect 47308 7531 47360 7540
rect 47308 7497 47317 7531
rect 47317 7497 47351 7531
rect 47351 7497 47360 7531
rect 47308 7488 47360 7497
rect 25504 7420 25556 7472
rect 35900 7420 35952 7472
rect 15476 7361 15493 7395
rect 15493 7361 15527 7395
rect 15527 7361 15528 7395
rect 15476 7352 15528 7361
rect 16580 7352 16632 7404
rect 19156 7352 19208 7404
rect 20720 7352 20772 7404
rect 26332 7352 26384 7404
rect 32312 7352 32364 7404
rect 43628 7420 43680 7472
rect 6736 7284 6788 7336
rect 15384 7284 15436 7336
rect 15660 7284 15712 7336
rect 28264 7284 28316 7336
rect 40500 7284 40552 7336
rect 42800 7284 42852 7336
rect 45376 7395 45428 7404
rect 45376 7361 45385 7395
rect 45385 7361 45419 7395
rect 45419 7361 45428 7395
rect 45376 7352 45428 7361
rect 45652 7395 45704 7404
rect 45652 7361 45661 7395
rect 45661 7361 45695 7395
rect 45695 7361 45704 7395
rect 45652 7352 45704 7361
rect 45744 7352 45796 7404
rect 46756 7395 46808 7404
rect 46756 7361 46765 7395
rect 46765 7361 46799 7395
rect 46799 7361 46808 7395
rect 46756 7352 46808 7361
rect 47124 7395 47176 7404
rect 47124 7361 47133 7395
rect 47133 7361 47167 7395
rect 47167 7361 47176 7395
rect 47124 7352 47176 7361
rect 47216 7284 47268 7336
rect 7656 7216 7708 7268
rect 11244 7148 11296 7200
rect 14832 7148 14884 7200
rect 42892 7216 42944 7268
rect 45468 7216 45520 7268
rect 46664 7216 46716 7268
rect 16304 7148 16356 7200
rect 29828 7148 29880 7200
rect 33324 7191 33376 7200
rect 33324 7157 33333 7191
rect 33333 7157 33367 7191
rect 33367 7157 33376 7191
rect 33324 7148 33376 7157
rect 41604 7191 41656 7200
rect 41604 7157 41613 7191
rect 41613 7157 41647 7191
rect 41647 7157 41656 7191
rect 41604 7148 41656 7157
rect 45928 7148 45980 7200
rect 46296 7148 46348 7200
rect 1950 7046 2002 7098
rect 2014 7046 2066 7098
rect 2078 7046 2130 7098
rect 2142 7046 2194 7098
rect 2206 7046 2258 7098
rect 7950 7046 8002 7098
rect 8014 7046 8066 7098
rect 8078 7046 8130 7098
rect 8142 7046 8194 7098
rect 8206 7046 8258 7098
rect 13950 7046 14002 7098
rect 14014 7046 14066 7098
rect 14078 7046 14130 7098
rect 14142 7046 14194 7098
rect 14206 7046 14258 7098
rect 19950 7046 20002 7098
rect 20014 7046 20066 7098
rect 20078 7046 20130 7098
rect 20142 7046 20194 7098
rect 20206 7046 20258 7098
rect 25950 7046 26002 7098
rect 26014 7046 26066 7098
rect 26078 7046 26130 7098
rect 26142 7046 26194 7098
rect 26206 7046 26258 7098
rect 31950 7046 32002 7098
rect 32014 7046 32066 7098
rect 32078 7046 32130 7098
rect 32142 7046 32194 7098
rect 32206 7046 32258 7098
rect 37950 7046 38002 7098
rect 38014 7046 38066 7098
rect 38078 7046 38130 7098
rect 38142 7046 38194 7098
rect 38206 7046 38258 7098
rect 43950 7046 44002 7098
rect 44014 7046 44066 7098
rect 44078 7046 44130 7098
rect 44142 7046 44194 7098
rect 44206 7046 44258 7098
rect 12532 6944 12584 6996
rect 19340 6944 19392 6996
rect 36912 6944 36964 6996
rect 45836 6944 45888 6996
rect 14832 6876 14884 6928
rect 33324 6876 33376 6928
rect 13636 6808 13688 6860
rect 16028 6740 16080 6792
rect 16396 6740 16448 6792
rect 17776 6808 17828 6860
rect 39396 6808 39448 6860
rect 43720 6808 43772 6860
rect 30288 6740 30340 6792
rect 31760 6740 31812 6792
rect 32864 6740 32916 6792
rect 45560 6740 45612 6792
rect 46112 6783 46164 6792
rect 46112 6749 46121 6783
rect 46121 6749 46155 6783
rect 46155 6749 46164 6783
rect 46112 6740 46164 6749
rect 46204 6740 46256 6792
rect 16764 6672 16816 6724
rect 17224 6672 17276 6724
rect 17132 6604 17184 6656
rect 23664 6647 23716 6656
rect 23664 6613 23673 6647
rect 23673 6613 23707 6647
rect 23707 6613 23716 6647
rect 23664 6604 23716 6613
rect 32772 6672 32824 6724
rect 29276 6604 29328 6656
rect 35348 6647 35400 6656
rect 35348 6613 35357 6647
rect 35357 6613 35391 6647
rect 35391 6613 35400 6647
rect 35348 6604 35400 6613
rect 46020 6647 46072 6656
rect 46020 6613 46029 6647
rect 46029 6613 46063 6647
rect 46063 6613 46072 6647
rect 46020 6604 46072 6613
rect 46296 6647 46348 6656
rect 46296 6613 46305 6647
rect 46305 6613 46339 6647
rect 46339 6613 46348 6647
rect 46296 6604 46348 6613
rect 46664 6647 46716 6656
rect 46664 6613 46673 6647
rect 46673 6613 46707 6647
rect 46707 6613 46716 6647
rect 46664 6604 46716 6613
rect 47032 6647 47084 6656
rect 47032 6613 47041 6647
rect 47041 6613 47075 6647
rect 47075 6613 47084 6647
rect 47032 6604 47084 6613
rect 47400 6647 47452 6656
rect 47400 6613 47409 6647
rect 47409 6613 47443 6647
rect 47443 6613 47452 6647
rect 47400 6604 47452 6613
rect 3010 6502 3062 6554
rect 3074 6502 3126 6554
rect 3138 6502 3190 6554
rect 3202 6502 3254 6554
rect 3266 6502 3318 6554
rect 9010 6502 9062 6554
rect 9074 6502 9126 6554
rect 9138 6502 9190 6554
rect 9202 6502 9254 6554
rect 9266 6502 9318 6554
rect 15010 6502 15062 6554
rect 15074 6502 15126 6554
rect 15138 6502 15190 6554
rect 15202 6502 15254 6554
rect 15266 6502 15318 6554
rect 21010 6502 21062 6554
rect 21074 6502 21126 6554
rect 21138 6502 21190 6554
rect 21202 6502 21254 6554
rect 21266 6502 21318 6554
rect 27010 6502 27062 6554
rect 27074 6502 27126 6554
rect 27138 6502 27190 6554
rect 27202 6502 27254 6554
rect 27266 6502 27318 6554
rect 33010 6502 33062 6554
rect 33074 6502 33126 6554
rect 33138 6502 33190 6554
rect 33202 6502 33254 6554
rect 33266 6502 33318 6554
rect 39010 6502 39062 6554
rect 39074 6502 39126 6554
rect 39138 6502 39190 6554
rect 39202 6502 39254 6554
rect 39266 6502 39318 6554
rect 45010 6502 45062 6554
rect 45074 6502 45126 6554
rect 45138 6502 45190 6554
rect 45202 6502 45254 6554
rect 45266 6502 45318 6554
rect 12716 6400 12768 6452
rect 17224 6400 17276 6452
rect 23664 6400 23716 6452
rect 10968 6332 11020 6384
rect 29276 6332 29328 6384
rect 33416 6332 33468 6384
rect 38568 6400 38620 6452
rect 40040 6332 40092 6384
rect 16856 6264 16908 6316
rect 24492 6264 24544 6316
rect 25136 6264 25188 6316
rect 25596 6264 25648 6316
rect 7840 6196 7892 6248
rect 25780 6196 25832 6248
rect 25872 6196 25924 6248
rect 32404 6264 32456 6316
rect 34336 6264 34388 6316
rect 26516 6196 26568 6248
rect 46020 6332 46072 6384
rect 46388 6307 46440 6316
rect 46388 6273 46397 6307
rect 46397 6273 46431 6307
rect 46431 6273 46440 6307
rect 46388 6264 46440 6273
rect 46940 6443 46992 6452
rect 46940 6409 46949 6443
rect 46949 6409 46983 6443
rect 46983 6409 46992 6443
rect 46940 6400 46992 6409
rect 47492 6400 47544 6452
rect 8392 6128 8444 6180
rect 6828 6060 6880 6112
rect 22468 6060 22520 6112
rect 24492 6103 24544 6112
rect 24492 6069 24501 6103
rect 24501 6069 24535 6103
rect 24535 6069 24544 6103
rect 24492 6060 24544 6069
rect 24676 6060 24728 6112
rect 34428 6128 34480 6180
rect 36176 6171 36228 6180
rect 36176 6137 36185 6171
rect 36185 6137 36219 6171
rect 36219 6137 36228 6171
rect 36176 6128 36228 6137
rect 36268 6128 36320 6180
rect 46204 6128 46256 6180
rect 25872 6060 25924 6112
rect 33140 6103 33192 6112
rect 33140 6069 33149 6103
rect 33149 6069 33183 6103
rect 33183 6069 33192 6103
rect 33140 6060 33192 6069
rect 46572 6103 46624 6112
rect 46572 6069 46581 6103
rect 46581 6069 46615 6103
rect 46615 6069 46624 6103
rect 46572 6060 46624 6069
rect 1950 5958 2002 6010
rect 2014 5958 2066 6010
rect 2078 5958 2130 6010
rect 2142 5958 2194 6010
rect 2206 5958 2258 6010
rect 7950 5958 8002 6010
rect 8014 5958 8066 6010
rect 8078 5958 8130 6010
rect 8142 5958 8194 6010
rect 8206 5958 8258 6010
rect 13950 5958 14002 6010
rect 14014 5958 14066 6010
rect 14078 5958 14130 6010
rect 14142 5958 14194 6010
rect 14206 5958 14258 6010
rect 19950 5958 20002 6010
rect 20014 5958 20066 6010
rect 20078 5958 20130 6010
rect 20142 5958 20194 6010
rect 20206 5958 20258 6010
rect 25950 5958 26002 6010
rect 26014 5958 26066 6010
rect 26078 5958 26130 6010
rect 26142 5958 26194 6010
rect 26206 5958 26258 6010
rect 31950 5958 32002 6010
rect 32014 5958 32066 6010
rect 32078 5958 32130 6010
rect 32142 5958 32194 6010
rect 32206 5958 32258 6010
rect 37950 5958 38002 6010
rect 38014 5958 38066 6010
rect 38078 5958 38130 6010
rect 38142 5958 38194 6010
rect 38206 5958 38258 6010
rect 43950 5958 44002 6010
rect 44014 5958 44066 6010
rect 44078 5958 44130 6010
rect 44142 5958 44194 6010
rect 44206 5958 44258 6010
rect 11060 5856 11112 5908
rect 17776 5899 17828 5908
rect 17776 5865 17785 5899
rect 17785 5865 17819 5899
rect 17819 5865 17828 5899
rect 17776 5856 17828 5865
rect 22468 5899 22520 5908
rect 22468 5865 22477 5899
rect 22477 5865 22511 5899
rect 22511 5865 22520 5899
rect 22468 5856 22520 5865
rect 27620 5856 27672 5908
rect 12624 5788 12676 5840
rect 31208 5856 31260 5908
rect 46388 5856 46440 5908
rect 47400 5899 47452 5908
rect 47400 5865 47409 5899
rect 47409 5865 47443 5899
rect 47443 5865 47452 5899
rect 47400 5856 47452 5865
rect 12808 5720 12860 5772
rect 14924 5695 14976 5704
rect 14924 5661 14933 5695
rect 14933 5661 14967 5695
rect 14967 5661 14976 5695
rect 14924 5652 14976 5661
rect 19340 5720 19392 5772
rect 36268 5788 36320 5840
rect 37188 5788 37240 5840
rect 17408 5559 17460 5568
rect 17408 5525 17417 5559
rect 17417 5525 17451 5559
rect 17451 5525 17460 5559
rect 17408 5516 17460 5525
rect 24400 5652 24452 5704
rect 30656 5720 30708 5772
rect 33140 5720 33192 5772
rect 43628 5720 43680 5772
rect 31024 5652 31076 5704
rect 31392 5652 31444 5704
rect 33968 5652 34020 5704
rect 39396 5652 39448 5704
rect 24952 5584 25004 5636
rect 31208 5584 31260 5636
rect 44456 5584 44508 5636
rect 47032 5559 47084 5568
rect 47032 5525 47041 5559
rect 47041 5525 47075 5559
rect 47075 5525 47084 5559
rect 47032 5516 47084 5525
rect 3010 5414 3062 5466
rect 3074 5414 3126 5466
rect 3138 5414 3190 5466
rect 3202 5414 3254 5466
rect 3266 5414 3318 5466
rect 9010 5414 9062 5466
rect 9074 5414 9126 5466
rect 9138 5414 9190 5466
rect 9202 5414 9254 5466
rect 9266 5414 9318 5466
rect 15010 5414 15062 5466
rect 15074 5414 15126 5466
rect 15138 5414 15190 5466
rect 15202 5414 15254 5466
rect 15266 5414 15318 5466
rect 21010 5414 21062 5466
rect 21074 5414 21126 5466
rect 21138 5414 21190 5466
rect 21202 5414 21254 5466
rect 21266 5414 21318 5466
rect 27010 5414 27062 5466
rect 27074 5414 27126 5466
rect 27138 5414 27190 5466
rect 27202 5414 27254 5466
rect 27266 5414 27318 5466
rect 33010 5414 33062 5466
rect 33074 5414 33126 5466
rect 33138 5414 33190 5466
rect 33202 5414 33254 5466
rect 33266 5414 33318 5466
rect 39010 5414 39062 5466
rect 39074 5414 39126 5466
rect 39138 5414 39190 5466
rect 39202 5414 39254 5466
rect 39266 5414 39318 5466
rect 45010 5414 45062 5466
rect 45074 5414 45126 5466
rect 45138 5414 45190 5466
rect 45202 5414 45254 5466
rect 45266 5414 45318 5466
rect 13728 5312 13780 5364
rect 23388 5312 23440 5364
rect 6000 5244 6052 5296
rect 9588 5176 9640 5228
rect 23572 5244 23624 5296
rect 21916 5176 21968 5228
rect 24768 5176 24820 5228
rect 18788 5108 18840 5160
rect 18144 5040 18196 5092
rect 20352 4972 20404 5024
rect 21732 5040 21784 5092
rect 33600 5176 33652 5228
rect 47308 5355 47360 5364
rect 47308 5321 47317 5355
rect 47317 5321 47351 5355
rect 47351 5321 47360 5355
rect 47308 5312 47360 5321
rect 37556 5151 37608 5160
rect 37556 5117 37565 5151
rect 37565 5117 37599 5151
rect 37599 5117 37608 5151
rect 37556 5108 37608 5117
rect 34428 5040 34480 5092
rect 44364 5040 44416 5092
rect 27620 4972 27672 5024
rect 46940 5015 46992 5024
rect 46940 4981 46949 5015
rect 46949 4981 46983 5015
rect 46983 4981 46992 5015
rect 46940 4972 46992 4981
rect 1950 4870 2002 4922
rect 2014 4870 2066 4922
rect 2078 4870 2130 4922
rect 2142 4870 2194 4922
rect 2206 4870 2258 4922
rect 7950 4870 8002 4922
rect 8014 4870 8066 4922
rect 8078 4870 8130 4922
rect 8142 4870 8194 4922
rect 8206 4870 8258 4922
rect 13950 4870 14002 4922
rect 14014 4870 14066 4922
rect 14078 4870 14130 4922
rect 14142 4870 14194 4922
rect 14206 4870 14258 4922
rect 19950 4870 20002 4922
rect 20014 4870 20066 4922
rect 20078 4870 20130 4922
rect 20142 4870 20194 4922
rect 20206 4870 20258 4922
rect 25950 4870 26002 4922
rect 26014 4870 26066 4922
rect 26078 4870 26130 4922
rect 26142 4870 26194 4922
rect 26206 4870 26258 4922
rect 31950 4870 32002 4922
rect 32014 4870 32066 4922
rect 32078 4870 32130 4922
rect 32142 4870 32194 4922
rect 32206 4870 32258 4922
rect 37950 4870 38002 4922
rect 38014 4870 38066 4922
rect 38078 4870 38130 4922
rect 38142 4870 38194 4922
rect 38206 4870 38258 4922
rect 43950 4870 44002 4922
rect 44014 4870 44066 4922
rect 44078 4870 44130 4922
rect 44142 4870 44194 4922
rect 44206 4870 44258 4922
rect 18052 4811 18104 4820
rect 18052 4777 18061 4811
rect 18061 4777 18095 4811
rect 18095 4777 18104 4811
rect 18052 4768 18104 4777
rect 19800 4768 19852 4820
rect 24952 4768 25004 4820
rect 8668 4700 8720 4752
rect 17224 4632 17276 4684
rect 47124 4768 47176 4820
rect 18236 4607 18288 4616
rect 18236 4573 18245 4607
rect 18245 4573 18279 4607
rect 18279 4573 18288 4607
rect 18236 4564 18288 4573
rect 22928 4632 22980 4684
rect 23112 4632 23164 4684
rect 47400 4743 47452 4752
rect 47400 4709 47409 4743
rect 47409 4709 47443 4743
rect 47443 4709 47452 4743
rect 47400 4700 47452 4709
rect 25504 4632 25556 4684
rect 23204 4564 23256 4616
rect 40040 4564 40092 4616
rect 8484 4496 8536 4548
rect 47124 4496 47176 4548
rect 24860 4471 24912 4480
rect 24860 4437 24869 4471
rect 24869 4437 24903 4471
rect 24903 4437 24912 4471
rect 24860 4428 24912 4437
rect 25228 4471 25280 4480
rect 25228 4437 25237 4471
rect 25237 4437 25271 4471
rect 25271 4437 25280 4471
rect 25228 4428 25280 4437
rect 47032 4471 47084 4480
rect 47032 4437 47041 4471
rect 47041 4437 47075 4471
rect 47075 4437 47084 4471
rect 47032 4428 47084 4437
rect 3010 4326 3062 4378
rect 3074 4326 3126 4378
rect 3138 4326 3190 4378
rect 3202 4326 3254 4378
rect 3266 4326 3318 4378
rect 9010 4326 9062 4378
rect 9074 4326 9126 4378
rect 9138 4326 9190 4378
rect 9202 4326 9254 4378
rect 9266 4326 9318 4378
rect 15010 4326 15062 4378
rect 15074 4326 15126 4378
rect 15138 4326 15190 4378
rect 15202 4326 15254 4378
rect 15266 4326 15318 4378
rect 21010 4326 21062 4378
rect 21074 4326 21126 4378
rect 21138 4326 21190 4378
rect 21202 4326 21254 4378
rect 21266 4326 21318 4378
rect 27010 4326 27062 4378
rect 27074 4326 27126 4378
rect 27138 4326 27190 4378
rect 27202 4326 27254 4378
rect 27266 4326 27318 4378
rect 33010 4326 33062 4378
rect 33074 4326 33126 4378
rect 33138 4326 33190 4378
rect 33202 4326 33254 4378
rect 33266 4326 33318 4378
rect 39010 4326 39062 4378
rect 39074 4326 39126 4378
rect 39138 4326 39190 4378
rect 39202 4326 39254 4378
rect 39266 4326 39318 4378
rect 45010 4326 45062 4378
rect 45074 4326 45126 4378
rect 45138 4326 45190 4378
rect 45202 4326 45254 4378
rect 45266 4326 45318 4378
rect 25228 4224 25280 4276
rect 42708 4224 42760 4276
rect 21456 4088 21508 4140
rect 12992 3952 13044 4004
rect 2596 3884 2648 3936
rect 15752 3884 15804 3936
rect 21824 4020 21876 4072
rect 17960 3995 18012 4004
rect 17960 3961 17969 3995
rect 17969 3961 18003 3995
rect 18003 3961 18012 3995
rect 17960 3952 18012 3961
rect 44364 4020 44416 4072
rect 47308 3995 47360 4004
rect 47308 3961 47317 3995
rect 47317 3961 47351 3995
rect 47351 3961 47360 3995
rect 47308 3952 47360 3961
rect 19524 3884 19576 3936
rect 20720 3884 20772 3936
rect 25872 3884 25924 3936
rect 37648 3884 37700 3936
rect 46756 3884 46808 3936
rect 46940 3927 46992 3936
rect 46940 3893 46949 3927
rect 46949 3893 46983 3927
rect 46983 3893 46992 3927
rect 46940 3884 46992 3893
rect 1950 3782 2002 3834
rect 2014 3782 2066 3834
rect 2078 3782 2130 3834
rect 2142 3782 2194 3834
rect 2206 3782 2258 3834
rect 7950 3782 8002 3834
rect 8014 3782 8066 3834
rect 8078 3782 8130 3834
rect 8142 3782 8194 3834
rect 8206 3782 8258 3834
rect 13950 3782 14002 3834
rect 14014 3782 14066 3834
rect 14078 3782 14130 3834
rect 14142 3782 14194 3834
rect 14206 3782 14258 3834
rect 19950 3782 20002 3834
rect 20014 3782 20066 3834
rect 20078 3782 20130 3834
rect 20142 3782 20194 3834
rect 20206 3782 20258 3834
rect 25950 3782 26002 3834
rect 26014 3782 26066 3834
rect 26078 3782 26130 3834
rect 26142 3782 26194 3834
rect 26206 3782 26258 3834
rect 31950 3782 32002 3834
rect 32014 3782 32066 3834
rect 32078 3782 32130 3834
rect 32142 3782 32194 3834
rect 32206 3782 32258 3834
rect 37950 3782 38002 3834
rect 38014 3782 38066 3834
rect 38078 3782 38130 3834
rect 38142 3782 38194 3834
rect 38206 3782 38258 3834
rect 43950 3782 44002 3834
rect 44014 3782 44066 3834
rect 44078 3782 44130 3834
rect 44142 3782 44194 3834
rect 44206 3782 44258 3834
rect 43352 3680 43404 3732
rect 12808 3612 12860 3664
rect 41788 3612 41840 3664
rect 47400 3655 47452 3664
rect 47400 3621 47409 3655
rect 47409 3621 47443 3655
rect 47443 3621 47452 3655
rect 47400 3612 47452 3621
rect 8852 3544 8904 3596
rect 2320 3408 2372 3460
rect 6920 3408 6972 3460
rect 22100 3476 22152 3528
rect 24768 3544 24820 3596
rect 29092 3544 29144 3596
rect 42708 3544 42760 3596
rect 22560 3408 22612 3460
rect 29460 3476 29512 3528
rect 44180 3476 44232 3528
rect 20904 3340 20956 3392
rect 23020 3340 23072 3392
rect 27436 3408 27488 3460
rect 40776 3408 40828 3460
rect 28540 3340 28592 3392
rect 33600 3340 33652 3392
rect 43812 3340 43864 3392
rect 47032 3383 47084 3392
rect 47032 3349 47041 3383
rect 47041 3349 47075 3383
rect 47075 3349 47084 3383
rect 47032 3340 47084 3349
rect 3010 3238 3062 3290
rect 3074 3238 3126 3290
rect 3138 3238 3190 3290
rect 3202 3238 3254 3290
rect 3266 3238 3318 3290
rect 9010 3238 9062 3290
rect 9074 3238 9126 3290
rect 9138 3238 9190 3290
rect 9202 3238 9254 3290
rect 9266 3238 9318 3290
rect 15010 3238 15062 3290
rect 15074 3238 15126 3290
rect 15138 3238 15190 3290
rect 15202 3238 15254 3290
rect 15266 3238 15318 3290
rect 21010 3238 21062 3290
rect 21074 3238 21126 3290
rect 21138 3238 21190 3290
rect 21202 3238 21254 3290
rect 21266 3238 21318 3290
rect 27010 3238 27062 3290
rect 27074 3238 27126 3290
rect 27138 3238 27190 3290
rect 27202 3238 27254 3290
rect 27266 3238 27318 3290
rect 33010 3238 33062 3290
rect 33074 3238 33126 3290
rect 33138 3238 33190 3290
rect 33202 3238 33254 3290
rect 33266 3238 33318 3290
rect 39010 3238 39062 3290
rect 39074 3238 39126 3290
rect 39138 3238 39190 3290
rect 39202 3238 39254 3290
rect 39266 3238 39318 3290
rect 45010 3238 45062 3290
rect 45074 3238 45126 3290
rect 45138 3238 45190 3290
rect 45202 3238 45254 3290
rect 45266 3238 45318 3290
rect 8852 3179 8904 3188
rect 8852 3145 8861 3179
rect 8861 3145 8895 3179
rect 8895 3145 8904 3179
rect 8852 3136 8904 3145
rect 12808 3179 12860 3188
rect 12808 3145 12817 3179
rect 12817 3145 12851 3179
rect 12851 3145 12860 3179
rect 12808 3136 12860 3145
rect 13544 3136 13596 3188
rect 23020 3136 23072 3188
rect 23112 3179 23164 3188
rect 23112 3145 23121 3179
rect 23121 3145 23155 3179
rect 23155 3145 23164 3179
rect 23112 3136 23164 3145
rect 26700 3136 26752 3188
rect 8300 3068 8352 3120
rect 9588 3068 9640 3120
rect 18144 3111 18196 3120
rect 18144 3077 18153 3111
rect 18153 3077 18187 3111
rect 18187 3077 18196 3111
rect 18144 3068 18196 3077
rect 19800 3068 19852 3120
rect 10600 3000 10652 3052
rect 12900 3000 12952 3052
rect 15384 3000 15436 3052
rect 11060 2975 11112 2984
rect 11060 2941 11069 2975
rect 11069 2941 11103 2975
rect 11103 2941 11112 2975
rect 11060 2932 11112 2941
rect 8576 2907 8628 2916
rect 8576 2873 8585 2907
rect 8585 2873 8619 2907
rect 8619 2873 8628 2907
rect 8576 2864 8628 2873
rect 9496 2864 9548 2916
rect 17500 2932 17552 2984
rect 22744 3043 22796 3052
rect 22744 3009 22753 3043
rect 22753 3009 22787 3043
rect 22787 3009 22796 3043
rect 22744 3000 22796 3009
rect 24400 3068 24452 3120
rect 25320 3043 25372 3052
rect 25320 3009 25329 3043
rect 25329 3009 25363 3043
rect 25363 3009 25372 3043
rect 25320 3000 25372 3009
rect 27528 3043 27580 3052
rect 27528 3009 27537 3043
rect 27537 3009 27571 3043
rect 27571 3009 27580 3043
rect 27528 3000 27580 3009
rect 29368 3136 29420 3188
rect 29460 3000 29512 3052
rect 32036 3136 32088 3188
rect 37740 3136 37792 3188
rect 38752 3179 38804 3188
rect 38752 3145 38761 3179
rect 38761 3145 38795 3179
rect 38795 3145 38804 3179
rect 38752 3136 38804 3145
rect 39672 3179 39724 3188
rect 39672 3145 39681 3179
rect 39681 3145 39715 3179
rect 39715 3145 39724 3179
rect 39672 3136 39724 3145
rect 40684 3136 40736 3188
rect 43260 3179 43312 3188
rect 43260 3145 43269 3179
rect 43269 3145 43303 3179
rect 43303 3145 43312 3179
rect 43260 3136 43312 3145
rect 43904 3136 43956 3188
rect 47308 3179 47360 3188
rect 47308 3145 47317 3179
rect 47317 3145 47351 3179
rect 47351 3145 47360 3179
rect 47308 3136 47360 3145
rect 44456 3068 44508 3120
rect 13268 2907 13320 2916
rect 13268 2873 13277 2907
rect 13277 2873 13311 2907
rect 13311 2873 13320 2907
rect 13268 2864 13320 2873
rect 1308 2796 1360 2848
rect 16856 2839 16908 2848
rect 16856 2805 16865 2839
rect 16865 2805 16899 2839
rect 16899 2805 16908 2839
rect 16856 2796 16908 2805
rect 31760 2932 31812 2984
rect 36452 3000 36504 3052
rect 37280 3043 37332 3052
rect 37280 3009 37289 3043
rect 37289 3009 37323 3043
rect 37323 3009 37332 3043
rect 37280 3000 37332 3009
rect 38568 3043 38620 3052
rect 38568 3009 38577 3043
rect 38577 3009 38611 3043
rect 38611 3009 38620 3043
rect 38568 3000 38620 3009
rect 39488 3043 39540 3052
rect 39488 3009 39497 3043
rect 39497 3009 39531 3043
rect 39531 3009 39540 3043
rect 39488 3000 39540 3009
rect 40316 3043 40368 3052
rect 40316 3009 40325 3043
rect 40325 3009 40359 3043
rect 40359 3009 40368 3043
rect 40316 3000 40368 3009
rect 43076 3043 43128 3052
rect 43076 3009 43085 3043
rect 43085 3009 43119 3043
rect 43119 3009 43128 3043
rect 43076 3000 43128 3009
rect 43812 3043 43864 3052
rect 43812 3009 43821 3043
rect 43821 3009 43855 3043
rect 43855 3009 43864 3043
rect 43812 3000 43864 3009
rect 46756 3043 46808 3052
rect 46756 3009 46765 3043
rect 46765 3009 46799 3043
rect 46799 3009 46808 3043
rect 46756 3000 46808 3009
rect 47124 3043 47176 3052
rect 47124 3009 47133 3043
rect 47133 3009 47167 3043
rect 47167 3009 47176 3043
rect 47124 3000 47176 3009
rect 42248 2932 42300 2984
rect 41880 2864 41932 2916
rect 19708 2796 19760 2848
rect 20444 2839 20496 2848
rect 20444 2805 20453 2839
rect 20453 2805 20487 2839
rect 20487 2805 20496 2839
rect 20444 2796 20496 2805
rect 20720 2839 20772 2848
rect 20720 2805 20729 2839
rect 20729 2805 20763 2839
rect 20763 2805 20772 2839
rect 20720 2796 20772 2805
rect 21088 2839 21140 2848
rect 21088 2805 21097 2839
rect 21097 2805 21131 2839
rect 21131 2805 21140 2839
rect 21088 2796 21140 2805
rect 26516 2796 26568 2848
rect 27436 2839 27488 2848
rect 27436 2805 27445 2839
rect 27445 2805 27479 2839
rect 27479 2805 27488 2839
rect 27436 2796 27488 2805
rect 29368 2796 29420 2848
rect 35808 2796 35860 2848
rect 36912 2839 36964 2848
rect 36912 2805 36921 2839
rect 36921 2805 36955 2839
rect 36955 2805 36964 2839
rect 36912 2796 36964 2805
rect 37648 2839 37700 2848
rect 37648 2805 37657 2839
rect 37657 2805 37691 2839
rect 37691 2805 37700 2839
rect 37648 2796 37700 2805
rect 37740 2796 37792 2848
rect 42984 2796 43036 2848
rect 46940 2839 46992 2848
rect 46940 2805 46949 2839
rect 46949 2805 46983 2839
rect 46983 2805 46992 2839
rect 46940 2796 46992 2805
rect 1950 2694 2002 2746
rect 2014 2694 2066 2746
rect 2078 2694 2130 2746
rect 2142 2694 2194 2746
rect 2206 2694 2258 2746
rect 7950 2694 8002 2746
rect 8014 2694 8066 2746
rect 8078 2694 8130 2746
rect 8142 2694 8194 2746
rect 8206 2694 8258 2746
rect 13950 2694 14002 2746
rect 14014 2694 14066 2746
rect 14078 2694 14130 2746
rect 14142 2694 14194 2746
rect 14206 2694 14258 2746
rect 19950 2694 20002 2746
rect 20014 2694 20066 2746
rect 20078 2694 20130 2746
rect 20142 2694 20194 2746
rect 20206 2694 20258 2746
rect 25950 2694 26002 2746
rect 26014 2694 26066 2746
rect 26078 2694 26130 2746
rect 26142 2694 26194 2746
rect 26206 2694 26258 2746
rect 31950 2694 32002 2746
rect 32014 2694 32066 2746
rect 32078 2694 32130 2746
rect 32142 2694 32194 2746
rect 32206 2694 32258 2746
rect 37950 2694 38002 2746
rect 38014 2694 38066 2746
rect 38078 2694 38130 2746
rect 38142 2694 38194 2746
rect 38206 2694 38258 2746
rect 43950 2694 44002 2746
rect 44014 2694 44066 2746
rect 44078 2694 44130 2746
rect 44142 2694 44194 2746
rect 44206 2694 44258 2746
rect 20444 2592 20496 2644
rect 42156 2592 42208 2644
rect 16856 2524 16908 2576
rect 45836 2635 45888 2644
rect 45836 2601 45845 2635
rect 45845 2601 45879 2635
rect 45879 2601 45888 2635
rect 45836 2592 45888 2601
rect 13268 2456 13320 2508
rect 33140 2456 33192 2508
rect 8576 2388 8628 2440
rect 36268 2388 36320 2440
rect 36452 2388 36504 2440
rect 45652 2431 45704 2440
rect 45652 2397 45661 2431
rect 45661 2397 45695 2431
rect 45695 2397 45704 2431
rect 45652 2388 45704 2397
rect 47308 2567 47360 2576
rect 47308 2533 47317 2567
rect 47317 2533 47351 2567
rect 47351 2533 47360 2567
rect 47308 2524 47360 2533
rect 21088 2320 21140 2372
rect 5632 2252 5684 2304
rect 27528 2252 27580 2304
rect 33140 2320 33192 2372
rect 46204 2295 46256 2304
rect 46204 2261 46213 2295
rect 46213 2261 46247 2295
rect 46247 2261 46256 2295
rect 46204 2252 46256 2261
rect 46572 2295 46624 2304
rect 46572 2261 46581 2295
rect 46581 2261 46615 2295
rect 46615 2261 46624 2295
rect 46572 2252 46624 2261
rect 46940 2295 46992 2304
rect 46940 2261 46949 2295
rect 46949 2261 46983 2295
rect 46983 2261 46992 2295
rect 46940 2252 46992 2261
rect 3010 2150 3062 2202
rect 3074 2150 3126 2202
rect 3138 2150 3190 2202
rect 3202 2150 3254 2202
rect 3266 2150 3318 2202
rect 9010 2150 9062 2202
rect 9074 2150 9126 2202
rect 9138 2150 9190 2202
rect 9202 2150 9254 2202
rect 9266 2150 9318 2202
rect 15010 2150 15062 2202
rect 15074 2150 15126 2202
rect 15138 2150 15190 2202
rect 15202 2150 15254 2202
rect 15266 2150 15318 2202
rect 21010 2150 21062 2202
rect 21074 2150 21126 2202
rect 21138 2150 21190 2202
rect 21202 2150 21254 2202
rect 21266 2150 21318 2202
rect 27010 2150 27062 2202
rect 27074 2150 27126 2202
rect 27138 2150 27190 2202
rect 27202 2150 27254 2202
rect 27266 2150 27318 2202
rect 33010 2150 33062 2202
rect 33074 2150 33126 2202
rect 33138 2150 33190 2202
rect 33202 2150 33254 2202
rect 33266 2150 33318 2202
rect 39010 2150 39062 2202
rect 39074 2150 39126 2202
rect 39138 2150 39190 2202
rect 39202 2150 39254 2202
rect 39266 2150 39318 2202
rect 45010 2150 45062 2202
rect 45074 2150 45126 2202
rect 45138 2150 45190 2202
rect 45202 2150 45254 2202
rect 45266 2150 45318 2202
rect 2872 2048 2924 2100
rect 25320 2048 25372 2100
rect 31300 2048 31352 2100
rect 43076 2048 43128 2100
rect 3700 144 3752 196
rect 6000 144 6052 196
rect 40316 144 40368 196
rect 39488 76 39540 128
rect 1492 8 1544 60
rect 38568 8 38620 60
<< metal2 >>
rect 1582 11194 1638 11250
rect 1950 11194 2006 11250
rect 2318 11194 2374 11250
rect 2686 11194 2742 11250
rect 3054 11194 3110 11250
rect 3422 11194 3478 11250
rect 3790 11194 3846 11250
rect 4158 11194 4214 11250
rect 4526 11194 4582 11250
rect 4894 11194 4950 11250
rect 5262 11194 5318 11250
rect 5630 11194 5686 11250
rect 5998 11194 6054 11250
rect 6366 11194 6422 11250
rect 6734 11194 6790 11250
rect 7102 11194 7158 11250
rect 7470 11194 7526 11250
rect 7838 11194 7894 11250
rect 8206 11194 8262 11250
rect 8574 11194 8630 11250
rect 8942 11194 8998 11250
rect 9310 11194 9366 11250
rect 9678 11194 9734 11250
rect 10046 11194 10102 11250
rect 10414 11194 10470 11250
rect 10782 11194 10838 11250
rect 11150 11194 11206 11250
rect 11518 11194 11574 11250
rect 11886 11194 11942 11250
rect 12254 11194 12310 11250
rect 12622 11194 12678 11250
rect 12990 11194 13046 11250
rect 13358 11194 13414 11250
rect 13544 11212 13596 11218
rect 1122 9480 1178 9489
rect 1122 9415 1178 9424
rect 202 9344 258 9353
rect 202 9279 258 9288
rect 216 7818 244 9279
rect 204 7812 256 7818
rect 204 7754 256 7760
rect 1136 7449 1164 9415
rect 1308 9376 1360 9382
rect 1308 9318 1360 9324
rect 1320 8265 1348 9318
rect 1306 8256 1362 8265
rect 1306 8191 1362 8200
rect 1596 8090 1624 11194
rect 1964 8634 1992 11194
rect 2332 8634 2360 11194
rect 2700 8634 2728 11194
rect 3068 9738 3096 11194
rect 2884 9710 3096 9738
rect 2884 8634 2912 9710
rect 3010 8732 3318 8741
rect 3010 8730 3016 8732
rect 3072 8730 3096 8732
rect 3152 8730 3176 8732
rect 3232 8730 3256 8732
rect 3312 8730 3318 8732
rect 3072 8678 3074 8730
rect 3254 8678 3256 8730
rect 3010 8676 3016 8678
rect 3072 8676 3096 8678
rect 3152 8676 3176 8678
rect 3232 8676 3256 8678
rect 3312 8676 3318 8678
rect 3010 8667 3318 8676
rect 3436 8634 3464 11194
rect 3516 9036 3568 9042
rect 3516 8978 3568 8984
rect 1952 8628 2004 8634
rect 1952 8570 2004 8576
rect 2320 8628 2372 8634
rect 2320 8570 2372 8576
rect 2688 8628 2740 8634
rect 2688 8570 2740 8576
rect 2872 8628 2924 8634
rect 2872 8570 2924 8576
rect 3424 8628 3476 8634
rect 3424 8570 3476 8576
rect 3528 8498 3556 8978
rect 2320 8492 2372 8498
rect 2320 8434 2372 8440
rect 2596 8492 2648 8498
rect 2596 8434 2648 8440
rect 3516 8492 3568 8498
rect 3516 8434 3568 8440
rect 1950 8188 2258 8197
rect 1950 8186 1956 8188
rect 2012 8186 2036 8188
rect 2092 8186 2116 8188
rect 2172 8186 2196 8188
rect 2252 8186 2258 8188
rect 2012 8134 2014 8186
rect 2194 8134 2196 8186
rect 1950 8132 1956 8134
rect 2012 8132 2036 8134
rect 2092 8132 2116 8134
rect 2172 8132 2196 8134
rect 2252 8132 2258 8134
rect 1950 8123 2258 8132
rect 1584 8084 1636 8090
rect 1584 8026 1636 8032
rect 1122 7440 1178 7449
rect 1122 7375 1178 7384
rect 1950 7100 2258 7109
rect 1950 7098 1956 7100
rect 2012 7098 2036 7100
rect 2092 7098 2116 7100
rect 2172 7098 2196 7100
rect 2252 7098 2258 7100
rect 2012 7046 2014 7098
rect 2194 7046 2196 7098
rect 1950 7044 1956 7046
rect 2012 7044 2036 7046
rect 2092 7044 2116 7046
rect 2172 7044 2196 7046
rect 2252 7044 2258 7046
rect 1950 7035 2258 7044
rect 1950 6012 2258 6021
rect 1950 6010 1956 6012
rect 2012 6010 2036 6012
rect 2092 6010 2116 6012
rect 2172 6010 2196 6012
rect 2252 6010 2258 6012
rect 2012 5958 2014 6010
rect 2194 5958 2196 6010
rect 1950 5956 1956 5958
rect 2012 5956 2036 5958
rect 2092 5956 2116 5958
rect 2172 5956 2196 5958
rect 2252 5956 2258 5958
rect 1950 5947 2258 5956
rect 1950 4924 2258 4933
rect 1950 4922 1956 4924
rect 2012 4922 2036 4924
rect 2092 4922 2116 4924
rect 2172 4922 2196 4924
rect 2252 4922 2258 4924
rect 2012 4870 2014 4922
rect 2194 4870 2196 4922
rect 1950 4868 1956 4870
rect 2012 4868 2036 4870
rect 2092 4868 2116 4870
rect 2172 4868 2196 4870
rect 2252 4868 2258 4870
rect 1950 4859 2258 4868
rect 1950 3836 2258 3845
rect 1950 3834 1956 3836
rect 2012 3834 2036 3836
rect 2092 3834 2116 3836
rect 2172 3834 2196 3836
rect 2252 3834 2258 3836
rect 2012 3782 2014 3834
rect 2194 3782 2196 3834
rect 1950 3780 1956 3782
rect 2012 3780 2036 3782
rect 2092 3780 2116 3782
rect 2172 3780 2196 3782
rect 2252 3780 2258 3782
rect 1950 3771 2258 3780
rect 2332 3466 2360 8434
rect 2412 7880 2464 7886
rect 2410 7848 2412 7857
rect 2464 7848 2466 7857
rect 2410 7783 2466 7792
rect 2608 3942 2636 8434
rect 3804 8090 3832 11194
rect 4172 8634 4200 11194
rect 4344 9308 4396 9314
rect 4344 9250 4396 9256
rect 4160 8628 4212 8634
rect 4160 8570 4212 8576
rect 4356 8498 4384 9250
rect 4540 8634 4568 11194
rect 4712 8968 4764 8974
rect 4712 8910 4764 8916
rect 4618 8800 4674 8809
rect 4618 8735 4674 8744
rect 4528 8628 4580 8634
rect 4528 8570 4580 8576
rect 4344 8492 4396 8498
rect 4344 8434 4396 8440
rect 3792 8084 3844 8090
rect 3792 8026 3844 8032
rect 4632 7993 4660 8735
rect 4724 8498 4752 8910
rect 4908 8634 4936 11194
rect 5170 9616 5226 9625
rect 5170 9551 5226 9560
rect 5080 8832 5132 8838
rect 5080 8774 5132 8780
rect 4896 8628 4948 8634
rect 4896 8570 4948 8576
rect 5092 8498 5120 8774
rect 4712 8492 4764 8498
rect 4712 8434 4764 8440
rect 5080 8492 5132 8498
rect 5080 8434 5132 8440
rect 4618 7984 4674 7993
rect 4618 7919 4674 7928
rect 5184 7886 5212 9551
rect 5276 8634 5304 11194
rect 5644 8634 5672 11194
rect 6012 8634 6040 11194
rect 6276 9240 6328 9246
rect 6276 9182 6328 9188
rect 6184 8900 6236 8906
rect 6184 8842 6236 8848
rect 6196 8634 6224 8842
rect 5264 8628 5316 8634
rect 5264 8570 5316 8576
rect 5632 8628 5684 8634
rect 5632 8570 5684 8576
rect 6000 8628 6052 8634
rect 6000 8570 6052 8576
rect 6184 8628 6236 8634
rect 6184 8570 6236 8576
rect 6288 8498 6316 9182
rect 6276 8492 6328 8498
rect 6276 8434 6328 8440
rect 6380 8090 6408 11194
rect 6748 8634 6776 11194
rect 7012 9104 7064 9110
rect 7012 9046 7064 9052
rect 6736 8628 6788 8634
rect 6736 8570 6788 8576
rect 6828 8492 6880 8498
rect 6880 8452 6960 8480
rect 6828 8434 6880 8440
rect 6828 8356 6880 8362
rect 6828 8298 6880 8304
rect 6368 8084 6420 8090
rect 6368 8026 6420 8032
rect 5356 8016 5408 8022
rect 5354 7984 5356 7993
rect 5408 7984 5410 7993
rect 5354 7919 5410 7928
rect 4160 7880 4212 7886
rect 4160 7822 4212 7828
rect 5172 7880 5224 7886
rect 5172 7822 5224 7828
rect 6736 7880 6788 7886
rect 6736 7822 6788 7828
rect 3010 7644 3318 7653
rect 3010 7642 3016 7644
rect 3072 7642 3096 7644
rect 3152 7642 3176 7644
rect 3232 7642 3256 7644
rect 3312 7642 3318 7644
rect 3072 7590 3074 7642
rect 3254 7590 3256 7642
rect 3010 7588 3016 7590
rect 3072 7588 3096 7590
rect 3152 7588 3176 7590
rect 3232 7588 3256 7590
rect 3312 7588 3318 7590
rect 3010 7579 3318 7588
rect 4172 7546 4200 7822
rect 4160 7540 4212 7546
rect 4160 7482 4212 7488
rect 6748 7342 6776 7822
rect 6736 7336 6788 7342
rect 5998 7304 6054 7313
rect 6736 7278 6788 7284
rect 5998 7239 6054 7248
rect 2778 6624 2834 6633
rect 2778 6559 2834 6568
rect 2686 5264 2742 5273
rect 2686 5199 2742 5208
rect 2700 5001 2728 5199
rect 2686 4992 2742 5001
rect 2686 4927 2742 4936
rect 2596 3936 2648 3942
rect 2596 3878 2648 3884
rect 2320 3460 2372 3466
rect 2320 3402 2372 3408
rect 1308 2848 1360 2854
rect 1308 2790 1360 2796
rect 1320 1465 1348 2790
rect 2792 2774 2820 6559
rect 3010 6556 3318 6565
rect 3010 6554 3016 6556
rect 3072 6554 3096 6556
rect 3152 6554 3176 6556
rect 3232 6554 3256 6556
rect 3312 6554 3318 6556
rect 3072 6502 3074 6554
rect 3254 6502 3256 6554
rect 3010 6500 3016 6502
rect 3072 6500 3096 6502
rect 3152 6500 3176 6502
rect 3232 6500 3256 6502
rect 3312 6500 3318 6502
rect 3010 6491 3318 6500
rect 5630 6216 5686 6225
rect 5630 6151 5686 6160
rect 3010 5468 3318 5477
rect 3010 5466 3016 5468
rect 3072 5466 3096 5468
rect 3152 5466 3176 5468
rect 3232 5466 3256 5468
rect 3312 5466 3318 5468
rect 3072 5414 3074 5466
rect 3254 5414 3256 5466
rect 3010 5412 3016 5414
rect 3072 5412 3096 5414
rect 3152 5412 3176 5414
rect 3232 5412 3256 5414
rect 3312 5412 3318 5414
rect 3010 5403 3318 5412
rect 3146 5264 3202 5273
rect 2884 5222 3146 5250
rect 2884 5137 2912 5222
rect 3146 5199 3202 5208
rect 2870 5128 2926 5137
rect 2870 5063 2926 5072
rect 3010 4380 3318 4389
rect 3010 4378 3016 4380
rect 3072 4378 3096 4380
rect 3152 4378 3176 4380
rect 3232 4378 3256 4380
rect 3312 4378 3318 4380
rect 3072 4326 3074 4378
rect 3254 4326 3256 4378
rect 3010 4324 3016 4326
rect 3072 4324 3096 4326
rect 3152 4324 3176 4326
rect 3232 4324 3256 4326
rect 3312 4324 3318 4326
rect 3010 4315 3318 4324
rect 3010 3292 3318 3301
rect 3010 3290 3016 3292
rect 3072 3290 3096 3292
rect 3152 3290 3176 3292
rect 3232 3290 3256 3292
rect 3312 3290 3318 3292
rect 3072 3238 3074 3290
rect 3254 3238 3256 3290
rect 3010 3236 3016 3238
rect 3072 3236 3096 3238
rect 3152 3236 3176 3238
rect 3232 3236 3256 3238
rect 3312 3236 3318 3238
rect 3010 3227 3318 3236
rect 1950 2748 2258 2757
rect 1950 2746 1956 2748
rect 2012 2746 2036 2748
rect 2092 2746 2116 2748
rect 2172 2746 2196 2748
rect 2252 2746 2258 2748
rect 2792 2746 2912 2774
rect 2012 2694 2014 2746
rect 2194 2694 2196 2746
rect 1950 2692 1956 2694
rect 2012 2692 2036 2694
rect 2092 2692 2116 2694
rect 2172 2692 2196 2694
rect 2252 2692 2258 2694
rect 1950 2683 2258 2692
rect 2884 2106 2912 2746
rect 5644 2310 5672 6151
rect 6012 5302 6040 7239
rect 6840 6118 6868 8298
rect 6828 6112 6880 6118
rect 6828 6054 6880 6060
rect 6000 5296 6052 5302
rect 6000 5238 6052 5244
rect 6932 3466 6960 8452
rect 7024 8294 7052 9046
rect 7116 8634 7144 11194
rect 7484 8634 7512 11194
rect 7656 9376 7708 9382
rect 7656 9318 7708 9324
rect 7668 8974 7696 9318
rect 7656 8968 7708 8974
rect 7656 8910 7708 8916
rect 7746 8936 7802 8945
rect 7746 8871 7802 8880
rect 7104 8628 7156 8634
rect 7104 8570 7156 8576
rect 7472 8628 7524 8634
rect 7472 8570 7524 8576
rect 7656 8492 7708 8498
rect 7656 8434 7708 8440
rect 7012 8288 7064 8294
rect 7012 8230 7064 8236
rect 7668 7274 7696 8434
rect 7760 7478 7788 8871
rect 7852 8634 7880 11194
rect 8220 8634 8248 11194
rect 8484 9036 8536 9042
rect 8484 8978 8536 8984
rect 7840 8628 7892 8634
rect 7840 8570 7892 8576
rect 8208 8628 8260 8634
rect 8208 8570 8260 8576
rect 7840 8492 7892 8498
rect 7840 8434 7892 8440
rect 8392 8492 8444 8498
rect 8392 8434 8444 8440
rect 7748 7472 7800 7478
rect 7748 7414 7800 7420
rect 7656 7268 7708 7274
rect 7656 7210 7708 7216
rect 7852 6254 7880 8434
rect 8298 8392 8354 8401
rect 8298 8327 8354 8336
rect 7950 8188 8258 8197
rect 7950 8186 7956 8188
rect 8012 8186 8036 8188
rect 8092 8186 8116 8188
rect 8172 8186 8196 8188
rect 8252 8186 8258 8188
rect 8012 8134 8014 8186
rect 8194 8134 8196 8186
rect 7950 8132 7956 8134
rect 8012 8132 8036 8134
rect 8092 8132 8116 8134
rect 8172 8132 8196 8134
rect 8252 8132 8258 8134
rect 7950 8123 8258 8132
rect 8312 7478 8340 8327
rect 8300 7472 8352 7478
rect 8300 7414 8352 7420
rect 7950 7100 8258 7109
rect 7950 7098 7956 7100
rect 8012 7098 8036 7100
rect 8092 7098 8116 7100
rect 8172 7098 8196 7100
rect 8252 7098 8258 7100
rect 8012 7046 8014 7098
rect 8194 7046 8196 7098
rect 7950 7044 7956 7046
rect 8012 7044 8036 7046
rect 8092 7044 8116 7046
rect 8172 7044 8196 7046
rect 8252 7044 8258 7046
rect 7950 7035 8258 7044
rect 7840 6248 7892 6254
rect 7840 6190 7892 6196
rect 8404 6186 8432 8434
rect 8392 6180 8444 6186
rect 8392 6122 8444 6128
rect 7950 6012 8258 6021
rect 7950 6010 7956 6012
rect 8012 6010 8036 6012
rect 8092 6010 8116 6012
rect 8172 6010 8196 6012
rect 8252 6010 8258 6012
rect 8012 5958 8014 6010
rect 8194 5958 8196 6010
rect 7950 5956 7956 5958
rect 8012 5956 8036 5958
rect 8092 5956 8116 5958
rect 8172 5956 8196 5958
rect 8252 5956 8258 5958
rect 7950 5947 8258 5956
rect 7470 5264 7526 5273
rect 7470 5199 7526 5208
rect 7484 4729 7512 5199
rect 7950 4924 8258 4933
rect 7950 4922 7956 4924
rect 8012 4922 8036 4924
rect 8092 4922 8116 4924
rect 8172 4922 8196 4924
rect 8252 4922 8258 4924
rect 8012 4870 8014 4922
rect 8194 4870 8196 4922
rect 7950 4868 7956 4870
rect 8012 4868 8036 4870
rect 8092 4868 8116 4870
rect 8172 4868 8196 4870
rect 8252 4868 8258 4870
rect 7950 4859 8258 4868
rect 7470 4720 7526 4729
rect 7470 4655 7526 4664
rect 8496 4554 8524 8978
rect 8588 8634 8616 11194
rect 8760 9376 8812 9382
rect 8760 9318 8812 9324
rect 8668 8832 8720 8838
rect 8668 8774 8720 8780
rect 8576 8628 8628 8634
rect 8576 8570 8628 8576
rect 8680 4758 8708 8774
rect 8772 8498 8800 9318
rect 8956 8786 8984 11194
rect 9324 8922 9352 11194
rect 9324 8894 9444 8922
rect 8864 8758 8984 8786
rect 8760 8492 8812 8498
rect 8760 8434 8812 8440
rect 8864 8090 8892 8758
rect 9010 8732 9318 8741
rect 9010 8730 9016 8732
rect 9072 8730 9096 8732
rect 9152 8730 9176 8732
rect 9232 8730 9256 8732
rect 9312 8730 9318 8732
rect 9072 8678 9074 8730
rect 9254 8678 9256 8730
rect 9010 8676 9016 8678
rect 9072 8676 9096 8678
rect 9152 8676 9176 8678
rect 9232 8676 9256 8678
rect 9312 8676 9318 8678
rect 9010 8667 9318 8676
rect 9416 8634 9444 8894
rect 9692 8634 9720 11194
rect 10060 8634 10088 11194
rect 10232 8832 10284 8838
rect 10232 8774 10284 8780
rect 9404 8628 9456 8634
rect 9404 8570 9456 8576
rect 9680 8628 9732 8634
rect 9680 8570 9732 8576
rect 10048 8628 10100 8634
rect 10048 8570 10100 8576
rect 10244 8498 10272 8774
rect 10428 8634 10456 11194
rect 10796 8634 10824 11194
rect 10874 10976 10930 10985
rect 10874 10911 10930 10920
rect 10416 8628 10468 8634
rect 10416 8570 10468 8576
rect 10784 8628 10836 8634
rect 10784 8570 10836 8576
rect 9496 8492 9548 8498
rect 9496 8434 9548 8440
rect 9864 8492 9916 8498
rect 9864 8434 9916 8440
rect 10232 8492 10284 8498
rect 10232 8434 10284 8440
rect 8852 8084 8904 8090
rect 8852 8026 8904 8032
rect 9010 7644 9318 7653
rect 9010 7642 9016 7644
rect 9072 7642 9096 7644
rect 9152 7642 9176 7644
rect 9232 7642 9256 7644
rect 9312 7642 9318 7644
rect 9072 7590 9074 7642
rect 9254 7590 9256 7642
rect 9010 7588 9016 7590
rect 9072 7588 9096 7590
rect 9152 7588 9176 7590
rect 9232 7588 9256 7590
rect 9312 7588 9318 7590
rect 9010 7579 9318 7588
rect 9010 6556 9318 6565
rect 9010 6554 9016 6556
rect 9072 6554 9096 6556
rect 9152 6554 9176 6556
rect 9232 6554 9256 6556
rect 9312 6554 9318 6556
rect 9072 6502 9074 6554
rect 9254 6502 9256 6554
rect 9010 6500 9016 6502
rect 9072 6500 9096 6502
rect 9152 6500 9176 6502
rect 9232 6500 9256 6502
rect 9312 6500 9318 6502
rect 9010 6491 9318 6500
rect 9508 6089 9536 8434
rect 9588 7880 9640 7886
rect 9588 7822 9640 7828
rect 9494 6080 9550 6089
rect 9494 6015 9550 6024
rect 9600 5658 9628 7822
rect 9876 6769 9904 8434
rect 10888 8090 10916 10911
rect 11164 8634 11192 11194
rect 11152 8628 11204 8634
rect 11152 8570 11204 8576
rect 11244 8560 11296 8566
rect 11244 8502 11296 8508
rect 11428 8560 11480 8566
rect 11428 8502 11480 8508
rect 10968 8492 11020 8498
rect 10968 8434 11020 8440
rect 10876 8084 10928 8090
rect 10876 8026 10928 8032
rect 9862 6760 9918 6769
rect 9862 6695 9918 6704
rect 10980 6390 11008 8434
rect 11152 8356 11204 8362
rect 11152 8298 11204 8304
rect 11164 7721 11192 8298
rect 11150 7712 11206 7721
rect 11150 7647 11206 7656
rect 11256 7206 11284 8502
rect 11440 8090 11468 8502
rect 11532 8090 11560 11194
rect 11796 11008 11848 11014
rect 11796 10950 11848 10956
rect 11428 8084 11480 8090
rect 11428 8026 11480 8032
rect 11520 8084 11572 8090
rect 11520 8026 11572 8032
rect 11808 7886 11836 10950
rect 11900 8634 11928 11194
rect 11978 10840 12034 10849
rect 11978 10775 12034 10784
rect 11888 8628 11940 8634
rect 11888 8570 11940 8576
rect 11992 7886 12020 10775
rect 12268 8634 12296 11194
rect 12636 8634 12664 11194
rect 13004 8634 13032 11194
rect 13372 8634 13400 11194
rect 13726 11194 13782 11250
rect 14094 11194 14150 11250
rect 14462 11194 14518 11250
rect 14830 11194 14886 11250
rect 15198 11194 15254 11250
rect 15566 11194 15622 11250
rect 15934 11194 15990 11250
rect 16302 11194 16358 11250
rect 16670 11194 16726 11250
rect 17038 11194 17094 11250
rect 17406 11194 17462 11250
rect 17774 11194 17830 11250
rect 18142 11194 18198 11250
rect 18510 11194 18566 11250
rect 18878 11194 18934 11250
rect 19246 11194 19302 11250
rect 19614 11194 19670 11250
rect 19982 11194 20038 11250
rect 20350 11194 20406 11250
rect 20718 11194 20774 11250
rect 21086 11194 21142 11250
rect 21454 11194 21510 11250
rect 21822 11194 21878 11250
rect 22190 11194 22246 11250
rect 22558 11194 22614 11250
rect 22926 11194 22982 11250
rect 23294 11194 23350 11250
rect 23662 11194 23718 11250
rect 24030 11194 24086 11250
rect 24398 11194 24454 11250
rect 24766 11194 24822 11250
rect 25134 11194 25190 11250
rect 25502 11194 25558 11250
rect 25870 11194 25926 11250
rect 26238 11194 26294 11250
rect 26606 11194 26662 11250
rect 26974 11194 27030 11250
rect 27342 11194 27398 11250
rect 27710 11194 27766 11250
rect 28078 11194 28134 11250
rect 28446 11194 28502 11250
rect 28814 11194 28870 11250
rect 29182 11194 29238 11250
rect 29550 11194 29606 11250
rect 29918 11194 29974 11250
rect 30286 11194 30342 11250
rect 30654 11194 30710 11250
rect 31022 11194 31078 11250
rect 31390 11194 31446 11250
rect 31758 11194 31814 11250
rect 32126 11194 32182 11250
rect 32494 11194 32550 11250
rect 32862 11194 32918 11250
rect 33230 11194 33286 11250
rect 33598 11194 33654 11250
rect 33966 11194 34022 11250
rect 34334 11194 34390 11250
rect 34702 11194 34758 11250
rect 35070 11194 35126 11250
rect 35438 11194 35494 11250
rect 35806 11194 35862 11250
rect 36174 11194 36230 11250
rect 36542 11194 36598 11250
rect 36910 11194 36966 11250
rect 37278 11194 37334 11250
rect 37646 11194 37702 11250
rect 38014 11194 38070 11250
rect 38382 11194 38438 11250
rect 38750 11194 38806 11250
rect 39118 11194 39174 11250
rect 39486 11212 39542 11250
rect 39486 11194 39488 11212
rect 13544 11154 13596 11160
rect 12256 8628 12308 8634
rect 12256 8570 12308 8576
rect 12624 8628 12676 8634
rect 12624 8570 12676 8576
rect 12992 8628 13044 8634
rect 12992 8570 13044 8576
rect 13360 8628 13412 8634
rect 13360 8570 13412 8576
rect 12716 8492 12768 8498
rect 12716 8434 12768 8440
rect 13176 8492 13228 8498
rect 13176 8434 13228 8440
rect 12624 8424 12676 8430
rect 12624 8366 12676 8372
rect 12440 8356 12492 8362
rect 12440 8298 12492 8304
rect 12452 8265 12480 8298
rect 12438 8256 12494 8265
rect 12438 8191 12494 8200
rect 12440 8084 12492 8090
rect 12440 8026 12492 8032
rect 12452 7954 12480 8026
rect 12440 7948 12492 7954
rect 12440 7890 12492 7896
rect 11796 7880 11848 7886
rect 11796 7822 11848 7828
rect 11980 7880 12032 7886
rect 11980 7822 12032 7828
rect 12532 7880 12584 7886
rect 12532 7822 12584 7828
rect 11244 7200 11296 7206
rect 11244 7142 11296 7148
rect 12544 7002 12572 7822
rect 12532 6996 12584 7002
rect 12532 6938 12584 6944
rect 10968 6384 11020 6390
rect 10968 6326 11020 6332
rect 11058 6352 11114 6361
rect 11058 6287 11114 6296
rect 11072 5914 11100 6287
rect 11060 5908 11112 5914
rect 11060 5850 11112 5856
rect 12636 5846 12664 8366
rect 12728 6458 12756 8434
rect 12806 8256 12862 8265
rect 12806 8191 12862 8200
rect 12716 6452 12768 6458
rect 12716 6394 12768 6400
rect 12624 5840 12676 5846
rect 12624 5782 12676 5788
rect 12820 5778 12848 8191
rect 12992 8084 13044 8090
rect 12992 8026 13044 8032
rect 12808 5772 12860 5778
rect 12808 5714 12860 5720
rect 9600 5630 9720 5658
rect 9010 5468 9318 5477
rect 9010 5466 9016 5468
rect 9072 5466 9096 5468
rect 9152 5466 9176 5468
rect 9232 5466 9256 5468
rect 9312 5466 9318 5468
rect 9072 5414 9074 5466
rect 9254 5414 9256 5466
rect 9010 5412 9016 5414
rect 9072 5412 9096 5414
rect 9152 5412 9176 5414
rect 9232 5412 9256 5414
rect 9312 5412 9318 5414
rect 9010 5403 9318 5412
rect 9692 5409 9720 5630
rect 9678 5400 9734 5409
rect 9678 5335 9734 5344
rect 9586 5264 9642 5273
rect 9586 5199 9588 5208
rect 9640 5199 9642 5208
rect 9588 5170 9640 5176
rect 8668 4752 8720 4758
rect 8668 4694 8720 4700
rect 8484 4548 8536 4554
rect 8484 4490 8536 4496
rect 9010 4380 9318 4389
rect 9010 4378 9016 4380
rect 9072 4378 9096 4380
rect 9152 4378 9176 4380
rect 9232 4378 9256 4380
rect 9312 4378 9318 4380
rect 9072 4326 9074 4378
rect 9254 4326 9256 4378
rect 9010 4324 9016 4326
rect 9072 4324 9096 4326
rect 9152 4324 9176 4326
rect 9232 4324 9256 4326
rect 9312 4324 9318 4326
rect 9010 4315 9318 4324
rect 13004 4010 13032 8026
rect 13188 7954 13216 8434
rect 13176 7948 13228 7954
rect 13176 7890 13228 7896
rect 13556 7886 13584 11154
rect 13740 8634 13768 11194
rect 13728 8628 13780 8634
rect 13728 8570 13780 8576
rect 13636 8492 13688 8498
rect 13636 8434 13688 8440
rect 13728 8492 13780 8498
rect 13728 8434 13780 8440
rect 13648 8022 13676 8434
rect 13740 8090 13768 8434
rect 14108 8378 14136 11194
rect 14476 8634 14504 11194
rect 14556 9036 14608 9042
rect 14556 8978 14608 8984
rect 14464 8628 14516 8634
rect 14464 8570 14516 8576
rect 14464 8492 14516 8498
rect 14464 8434 14516 8440
rect 14108 8350 14320 8378
rect 13950 8188 14258 8197
rect 13950 8186 13956 8188
rect 14012 8186 14036 8188
rect 14092 8186 14116 8188
rect 14172 8186 14196 8188
rect 14252 8186 14258 8188
rect 14012 8134 14014 8186
rect 14194 8134 14196 8186
rect 13950 8132 13956 8134
rect 14012 8132 14036 8134
rect 14092 8132 14116 8134
rect 14172 8132 14196 8134
rect 14252 8132 14258 8134
rect 13950 8123 14258 8132
rect 14292 8090 14320 8350
rect 13728 8084 13780 8090
rect 13728 8026 13780 8032
rect 14280 8084 14332 8090
rect 14280 8026 14332 8032
rect 14476 8022 14504 8434
rect 13636 8016 13688 8022
rect 13636 7958 13688 7964
rect 14464 8016 14516 8022
rect 14464 7958 14516 7964
rect 14568 7886 14596 8978
rect 14648 8900 14700 8906
rect 14648 8842 14700 8848
rect 14660 8566 14688 8842
rect 14844 8634 14872 11194
rect 14924 11144 14976 11150
rect 14924 11086 14976 11092
rect 14832 8628 14884 8634
rect 14832 8570 14884 8576
rect 14648 8560 14700 8566
rect 14648 8502 14700 8508
rect 13544 7880 13596 7886
rect 13544 7822 13596 7828
rect 14556 7880 14608 7886
rect 14556 7822 14608 7828
rect 14280 7812 14332 7818
rect 14280 7754 14332 7760
rect 14292 7721 14320 7754
rect 14278 7712 14334 7721
rect 14278 7647 14334 7656
rect 13728 7540 13780 7546
rect 13728 7482 13780 7488
rect 13542 6896 13598 6905
rect 13542 6831 13598 6840
rect 13636 6860 13688 6866
rect 12992 4004 13044 4010
rect 12992 3946 13044 3952
rect 7950 3836 8258 3845
rect 7950 3834 7956 3836
rect 8012 3834 8036 3836
rect 8092 3834 8116 3836
rect 8172 3834 8196 3836
rect 8252 3834 8258 3836
rect 8012 3782 8014 3834
rect 8194 3782 8196 3834
rect 7950 3780 7956 3782
rect 8012 3780 8036 3782
rect 8092 3780 8116 3782
rect 8172 3780 8196 3782
rect 8252 3780 8258 3782
rect 7950 3771 8258 3780
rect 12808 3664 12860 3670
rect 12808 3606 12860 3612
rect 8852 3596 8904 3602
rect 8852 3538 8904 3544
rect 6920 3460 6972 3466
rect 6920 3402 6972 3408
rect 8864 3194 8892 3538
rect 9010 3292 9318 3301
rect 9010 3290 9016 3292
rect 9072 3290 9096 3292
rect 9152 3290 9176 3292
rect 9232 3290 9256 3292
rect 9312 3290 9318 3292
rect 9072 3238 9074 3290
rect 9254 3238 9256 3290
rect 9010 3236 9016 3238
rect 9072 3236 9096 3238
rect 9152 3236 9176 3238
rect 9232 3236 9256 3238
rect 9312 3236 9318 3238
rect 9010 3227 9318 3236
rect 9402 3224 9458 3233
rect 8852 3188 8904 3194
rect 12820 3194 12848 3606
rect 13556 3194 13584 6831
rect 13636 6802 13688 6808
rect 13648 4593 13676 6802
rect 13740 5370 13768 7482
rect 14936 7410 14964 11086
rect 15212 9738 15240 11194
rect 15212 9710 15424 9738
rect 15010 8732 15318 8741
rect 15010 8730 15016 8732
rect 15072 8730 15096 8732
rect 15152 8730 15176 8732
rect 15232 8730 15256 8732
rect 15312 8730 15318 8732
rect 15072 8678 15074 8730
rect 15254 8678 15256 8730
rect 15010 8676 15016 8678
rect 15072 8676 15096 8678
rect 15152 8676 15176 8678
rect 15232 8676 15256 8678
rect 15312 8676 15318 8678
rect 15010 8667 15318 8676
rect 15396 8634 15424 9710
rect 15476 9104 15528 9110
rect 15476 9046 15528 9052
rect 15488 8906 15516 9046
rect 15476 8900 15528 8906
rect 15476 8842 15528 8848
rect 15580 8634 15608 11194
rect 15660 9104 15712 9110
rect 15660 9046 15712 9052
rect 15384 8628 15436 8634
rect 15384 8570 15436 8576
rect 15568 8628 15620 8634
rect 15568 8570 15620 8576
rect 15108 8492 15160 8498
rect 15108 8434 15160 8440
rect 15476 8492 15528 8498
rect 15476 8434 15528 8440
rect 15120 8090 15148 8434
rect 15108 8084 15160 8090
rect 15108 8026 15160 8032
rect 15010 7644 15318 7653
rect 15010 7642 15016 7644
rect 15072 7642 15096 7644
rect 15152 7642 15176 7644
rect 15232 7642 15256 7644
rect 15312 7642 15318 7644
rect 15072 7590 15074 7642
rect 15254 7590 15256 7642
rect 15010 7588 15016 7590
rect 15072 7588 15096 7590
rect 15152 7588 15176 7590
rect 15232 7588 15256 7590
rect 15312 7588 15318 7590
rect 15010 7579 15318 7588
rect 15488 7546 15516 8434
rect 15568 7744 15620 7750
rect 15566 7712 15568 7721
rect 15620 7712 15622 7721
rect 15566 7647 15622 7656
rect 15476 7540 15528 7546
rect 15476 7482 15528 7488
rect 15672 7460 15700 9046
rect 15752 8900 15804 8906
rect 15752 8842 15804 8848
rect 15580 7432 15700 7460
rect 14924 7404 14976 7410
rect 14924 7346 14976 7352
rect 15476 7404 15528 7410
rect 15580 7392 15608 7432
rect 15528 7364 15608 7392
rect 15476 7346 15528 7352
rect 15384 7336 15436 7342
rect 15660 7336 15712 7342
rect 15436 7284 15660 7290
rect 15384 7278 15712 7284
rect 15396 7262 15700 7278
rect 14832 7200 14884 7206
rect 14832 7142 14884 7148
rect 13950 7100 14258 7109
rect 13950 7098 13956 7100
rect 14012 7098 14036 7100
rect 14092 7098 14116 7100
rect 14172 7098 14196 7100
rect 14252 7098 14258 7100
rect 14012 7046 14014 7098
rect 14194 7046 14196 7098
rect 13950 7044 13956 7046
rect 14012 7044 14036 7046
rect 14092 7044 14116 7046
rect 14172 7044 14196 7046
rect 14252 7044 14258 7046
rect 13950 7035 14258 7044
rect 14844 6934 14872 7142
rect 14832 6928 14884 6934
rect 14832 6870 14884 6876
rect 15010 6556 15318 6565
rect 15010 6554 15016 6556
rect 15072 6554 15096 6556
rect 15152 6554 15176 6556
rect 15232 6554 15256 6556
rect 15312 6554 15318 6556
rect 15072 6502 15074 6554
rect 15254 6502 15256 6554
rect 15010 6500 15016 6502
rect 15072 6500 15096 6502
rect 15152 6500 15176 6502
rect 15232 6500 15256 6502
rect 15312 6500 15318 6502
rect 15010 6491 15318 6500
rect 13950 6012 14258 6021
rect 13950 6010 13956 6012
rect 14012 6010 14036 6012
rect 14092 6010 14116 6012
rect 14172 6010 14196 6012
rect 14252 6010 14258 6012
rect 14012 5958 14014 6010
rect 14194 5958 14196 6010
rect 13950 5956 13956 5958
rect 14012 5956 14036 5958
rect 14092 5956 14116 5958
rect 14172 5956 14196 5958
rect 14252 5956 14258 5958
rect 13950 5947 14258 5956
rect 14924 5704 14976 5710
rect 14922 5672 14924 5681
rect 14976 5672 14978 5681
rect 14922 5607 14978 5616
rect 15010 5468 15318 5477
rect 15010 5466 15016 5468
rect 15072 5466 15096 5468
rect 15152 5466 15176 5468
rect 15232 5466 15256 5468
rect 15312 5466 15318 5468
rect 15072 5414 15074 5466
rect 15254 5414 15256 5466
rect 15010 5412 15016 5414
rect 15072 5412 15096 5414
rect 15152 5412 15176 5414
rect 15232 5412 15256 5414
rect 15312 5412 15318 5414
rect 14830 5400 14886 5409
rect 15010 5403 15318 5412
rect 13728 5364 13780 5370
rect 14830 5335 14886 5344
rect 13728 5306 13780 5312
rect 14844 5137 14872 5335
rect 14830 5128 14886 5137
rect 14830 5063 14886 5072
rect 13950 4924 14258 4933
rect 13950 4922 13956 4924
rect 14012 4922 14036 4924
rect 14092 4922 14116 4924
rect 14172 4922 14196 4924
rect 14252 4922 14258 4924
rect 14012 4870 14014 4922
rect 14194 4870 14196 4922
rect 13950 4868 13956 4870
rect 14012 4868 14036 4870
rect 14092 4868 14116 4870
rect 14172 4868 14196 4870
rect 14252 4868 14258 4870
rect 13950 4859 14258 4868
rect 13634 4584 13690 4593
rect 13634 4519 13690 4528
rect 15010 4380 15318 4389
rect 15010 4378 15016 4380
rect 15072 4378 15096 4380
rect 15152 4378 15176 4380
rect 15232 4378 15256 4380
rect 15312 4378 15318 4380
rect 15072 4326 15074 4378
rect 15254 4326 15256 4378
rect 15010 4324 15016 4326
rect 15072 4324 15096 4326
rect 15152 4324 15176 4326
rect 15232 4324 15256 4326
rect 15312 4324 15318 4326
rect 15010 4315 15318 4324
rect 15764 3942 15792 8842
rect 15948 8634 15976 11194
rect 16026 10704 16082 10713
rect 16026 10639 16082 10648
rect 15936 8628 15988 8634
rect 15936 8570 15988 8576
rect 15844 8492 15896 8498
rect 15844 8434 15896 8440
rect 15856 7546 15884 8434
rect 15844 7540 15896 7546
rect 15844 7482 15896 7488
rect 16040 6798 16068 10639
rect 16316 8634 16344 11194
rect 16394 11112 16450 11121
rect 16394 11047 16450 11056
rect 16304 8628 16356 8634
rect 16304 8570 16356 8576
rect 16212 8492 16264 8498
rect 16212 8434 16264 8440
rect 16224 7546 16252 8434
rect 16304 7948 16356 7954
rect 16304 7890 16356 7896
rect 16212 7540 16264 7546
rect 16212 7482 16264 7488
rect 16316 7206 16344 7890
rect 16304 7200 16356 7206
rect 16304 7142 16356 7148
rect 16408 6798 16436 11047
rect 16488 8424 16540 8430
rect 16488 8366 16540 8372
rect 16500 7478 16528 8366
rect 16684 8090 16712 11194
rect 16856 9376 16908 9382
rect 16856 9318 16908 9324
rect 16672 8084 16724 8090
rect 16672 8026 16724 8032
rect 16764 7880 16816 7886
rect 16764 7822 16816 7828
rect 16488 7472 16540 7478
rect 16488 7414 16540 7420
rect 16578 7440 16634 7449
rect 16578 7375 16580 7384
rect 16632 7375 16634 7384
rect 16580 7346 16632 7352
rect 16028 6792 16080 6798
rect 16028 6734 16080 6740
rect 16396 6792 16448 6798
rect 16396 6734 16448 6740
rect 16776 6730 16804 7822
rect 16764 6724 16816 6730
rect 16764 6666 16816 6672
rect 16868 6322 16896 9318
rect 16948 8492 17000 8498
rect 16948 8434 17000 8440
rect 16960 7546 16988 8434
rect 17052 8090 17080 11194
rect 17420 8634 17448 11194
rect 17408 8628 17460 8634
rect 17408 8570 17460 8576
rect 17592 8492 17644 8498
rect 17592 8434 17644 8440
rect 17604 8090 17632 8434
rect 17788 8430 17816 11194
rect 18052 8628 18104 8634
rect 18156 8616 18184 11194
rect 18236 11076 18288 11082
rect 18236 11018 18288 11024
rect 18104 8588 18184 8616
rect 18052 8570 18104 8576
rect 17960 8492 18012 8498
rect 17960 8434 18012 8440
rect 18144 8492 18196 8498
rect 18144 8434 18196 8440
rect 17776 8424 17828 8430
rect 17776 8366 17828 8372
rect 17972 8090 18000 8434
rect 18052 8356 18104 8362
rect 18052 8298 18104 8304
rect 17040 8084 17092 8090
rect 17040 8026 17092 8032
rect 17592 8084 17644 8090
rect 17592 8026 17644 8032
rect 17960 8084 18012 8090
rect 17960 8026 18012 8032
rect 18064 8022 18092 8298
rect 18052 8016 18104 8022
rect 18052 7958 18104 7964
rect 17132 7880 17184 7886
rect 17132 7822 17184 7828
rect 16948 7540 17000 7546
rect 16948 7482 17000 7488
rect 17144 6662 17172 7822
rect 17868 7744 17920 7750
rect 17868 7686 17920 7692
rect 17776 6860 17828 6866
rect 17776 6802 17828 6808
rect 17224 6724 17276 6730
rect 17224 6666 17276 6672
rect 17132 6656 17184 6662
rect 17132 6598 17184 6604
rect 17236 6458 17264 6666
rect 17224 6452 17276 6458
rect 17224 6394 17276 6400
rect 16856 6316 16908 6322
rect 16856 6258 16908 6264
rect 17788 5914 17816 6802
rect 17776 5908 17828 5914
rect 17776 5850 17828 5856
rect 17408 5568 17460 5574
rect 17408 5510 17460 5516
rect 17420 5001 17448 5510
rect 17406 4992 17462 5001
rect 17406 4927 17462 4936
rect 17880 4729 17908 7686
rect 18156 6610 18184 8434
rect 18248 7886 18276 11018
rect 18328 10940 18380 10946
rect 18328 10882 18380 10888
rect 18340 7886 18368 10882
rect 18524 8634 18552 11194
rect 18512 8628 18564 8634
rect 18512 8570 18564 8576
rect 18892 8362 18920 11194
rect 19156 9240 19208 9246
rect 19156 9182 19208 9188
rect 18972 8832 19024 8838
rect 18972 8774 19024 8780
rect 18880 8356 18932 8362
rect 18880 8298 18932 8304
rect 18880 7948 18932 7954
rect 18880 7890 18932 7896
rect 18236 7880 18288 7886
rect 18236 7822 18288 7828
rect 18328 7880 18380 7886
rect 18328 7822 18380 7828
rect 18788 7744 18840 7750
rect 18788 7686 18840 7692
rect 18064 6582 18184 6610
rect 18064 4826 18092 6582
rect 18234 6352 18290 6361
rect 18234 6287 18290 6296
rect 18144 5092 18196 5098
rect 18144 5034 18196 5040
rect 18052 4820 18104 4826
rect 18052 4762 18104 4768
rect 17866 4720 17922 4729
rect 17224 4684 17276 4690
rect 17866 4655 17922 4664
rect 17224 4626 17276 4632
rect 15752 3936 15804 3942
rect 14830 3904 14886 3913
rect 15752 3878 15804 3884
rect 13950 3836 14258 3845
rect 14830 3839 14886 3848
rect 13950 3834 13956 3836
rect 14012 3834 14036 3836
rect 14092 3834 14116 3836
rect 14172 3834 14196 3836
rect 14252 3834 14258 3836
rect 14012 3782 14014 3834
rect 14194 3782 14196 3834
rect 13950 3780 13956 3782
rect 14012 3780 14036 3782
rect 14092 3780 14116 3782
rect 14172 3780 14196 3782
rect 14252 3780 14258 3782
rect 13950 3771 14258 3780
rect 14844 3233 14872 3839
rect 15010 3292 15318 3301
rect 15010 3290 15016 3292
rect 15072 3290 15096 3292
rect 15152 3290 15176 3292
rect 15232 3290 15256 3292
rect 15312 3290 15318 3292
rect 15072 3238 15074 3290
rect 15254 3238 15256 3290
rect 15010 3236 15016 3238
rect 15072 3236 15096 3238
rect 15152 3236 15176 3238
rect 15232 3236 15256 3238
rect 15312 3236 15318 3238
rect 14830 3224 14886 3233
rect 15010 3227 15318 3236
rect 9402 3159 9458 3168
rect 12808 3188 12860 3194
rect 8852 3130 8904 3136
rect 8300 3120 8352 3126
rect 8300 3062 8352 3068
rect 7950 2748 8258 2757
rect 7950 2746 7956 2748
rect 8012 2746 8036 2748
rect 8092 2746 8116 2748
rect 8172 2746 8196 2748
rect 8252 2746 8258 2748
rect 8012 2694 8014 2746
rect 8194 2694 8196 2746
rect 7950 2692 7956 2694
rect 8012 2692 8036 2694
rect 8092 2692 8116 2694
rect 8172 2692 8196 2694
rect 8252 2692 8258 2694
rect 7950 2683 8258 2692
rect 5632 2304 5684 2310
rect 5632 2246 5684 2252
rect 3010 2204 3318 2213
rect 3010 2202 3016 2204
rect 3072 2202 3096 2204
rect 3152 2202 3176 2204
rect 3232 2202 3256 2204
rect 3312 2202 3318 2204
rect 3072 2150 3074 2202
rect 3254 2150 3256 2202
rect 3010 2148 3016 2150
rect 3072 2148 3096 2150
rect 3152 2148 3176 2150
rect 3232 2148 3256 2150
rect 3312 2148 3318 2150
rect 3010 2139 3318 2148
rect 2872 2100 2924 2106
rect 2872 2042 2924 2048
rect 1306 1456 1362 1465
rect 1306 1391 1362 1400
rect 3700 196 3752 202
rect 3700 138 3752 144
rect 6000 196 6052 202
rect 6000 138 6052 144
rect 1412 66 1532 82
rect 1412 60 1544 66
rect 1412 56 1492 60
rect 1398 54 1492 56
rect 1398 0 1454 54
rect 3712 56 3740 138
rect 6012 56 6040 138
rect 8312 56 8340 3062
rect 9416 2961 9444 3159
rect 12808 3130 12860 3136
rect 13544 3188 13596 3194
rect 14830 3159 14886 3168
rect 13544 3130 13596 3136
rect 9588 3120 9640 3126
rect 17236 3097 17264 4626
rect 17958 4040 18014 4049
rect 17958 3975 17960 3984
rect 18012 3975 18014 3984
rect 17960 3946 18012 3952
rect 18156 3126 18184 5034
rect 18248 4622 18276 6287
rect 18800 5166 18828 7686
rect 18892 7478 18920 7890
rect 18984 7750 19012 8774
rect 18972 7744 19024 7750
rect 18972 7686 19024 7692
rect 18880 7472 18932 7478
rect 18880 7414 18932 7420
rect 19168 7410 19196 9182
rect 19260 8634 19288 11194
rect 19522 9752 19578 9761
rect 19522 9687 19578 9696
rect 19248 8628 19300 8634
rect 19248 8570 19300 8576
rect 19432 8560 19484 8566
rect 19432 8502 19484 8508
rect 19444 8090 19472 8502
rect 19432 8084 19484 8090
rect 19432 8026 19484 8032
rect 19156 7404 19208 7410
rect 19156 7346 19208 7352
rect 19340 6996 19392 7002
rect 19340 6938 19392 6944
rect 19352 5778 19380 6938
rect 19340 5772 19392 5778
rect 19340 5714 19392 5720
rect 18788 5160 18840 5166
rect 18788 5102 18840 5108
rect 18236 4616 18288 4622
rect 18236 4558 18288 4564
rect 19536 3942 19564 9687
rect 19628 8634 19656 11194
rect 19798 9208 19854 9217
rect 19798 9143 19854 9152
rect 19708 8832 19760 8838
rect 19708 8774 19760 8780
rect 19720 8634 19748 8774
rect 19616 8628 19668 8634
rect 19616 8570 19668 8576
rect 19708 8628 19760 8634
rect 19708 8570 19760 8576
rect 19708 8356 19760 8362
rect 19708 8298 19760 8304
rect 19720 8090 19748 8298
rect 19708 8084 19760 8090
rect 19708 8026 19760 8032
rect 19812 7886 19840 9143
rect 19996 8634 20024 11194
rect 20260 9376 20312 9382
rect 20260 9318 20312 9324
rect 19984 8628 20036 8634
rect 19984 8570 20036 8576
rect 20272 8378 20300 9318
rect 20364 8634 20392 11194
rect 20732 9761 20760 11194
rect 20718 9752 20774 9761
rect 20718 9687 20774 9696
rect 20442 9344 20498 9353
rect 20442 9279 20498 9288
rect 20352 8628 20404 8634
rect 20352 8570 20404 8576
rect 20272 8350 20392 8378
rect 19950 8188 20258 8197
rect 19950 8186 19956 8188
rect 20012 8186 20036 8188
rect 20092 8186 20116 8188
rect 20172 8186 20196 8188
rect 20252 8186 20258 8188
rect 20012 8134 20014 8186
rect 20194 8134 20196 8186
rect 19950 8132 19956 8134
rect 20012 8132 20036 8134
rect 20092 8132 20116 8134
rect 20172 8132 20196 8134
rect 20252 8132 20258 8134
rect 19950 8123 20258 8132
rect 19800 7880 19852 7886
rect 19800 7822 19852 7828
rect 19950 7100 20258 7109
rect 19950 7098 19956 7100
rect 20012 7098 20036 7100
rect 20092 7098 20116 7100
rect 20172 7098 20196 7100
rect 20252 7098 20258 7100
rect 20012 7046 20014 7098
rect 20194 7046 20196 7098
rect 19950 7044 19956 7046
rect 20012 7044 20036 7046
rect 20092 7044 20116 7046
rect 20172 7044 20196 7046
rect 20252 7044 20258 7046
rect 19950 7035 20258 7044
rect 19950 6012 20258 6021
rect 19950 6010 19956 6012
rect 20012 6010 20036 6012
rect 20092 6010 20116 6012
rect 20172 6010 20196 6012
rect 20252 6010 20258 6012
rect 20012 5958 20014 6010
rect 20194 5958 20196 6010
rect 19950 5956 19956 5958
rect 20012 5956 20036 5958
rect 20092 5956 20116 5958
rect 20172 5956 20196 5958
rect 20252 5956 20258 5958
rect 19950 5947 20258 5956
rect 19798 5808 19854 5817
rect 19798 5743 19854 5752
rect 19812 4826 19840 5743
rect 20364 5030 20392 8350
rect 20456 7886 20484 9279
rect 21100 8922 21128 11194
rect 20916 8894 21128 8922
rect 20444 7880 20496 7886
rect 20444 7822 20496 7828
rect 20536 7880 20588 7886
rect 20536 7822 20588 7828
rect 20548 6497 20576 7822
rect 20626 7712 20682 7721
rect 20626 7647 20682 7656
rect 20640 7177 20668 7647
rect 20718 7576 20774 7585
rect 20718 7511 20774 7520
rect 20732 7410 20760 7511
rect 20720 7404 20772 7410
rect 20720 7346 20772 7352
rect 20626 7168 20682 7177
rect 20626 7103 20682 7112
rect 20534 6488 20590 6497
rect 20534 6423 20590 6432
rect 20352 5024 20404 5030
rect 20352 4966 20404 4972
rect 19950 4924 20258 4933
rect 19950 4922 19956 4924
rect 20012 4922 20036 4924
rect 20092 4922 20116 4924
rect 20172 4922 20196 4924
rect 20252 4922 20258 4924
rect 20012 4870 20014 4922
rect 20194 4870 20196 4922
rect 19950 4868 19956 4870
rect 20012 4868 20036 4870
rect 20092 4868 20116 4870
rect 20172 4868 20196 4870
rect 20252 4868 20258 4870
rect 19950 4859 20258 4868
rect 19800 4820 19852 4826
rect 19800 4762 19852 4768
rect 19524 3936 19576 3942
rect 19524 3878 19576 3884
rect 20720 3936 20772 3942
rect 20720 3878 20772 3884
rect 19950 3836 20258 3845
rect 19950 3834 19956 3836
rect 20012 3834 20036 3836
rect 20092 3834 20116 3836
rect 20172 3834 20196 3836
rect 20252 3834 20258 3836
rect 20012 3782 20014 3834
rect 20194 3782 20196 3834
rect 19950 3780 19956 3782
rect 20012 3780 20036 3782
rect 20092 3780 20116 3782
rect 20172 3780 20196 3782
rect 20252 3780 20258 3782
rect 19950 3771 20258 3780
rect 20732 3505 20760 3878
rect 20718 3496 20774 3505
rect 20718 3431 20774 3440
rect 20916 3398 20944 8894
rect 21010 8732 21318 8741
rect 21010 8730 21016 8732
rect 21072 8730 21096 8732
rect 21152 8730 21176 8732
rect 21232 8730 21256 8732
rect 21312 8730 21318 8732
rect 21072 8678 21074 8730
rect 21254 8678 21256 8730
rect 21010 8676 21016 8678
rect 21072 8676 21096 8678
rect 21152 8676 21176 8678
rect 21232 8676 21256 8678
rect 21312 8676 21318 8678
rect 21010 8667 21318 8676
rect 21364 8084 21416 8090
rect 21364 8026 21416 8032
rect 21376 7818 21404 8026
rect 21364 7812 21416 7818
rect 21364 7754 21416 7760
rect 21010 7644 21318 7653
rect 21010 7642 21016 7644
rect 21072 7642 21096 7644
rect 21152 7642 21176 7644
rect 21232 7642 21256 7644
rect 21312 7642 21318 7644
rect 21072 7590 21074 7642
rect 21254 7590 21256 7642
rect 21010 7588 21016 7590
rect 21072 7588 21096 7590
rect 21152 7588 21176 7590
rect 21232 7588 21256 7590
rect 21312 7588 21318 7590
rect 21010 7579 21318 7588
rect 21010 6556 21318 6565
rect 21010 6554 21016 6556
rect 21072 6554 21096 6556
rect 21152 6554 21176 6556
rect 21232 6554 21256 6556
rect 21312 6554 21318 6556
rect 21072 6502 21074 6554
rect 21254 6502 21256 6554
rect 21010 6500 21016 6502
rect 21072 6500 21096 6502
rect 21152 6500 21176 6502
rect 21232 6500 21256 6502
rect 21312 6500 21318 6502
rect 21010 6491 21318 6500
rect 21010 5468 21318 5477
rect 21010 5466 21016 5468
rect 21072 5466 21096 5468
rect 21152 5466 21176 5468
rect 21232 5466 21256 5468
rect 21312 5466 21318 5468
rect 21072 5414 21074 5466
rect 21254 5414 21256 5466
rect 21010 5412 21016 5414
rect 21072 5412 21096 5414
rect 21152 5412 21176 5414
rect 21232 5412 21256 5414
rect 21312 5412 21318 5414
rect 21010 5403 21318 5412
rect 21010 4380 21318 4389
rect 21010 4378 21016 4380
rect 21072 4378 21096 4380
rect 21152 4378 21176 4380
rect 21232 4378 21256 4380
rect 21312 4378 21318 4380
rect 21072 4326 21074 4378
rect 21254 4326 21256 4378
rect 21010 4324 21016 4326
rect 21072 4324 21096 4326
rect 21152 4324 21176 4326
rect 21232 4324 21256 4326
rect 21312 4324 21318 4326
rect 21010 4315 21318 4324
rect 21468 4146 21496 11194
rect 21640 7880 21692 7886
rect 21640 7822 21692 7828
rect 21652 7750 21680 7822
rect 21640 7744 21692 7750
rect 21640 7686 21692 7692
rect 21732 7744 21784 7750
rect 21732 7686 21784 7692
rect 21744 5098 21772 7686
rect 21732 5092 21784 5098
rect 21732 5034 21784 5040
rect 21456 4140 21508 4146
rect 21456 4082 21508 4088
rect 21836 4078 21864 11194
rect 21916 10736 21968 10742
rect 21916 10678 21968 10684
rect 21928 5234 21956 10678
rect 22204 6361 22232 11194
rect 22190 6352 22246 6361
rect 22190 6287 22246 6296
rect 22468 6112 22520 6118
rect 22468 6054 22520 6060
rect 22480 5914 22508 6054
rect 22468 5908 22520 5914
rect 22468 5850 22520 5856
rect 21916 5228 21968 5234
rect 21916 5170 21968 5176
rect 21824 4072 21876 4078
rect 21824 4014 21876 4020
rect 22100 3528 22152 3534
rect 22100 3470 22152 3476
rect 20904 3392 20956 3398
rect 20904 3334 20956 3340
rect 21010 3292 21318 3301
rect 21010 3290 21016 3292
rect 21072 3290 21096 3292
rect 21152 3290 21176 3292
rect 21232 3290 21256 3292
rect 21312 3290 21318 3292
rect 21072 3238 21074 3290
rect 21254 3238 21256 3290
rect 21010 3236 21016 3238
rect 21072 3236 21096 3238
rect 21152 3236 21176 3238
rect 21232 3236 21256 3238
rect 21312 3236 21318 3238
rect 21010 3227 21318 3236
rect 18144 3120 18196 3126
rect 9588 3062 9640 3068
rect 17222 3088 17278 3097
rect 9402 2952 9458 2961
rect 8576 2916 8628 2922
rect 9402 2887 9458 2896
rect 9496 2916 9548 2922
rect 8576 2858 8628 2864
rect 9496 2858 9548 2864
rect 8588 2446 8616 2858
rect 9508 2553 9536 2858
rect 9494 2544 9550 2553
rect 9494 2479 9550 2488
rect 8576 2440 8628 2446
rect 8576 2382 8628 2388
rect 9010 2204 9318 2213
rect 9010 2202 9016 2204
rect 9072 2202 9096 2204
rect 9152 2202 9176 2204
rect 9232 2202 9256 2204
rect 9312 2202 9318 2204
rect 9072 2150 9074 2202
rect 9254 2150 9256 2202
rect 9010 2148 9016 2150
rect 9072 2148 9096 2150
rect 9152 2148 9176 2150
rect 9232 2148 9256 2150
rect 9312 2148 9318 2150
rect 9010 2139 9318 2148
rect 9600 1737 9628 3062
rect 10600 3052 10652 3058
rect 10600 2994 10652 3000
rect 12900 3052 12952 3058
rect 12900 2994 12952 3000
rect 15384 3052 15436 3058
rect 18144 3062 18196 3068
rect 19800 3120 19852 3126
rect 19800 3062 19852 3068
rect 17222 3023 17278 3032
rect 15384 2994 15436 3000
rect 9586 1728 9642 1737
rect 9586 1663 9642 1672
rect 10612 56 10640 2994
rect 11060 2984 11112 2990
rect 11058 2952 11060 2961
rect 11112 2952 11114 2961
rect 11058 2887 11114 2896
rect 12912 56 12940 2994
rect 13268 2916 13320 2922
rect 13268 2858 13320 2864
rect 13280 2514 13308 2858
rect 13950 2748 14258 2757
rect 13950 2746 13956 2748
rect 14012 2746 14036 2748
rect 14092 2746 14116 2748
rect 14172 2746 14196 2748
rect 14252 2746 14258 2748
rect 14012 2694 14014 2746
rect 14194 2694 14196 2746
rect 13950 2692 13956 2694
rect 14012 2692 14036 2694
rect 14092 2692 14116 2694
rect 14172 2692 14196 2694
rect 14252 2692 14258 2694
rect 13950 2683 14258 2692
rect 13268 2508 13320 2514
rect 13268 2450 13320 2456
rect 15010 2204 15318 2213
rect 15010 2202 15016 2204
rect 15072 2202 15096 2204
rect 15152 2202 15176 2204
rect 15232 2202 15256 2204
rect 15312 2202 15318 2204
rect 15072 2150 15074 2202
rect 15254 2150 15256 2202
rect 15010 2148 15016 2150
rect 15072 2148 15096 2150
rect 15152 2148 15176 2150
rect 15232 2148 15256 2150
rect 15312 2148 15318 2150
rect 15010 2139 15318 2148
rect 15212 56 15332 82
rect 1492 2 1544 8
rect 3698 0 3754 56
rect 5998 0 6054 56
rect 8298 0 8354 56
rect 10598 0 10654 56
rect 12898 0 12954 56
rect 15198 54 15332 56
rect 15198 0 15254 54
rect 15304 42 15332 54
rect 15396 42 15424 2994
rect 17500 2984 17552 2990
rect 17500 2926 17552 2932
rect 16856 2848 16908 2854
rect 16856 2790 16908 2796
rect 16868 2582 16896 2790
rect 16856 2576 16908 2582
rect 16856 2518 16908 2524
rect 17512 56 17540 2926
rect 19708 2848 19760 2854
rect 19708 2790 19760 2796
rect 19720 2009 19748 2790
rect 19706 2000 19762 2009
rect 19706 1935 19762 1944
rect 19812 56 19840 3062
rect 20444 2848 20496 2854
rect 20444 2790 20496 2796
rect 20720 2848 20772 2854
rect 20720 2790 20772 2796
rect 21088 2848 21140 2854
rect 21088 2790 21140 2796
rect 19950 2748 20258 2757
rect 19950 2746 19956 2748
rect 20012 2746 20036 2748
rect 20092 2746 20116 2748
rect 20172 2746 20196 2748
rect 20252 2746 20258 2748
rect 20012 2694 20014 2746
rect 20194 2694 20196 2746
rect 19950 2692 19956 2694
rect 20012 2692 20036 2694
rect 20092 2692 20116 2694
rect 20172 2692 20196 2694
rect 20252 2692 20258 2694
rect 19950 2683 20258 2692
rect 20456 2650 20484 2790
rect 20444 2644 20496 2650
rect 20444 2586 20496 2592
rect 20732 2417 20760 2790
rect 20718 2408 20774 2417
rect 21100 2378 21128 2790
rect 20718 2343 20774 2352
rect 21088 2372 21140 2378
rect 21088 2314 21140 2320
rect 21010 2204 21318 2213
rect 21010 2202 21016 2204
rect 21072 2202 21096 2204
rect 21152 2202 21176 2204
rect 21232 2202 21256 2204
rect 21312 2202 21318 2204
rect 21072 2150 21074 2202
rect 21254 2150 21256 2202
rect 21010 2148 21016 2150
rect 21072 2148 21096 2150
rect 21152 2148 21176 2150
rect 21232 2148 21256 2150
rect 21312 2148 21318 2150
rect 21010 2139 21318 2148
rect 22112 56 22140 3470
rect 22572 3466 22600 11194
rect 22652 8084 22704 8090
rect 22652 8026 22704 8032
rect 22664 7750 22692 8026
rect 22652 7744 22704 7750
rect 22652 7686 22704 7692
rect 22742 7032 22798 7041
rect 22742 6967 22798 6976
rect 22560 3460 22612 3466
rect 22560 3402 22612 3408
rect 22756 3058 22784 6967
rect 22940 4690 22968 11194
rect 23308 7970 23336 11194
rect 23388 9172 23440 9178
rect 23388 9114 23440 9120
rect 23216 7942 23336 7970
rect 22928 4684 22980 4690
rect 22928 4626 22980 4632
rect 23112 4684 23164 4690
rect 23112 4626 23164 4632
rect 23020 3392 23072 3398
rect 23020 3334 23072 3340
rect 23032 3194 23060 3334
rect 23124 3194 23152 4626
rect 23216 4622 23244 7942
rect 23400 5370 23428 9114
rect 23676 8242 23704 11194
rect 24044 10742 24072 11194
rect 24032 10736 24084 10742
rect 24032 10678 24084 10684
rect 23584 8214 23704 8242
rect 23388 5364 23440 5370
rect 23388 5306 23440 5312
rect 23584 5302 23612 8214
rect 24124 8084 24176 8090
rect 24124 8026 24176 8032
rect 24136 7954 24164 8026
rect 24124 7948 24176 7954
rect 24124 7890 24176 7896
rect 23664 6656 23716 6662
rect 23664 6598 23716 6604
rect 23676 6458 23704 6598
rect 23664 6452 23716 6458
rect 23664 6394 23716 6400
rect 24412 5710 24440 11194
rect 24492 6316 24544 6322
rect 24492 6258 24544 6264
rect 24504 6118 24532 6258
rect 24492 6112 24544 6118
rect 24492 6054 24544 6060
rect 24676 6112 24728 6118
rect 24676 6054 24728 6060
rect 24400 5704 24452 5710
rect 24400 5646 24452 5652
rect 23572 5296 23624 5302
rect 23572 5238 23624 5244
rect 23204 4616 23256 4622
rect 23204 4558 23256 4564
rect 24688 4185 24716 6054
rect 24780 5234 24808 11194
rect 25148 6322 25176 11194
rect 25516 8786 25544 11194
rect 25780 9308 25832 9314
rect 25780 9250 25832 9256
rect 25516 8758 25636 8786
rect 25504 7472 25556 7478
rect 25504 7414 25556 7420
rect 25136 6316 25188 6322
rect 25136 6258 25188 6264
rect 24952 5636 25004 5642
rect 24952 5578 25004 5584
rect 24768 5228 24820 5234
rect 24768 5170 24820 5176
rect 24964 4826 24992 5578
rect 24952 4820 25004 4826
rect 24952 4762 25004 4768
rect 25516 4690 25544 7414
rect 25608 6322 25636 8758
rect 25792 7818 25820 9250
rect 25780 7812 25832 7818
rect 25780 7754 25832 7760
rect 25596 6316 25648 6322
rect 25596 6258 25648 6264
rect 25884 6254 25912 11194
rect 26252 9330 26280 11194
rect 26252 9302 26372 9330
rect 25950 8188 26258 8197
rect 25950 8186 25956 8188
rect 26012 8186 26036 8188
rect 26092 8186 26116 8188
rect 26172 8186 26196 8188
rect 26252 8186 26258 8188
rect 26012 8134 26014 8186
rect 26194 8134 26196 8186
rect 25950 8132 25956 8134
rect 26012 8132 26036 8134
rect 26092 8132 26116 8134
rect 26172 8132 26196 8134
rect 26252 8132 26258 8134
rect 25950 8123 26258 8132
rect 26344 7410 26372 9302
rect 26620 7886 26648 11194
rect 26988 9602 27016 11194
rect 26896 9574 27016 9602
rect 26792 9240 26844 9246
rect 26792 9182 26844 9188
rect 26804 8974 26832 9182
rect 26792 8968 26844 8974
rect 26792 8910 26844 8916
rect 26896 7886 26924 9574
rect 27010 8732 27318 8741
rect 27010 8730 27016 8732
rect 27072 8730 27096 8732
rect 27152 8730 27176 8732
rect 27232 8730 27256 8732
rect 27312 8730 27318 8732
rect 27072 8678 27074 8730
rect 27254 8678 27256 8730
rect 27010 8676 27016 8678
rect 27072 8676 27096 8678
rect 27152 8676 27176 8678
rect 27232 8676 27256 8678
rect 27312 8676 27318 8678
rect 27010 8667 27318 8676
rect 27356 7886 27384 11194
rect 27724 7954 27752 11194
rect 27712 7948 27764 7954
rect 27712 7890 27764 7896
rect 26608 7880 26660 7886
rect 26608 7822 26660 7828
rect 26884 7880 26936 7886
rect 26884 7822 26936 7828
rect 27344 7880 27396 7886
rect 27344 7822 27396 7828
rect 27010 7644 27318 7653
rect 27010 7642 27016 7644
rect 27072 7642 27096 7644
rect 27152 7642 27176 7644
rect 27232 7642 27256 7644
rect 27312 7642 27318 7644
rect 27072 7590 27074 7642
rect 27254 7590 27256 7642
rect 27010 7588 27016 7590
rect 27072 7588 27096 7590
rect 27152 7588 27176 7590
rect 27232 7588 27256 7590
rect 27312 7588 27318 7590
rect 27010 7579 27318 7588
rect 26332 7404 26384 7410
rect 26332 7346 26384 7352
rect 28092 7313 28120 11194
rect 28460 10849 28488 11194
rect 28828 10985 28856 11194
rect 29196 11014 29224 11194
rect 29184 11008 29236 11014
rect 28814 10976 28870 10985
rect 29184 10950 29236 10956
rect 28814 10911 28870 10920
rect 28446 10840 28502 10849
rect 28446 10775 28502 10784
rect 29092 8560 29144 8566
rect 29092 8502 29144 8508
rect 28264 7744 28316 7750
rect 28264 7686 28316 7692
rect 28276 7342 28304 7686
rect 28264 7336 28316 7342
rect 28078 7304 28134 7313
rect 28264 7278 28316 7284
rect 28078 7239 28134 7248
rect 25950 7100 26258 7109
rect 25950 7098 25956 7100
rect 26012 7098 26036 7100
rect 26092 7098 26116 7100
rect 26172 7098 26196 7100
rect 26252 7098 26258 7100
rect 26012 7046 26014 7098
rect 26194 7046 26196 7098
rect 25950 7044 25956 7046
rect 26012 7044 26036 7046
rect 26092 7044 26116 7046
rect 26172 7044 26196 7046
rect 26252 7044 26258 7046
rect 25950 7035 26258 7044
rect 27010 6556 27318 6565
rect 27010 6554 27016 6556
rect 27072 6554 27096 6556
rect 27152 6554 27176 6556
rect 27232 6554 27256 6556
rect 27312 6554 27318 6556
rect 27072 6502 27074 6554
rect 27254 6502 27256 6554
rect 27010 6500 27016 6502
rect 27072 6500 27096 6502
rect 27152 6500 27176 6502
rect 27232 6500 27256 6502
rect 27312 6500 27318 6502
rect 27010 6491 27318 6500
rect 25780 6248 25832 6254
rect 25780 6190 25832 6196
rect 25872 6248 25924 6254
rect 25872 6190 25924 6196
rect 26516 6248 26568 6254
rect 26516 6190 26568 6196
rect 25792 6066 25820 6190
rect 25872 6112 25924 6118
rect 25792 6060 25872 6066
rect 25792 6054 25924 6060
rect 25792 6038 25912 6054
rect 25950 6012 26258 6021
rect 25950 6010 25956 6012
rect 26012 6010 26036 6012
rect 26092 6010 26116 6012
rect 26172 6010 26196 6012
rect 26252 6010 26258 6012
rect 26012 5958 26014 6010
rect 26194 5958 26196 6010
rect 25950 5956 25956 5958
rect 26012 5956 26036 5958
rect 26092 5956 26116 5958
rect 26172 5956 26196 5958
rect 26252 5956 26258 5958
rect 25950 5947 26258 5956
rect 25950 4924 26258 4933
rect 25950 4922 25956 4924
rect 26012 4922 26036 4924
rect 26092 4922 26116 4924
rect 26172 4922 26196 4924
rect 26252 4922 26258 4924
rect 26012 4870 26014 4922
rect 26194 4870 26196 4922
rect 25950 4868 25956 4870
rect 26012 4868 26036 4870
rect 26092 4868 26116 4870
rect 26172 4868 26196 4870
rect 26252 4868 26258 4870
rect 25950 4859 26258 4868
rect 25504 4684 25556 4690
rect 25504 4626 25556 4632
rect 24860 4480 24912 4486
rect 24860 4422 24912 4428
rect 25228 4480 25280 4486
rect 25228 4422 25280 4428
rect 24674 4176 24730 4185
rect 24674 4111 24730 4120
rect 24766 4040 24822 4049
rect 24766 3975 24822 3984
rect 24780 3602 24808 3975
rect 24872 3641 24900 4422
rect 25240 4282 25268 4422
rect 25228 4276 25280 4282
rect 25228 4218 25280 4224
rect 25872 3936 25924 3942
rect 25872 3878 25924 3884
rect 24858 3632 24914 3641
rect 24768 3596 24820 3602
rect 24858 3567 24914 3576
rect 24768 3538 24820 3544
rect 25884 3505 25912 3878
rect 25950 3836 26258 3845
rect 25950 3834 25956 3836
rect 26012 3834 26036 3836
rect 26092 3834 26116 3836
rect 26172 3834 26196 3836
rect 26252 3834 26258 3836
rect 26012 3782 26014 3834
rect 26194 3782 26196 3834
rect 25950 3780 25956 3782
rect 26012 3780 26036 3782
rect 26092 3780 26116 3782
rect 26172 3780 26196 3782
rect 26252 3780 26258 3782
rect 25950 3771 26258 3780
rect 25870 3496 25926 3505
rect 25870 3431 25926 3440
rect 23020 3188 23072 3194
rect 23020 3130 23072 3136
rect 23112 3188 23164 3194
rect 23112 3130 23164 3136
rect 24400 3120 24452 3126
rect 24400 3062 24452 3068
rect 22744 3052 22796 3058
rect 22744 2994 22796 3000
rect 24412 56 24440 3062
rect 25320 3052 25372 3058
rect 25320 2994 25372 3000
rect 25332 2106 25360 2994
rect 26528 2854 26556 6190
rect 27620 5908 27672 5914
rect 27620 5850 27672 5856
rect 27010 5468 27318 5477
rect 27010 5466 27016 5468
rect 27072 5466 27096 5468
rect 27152 5466 27176 5468
rect 27232 5466 27256 5468
rect 27312 5466 27318 5468
rect 27072 5414 27074 5466
rect 27254 5414 27256 5466
rect 27010 5412 27016 5414
rect 27072 5412 27096 5414
rect 27152 5412 27176 5414
rect 27232 5412 27256 5414
rect 27312 5412 27318 5414
rect 27010 5403 27318 5412
rect 27632 5030 27660 5850
rect 27620 5024 27672 5030
rect 27620 4966 27672 4972
rect 27010 4380 27318 4389
rect 27010 4378 27016 4380
rect 27072 4378 27096 4380
rect 27152 4378 27176 4380
rect 27232 4378 27256 4380
rect 27312 4378 27318 4380
rect 27072 4326 27074 4378
rect 27254 4326 27256 4378
rect 27010 4324 27016 4326
rect 27072 4324 27096 4326
rect 27152 4324 27176 4326
rect 27232 4324 27256 4326
rect 27312 4324 27318 4326
rect 27010 4315 27318 4324
rect 28998 3632 29054 3641
rect 29104 3602 29132 8502
rect 29564 7954 29592 11194
rect 29552 7948 29604 7954
rect 29552 7890 29604 7896
rect 29932 7886 29960 11194
rect 30194 9072 30250 9081
rect 30194 9007 30250 9016
rect 30208 8090 30236 9007
rect 30196 8084 30248 8090
rect 30196 8026 30248 8032
rect 29920 7880 29972 7886
rect 29920 7822 29972 7828
rect 29828 7812 29880 7818
rect 29828 7754 29880 7760
rect 29840 7206 29868 7754
rect 29828 7200 29880 7206
rect 29828 7142 29880 7148
rect 30300 6798 30328 11194
rect 30564 7744 30616 7750
rect 30564 7686 30616 7692
rect 30576 7546 30604 7686
rect 30564 7540 30616 7546
rect 30564 7482 30616 7488
rect 30288 6792 30340 6798
rect 30288 6734 30340 6740
rect 29276 6656 29328 6662
rect 29276 6598 29328 6604
rect 29288 6390 29316 6598
rect 29276 6384 29328 6390
rect 29276 6326 29328 6332
rect 30668 5778 30696 11194
rect 30748 8424 30800 8430
rect 30748 8366 30800 8372
rect 30760 7818 30788 8366
rect 30748 7812 30800 7818
rect 30748 7754 30800 7760
rect 30656 5772 30708 5778
rect 30656 5714 30708 5720
rect 31036 5710 31064 11194
rect 31208 5908 31260 5914
rect 31208 5850 31260 5856
rect 31024 5704 31076 5710
rect 31024 5646 31076 5652
rect 31220 5642 31248 5850
rect 31404 5710 31432 11194
rect 31772 6798 31800 11194
rect 32140 9330 32168 11194
rect 32140 9302 32352 9330
rect 31950 8188 32258 8197
rect 31950 8186 31956 8188
rect 32012 8186 32036 8188
rect 32092 8186 32116 8188
rect 32172 8186 32196 8188
rect 32252 8186 32258 8188
rect 32012 8134 32014 8186
rect 32194 8134 32196 8186
rect 31950 8132 31956 8134
rect 32012 8132 32036 8134
rect 32092 8132 32116 8134
rect 32172 8132 32196 8134
rect 32252 8132 32258 8134
rect 31950 8123 32258 8132
rect 32324 7410 32352 9302
rect 32404 8900 32456 8906
rect 32404 8842 32456 8848
rect 32312 7404 32364 7410
rect 32312 7346 32364 7352
rect 31950 7100 32258 7109
rect 31950 7098 31956 7100
rect 32012 7098 32036 7100
rect 32092 7098 32116 7100
rect 32172 7098 32196 7100
rect 32252 7098 32258 7100
rect 32012 7046 32014 7098
rect 32194 7046 32196 7098
rect 31950 7044 31956 7046
rect 32012 7044 32036 7046
rect 32092 7044 32116 7046
rect 32172 7044 32196 7046
rect 32252 7044 32258 7046
rect 31950 7035 32258 7044
rect 31760 6792 31812 6798
rect 31760 6734 31812 6740
rect 32416 6322 32444 8842
rect 32508 7886 32536 11194
rect 32496 7880 32548 7886
rect 32496 7822 32548 7828
rect 32876 6798 32904 11194
rect 33244 8922 33272 11194
rect 33244 8894 33456 8922
rect 33010 8732 33318 8741
rect 33010 8730 33016 8732
rect 33072 8730 33096 8732
rect 33152 8730 33176 8732
rect 33232 8730 33256 8732
rect 33312 8730 33318 8732
rect 33072 8678 33074 8730
rect 33254 8678 33256 8730
rect 33010 8676 33016 8678
rect 33072 8676 33096 8678
rect 33152 8676 33176 8678
rect 33232 8676 33256 8678
rect 33312 8676 33318 8678
rect 33010 8667 33318 8676
rect 33010 7644 33318 7653
rect 33010 7642 33016 7644
rect 33072 7642 33096 7644
rect 33152 7642 33176 7644
rect 33232 7642 33256 7644
rect 33312 7642 33318 7644
rect 33072 7590 33074 7642
rect 33254 7590 33256 7642
rect 33010 7588 33016 7590
rect 33072 7588 33096 7590
rect 33152 7588 33176 7590
rect 33232 7588 33256 7590
rect 33312 7588 33318 7590
rect 33010 7579 33318 7588
rect 33324 7200 33376 7206
rect 33324 7142 33376 7148
rect 33336 6934 33364 7142
rect 33324 6928 33376 6934
rect 33324 6870 33376 6876
rect 32864 6792 32916 6798
rect 32864 6734 32916 6740
rect 32772 6724 32824 6730
rect 32772 6666 32824 6672
rect 32404 6316 32456 6322
rect 32404 6258 32456 6264
rect 31950 6012 32258 6021
rect 31950 6010 31956 6012
rect 32012 6010 32036 6012
rect 32092 6010 32116 6012
rect 32172 6010 32196 6012
rect 32252 6010 32258 6012
rect 32012 5958 32014 6010
rect 32194 5958 32196 6010
rect 31950 5956 31956 5958
rect 32012 5956 32036 5958
rect 32092 5956 32116 5958
rect 32172 5956 32196 5958
rect 32252 5956 32258 5958
rect 31950 5947 32258 5956
rect 31392 5704 31444 5710
rect 31392 5646 31444 5652
rect 31208 5636 31260 5642
rect 31208 5578 31260 5584
rect 32784 5273 32812 6666
rect 33010 6556 33318 6565
rect 33010 6554 33016 6556
rect 33072 6554 33096 6556
rect 33152 6554 33176 6556
rect 33232 6554 33256 6556
rect 33312 6554 33318 6556
rect 33072 6502 33074 6554
rect 33254 6502 33256 6554
rect 33010 6500 33016 6502
rect 33072 6500 33096 6502
rect 33152 6500 33176 6502
rect 33232 6500 33256 6502
rect 33312 6500 33318 6502
rect 33010 6491 33318 6500
rect 33428 6390 33456 8894
rect 33416 6384 33468 6390
rect 33416 6326 33468 6332
rect 33140 6112 33192 6118
rect 33140 6054 33192 6060
rect 33152 5778 33180 6054
rect 33140 5772 33192 5778
rect 33140 5714 33192 5720
rect 33010 5468 33318 5477
rect 33010 5466 33016 5468
rect 33072 5466 33096 5468
rect 33152 5466 33176 5468
rect 33232 5466 33256 5468
rect 33312 5466 33318 5468
rect 33072 5414 33074 5466
rect 33254 5414 33256 5466
rect 33010 5412 33016 5414
rect 33072 5412 33096 5414
rect 33152 5412 33176 5414
rect 33232 5412 33256 5414
rect 33312 5412 33318 5414
rect 33010 5403 33318 5412
rect 32770 5264 32826 5273
rect 33612 5234 33640 11194
rect 33980 5710 34008 11194
rect 34348 6322 34376 11194
rect 34426 9888 34482 9897
rect 34426 9823 34482 9832
rect 34440 9178 34468 9823
rect 34428 9172 34480 9178
rect 34428 9114 34480 9120
rect 34716 7954 34744 11194
rect 35084 8090 35112 11194
rect 35452 9353 35480 11194
rect 35438 9344 35494 9353
rect 35438 9279 35494 9288
rect 35820 9217 35848 11194
rect 36188 10946 36216 11194
rect 36556 11082 36584 11194
rect 36544 11076 36596 11082
rect 36544 11018 36596 11024
rect 36176 10940 36228 10946
rect 36176 10882 36228 10888
rect 35806 9208 35862 9217
rect 35806 9143 35862 9152
rect 36924 8974 36952 11194
rect 37292 11121 37320 11194
rect 37278 11112 37334 11121
rect 37278 11047 37334 11056
rect 37660 10713 37688 11194
rect 37646 10704 37702 10713
rect 37646 10639 37702 10648
rect 37278 9480 37334 9489
rect 37278 9415 37334 9424
rect 36912 8968 36964 8974
rect 36450 8936 36506 8945
rect 36912 8910 36964 8916
rect 36450 8871 36506 8880
rect 35808 8424 35860 8430
rect 35808 8366 35860 8372
rect 35072 8084 35124 8090
rect 35072 8026 35124 8032
rect 34704 7948 34756 7954
rect 34704 7890 34756 7896
rect 35346 6760 35402 6769
rect 35346 6695 35402 6704
rect 35360 6662 35388 6695
rect 35348 6656 35400 6662
rect 35348 6598 35400 6604
rect 34336 6316 34388 6322
rect 34336 6258 34388 6264
rect 34428 6180 34480 6186
rect 34428 6122 34480 6128
rect 33968 5704 34020 5710
rect 33968 5646 34020 5652
rect 32770 5199 32826 5208
rect 33600 5228 33652 5234
rect 33600 5170 33652 5176
rect 34440 5098 34468 6122
rect 34428 5092 34480 5098
rect 34428 5034 34480 5040
rect 31950 4924 32258 4933
rect 31950 4922 31956 4924
rect 32012 4922 32036 4924
rect 32092 4922 32116 4924
rect 32172 4922 32196 4924
rect 32252 4922 32258 4924
rect 32012 4870 32014 4922
rect 32194 4870 32196 4922
rect 31950 4868 31956 4870
rect 32012 4868 32036 4870
rect 32092 4868 32116 4870
rect 32172 4868 32196 4870
rect 32252 4868 32258 4870
rect 31950 4859 32258 4868
rect 33010 4380 33318 4389
rect 33010 4378 33016 4380
rect 33072 4378 33096 4380
rect 33152 4378 33176 4380
rect 33232 4378 33256 4380
rect 33312 4378 33318 4380
rect 33072 4326 33074 4378
rect 33254 4326 33256 4378
rect 33010 4324 33016 4326
rect 33072 4324 33096 4326
rect 33152 4324 33176 4326
rect 33232 4324 33256 4326
rect 33312 4324 33318 4326
rect 33010 4315 33318 4324
rect 31950 3836 32258 3845
rect 31950 3834 31956 3836
rect 32012 3834 32036 3836
rect 32092 3834 32116 3836
rect 32172 3834 32196 3836
rect 32252 3834 32258 3836
rect 32012 3782 32014 3834
rect 32194 3782 32196 3834
rect 31950 3780 31956 3782
rect 32012 3780 32036 3782
rect 32092 3780 32116 3782
rect 32172 3780 32196 3782
rect 32252 3780 32258 3782
rect 31950 3771 32258 3780
rect 28998 3567 29054 3576
rect 29092 3596 29144 3602
rect 27436 3460 27488 3466
rect 27436 3402 27488 3408
rect 27010 3292 27318 3301
rect 27010 3290 27016 3292
rect 27072 3290 27096 3292
rect 27152 3290 27176 3292
rect 27232 3290 27256 3292
rect 27312 3290 27318 3292
rect 27072 3238 27074 3290
rect 27254 3238 27256 3290
rect 27010 3236 27016 3238
rect 27072 3236 27096 3238
rect 27152 3236 27176 3238
rect 27232 3236 27256 3238
rect 27312 3236 27318 3238
rect 27010 3227 27318 3236
rect 26700 3188 26752 3194
rect 26700 3130 26752 3136
rect 26516 2848 26568 2854
rect 26516 2790 26568 2796
rect 25950 2748 26258 2757
rect 25950 2746 25956 2748
rect 26012 2746 26036 2748
rect 26092 2746 26116 2748
rect 26172 2746 26196 2748
rect 26252 2746 26258 2748
rect 26012 2694 26014 2746
rect 26194 2694 26196 2746
rect 25950 2692 25956 2694
rect 26012 2692 26036 2694
rect 26092 2692 26116 2694
rect 26172 2692 26196 2694
rect 26252 2692 26258 2694
rect 25950 2683 26258 2692
rect 25320 2100 25372 2106
rect 25320 2042 25372 2048
rect 26712 56 26740 3130
rect 27448 2854 27476 3402
rect 28540 3392 28592 3398
rect 28540 3334 28592 3340
rect 28552 3097 28580 3334
rect 28538 3088 28594 3097
rect 27528 3052 27580 3058
rect 28538 3023 28594 3032
rect 27528 2994 27580 3000
rect 27436 2848 27488 2854
rect 27436 2790 27488 2796
rect 27540 2310 27568 2994
rect 27528 2304 27580 2310
rect 27528 2246 27580 2252
rect 27010 2204 27318 2213
rect 27010 2202 27016 2204
rect 27072 2202 27096 2204
rect 27152 2202 27176 2204
rect 27232 2202 27256 2204
rect 27312 2202 27318 2204
rect 27072 2150 27074 2202
rect 27254 2150 27256 2202
rect 27010 2148 27016 2150
rect 27072 2148 27096 2150
rect 27152 2148 27176 2150
rect 27232 2148 27256 2150
rect 27312 2148 27318 2150
rect 27010 2139 27318 2148
rect 29012 56 29040 3567
rect 29092 3538 29144 3544
rect 29460 3528 29512 3534
rect 29460 3470 29512 3476
rect 29368 3188 29420 3194
rect 29368 3130 29420 3136
rect 29380 2854 29408 3130
rect 29472 3058 29500 3470
rect 33600 3392 33652 3398
rect 33600 3334 33652 3340
rect 33010 3292 33318 3301
rect 33010 3290 33016 3292
rect 33072 3290 33096 3292
rect 33152 3290 33176 3292
rect 33232 3290 33256 3292
rect 33312 3290 33318 3292
rect 33072 3238 33074 3290
rect 33254 3238 33256 3290
rect 33010 3236 33016 3238
rect 33072 3236 33096 3238
rect 33152 3236 33176 3238
rect 33232 3236 33256 3238
rect 33312 3236 33318 3238
rect 33010 3227 33318 3236
rect 32036 3188 32088 3194
rect 32036 3130 32088 3136
rect 29460 3052 29512 3058
rect 29460 2994 29512 3000
rect 31760 2984 31812 2990
rect 32048 2972 32076 3130
rect 31812 2944 32076 2972
rect 31760 2926 31812 2932
rect 29368 2848 29420 2854
rect 29368 2790 29420 2796
rect 31950 2748 32258 2757
rect 31950 2746 31956 2748
rect 32012 2746 32036 2748
rect 32092 2746 32116 2748
rect 32172 2746 32196 2748
rect 32252 2746 32258 2748
rect 32012 2694 32014 2746
rect 32194 2694 32196 2746
rect 31950 2692 31956 2694
rect 32012 2692 32036 2694
rect 32092 2692 32116 2694
rect 32172 2692 32196 2694
rect 32252 2692 32258 2694
rect 31950 2683 32258 2692
rect 33140 2508 33192 2514
rect 33140 2450 33192 2456
rect 33152 2378 33180 2450
rect 33140 2372 33192 2378
rect 33140 2314 33192 2320
rect 33010 2204 33318 2213
rect 33010 2202 33016 2204
rect 33072 2202 33096 2204
rect 33152 2202 33176 2204
rect 33232 2202 33256 2204
rect 33312 2202 33318 2204
rect 33072 2150 33074 2202
rect 33254 2150 33256 2202
rect 33010 2148 33016 2150
rect 33072 2148 33096 2150
rect 33152 2148 33176 2150
rect 33232 2148 33256 2150
rect 33312 2148 33318 2150
rect 33010 2139 33318 2148
rect 31300 2100 31352 2106
rect 31300 2042 31352 2048
rect 31312 56 31340 2042
rect 33612 56 33640 3334
rect 35820 2854 35848 8366
rect 35900 7472 35952 7478
rect 35900 7414 35952 7420
rect 35808 2848 35860 2854
rect 35808 2790 35860 2796
rect 35912 56 35940 7414
rect 36174 6216 36230 6225
rect 36174 6151 36176 6160
rect 36228 6151 36230 6160
rect 36268 6180 36320 6186
rect 36176 6122 36228 6128
rect 36268 6122 36320 6128
rect 36280 5846 36308 6122
rect 36268 5840 36320 5846
rect 36268 5782 36320 5788
rect 36464 3058 36492 8871
rect 37188 8492 37240 8498
rect 37188 8434 37240 8440
rect 36912 6996 36964 7002
rect 36912 6938 36964 6944
rect 36452 3052 36504 3058
rect 36452 2994 36504 3000
rect 36924 2854 36952 6938
rect 37200 5846 37228 8434
rect 37188 5840 37240 5846
rect 37188 5782 37240 5788
rect 37292 3058 37320 9415
rect 38028 9330 38056 11194
rect 37844 9302 38056 9330
rect 37844 7449 37872 9302
rect 38396 9110 38424 11194
rect 38764 11150 38792 11194
rect 38752 11144 38804 11150
rect 38752 11086 38804 11092
rect 38384 9104 38436 9110
rect 38384 9046 38436 9052
rect 39132 9042 39160 11194
rect 39540 11194 39542 11212
rect 39854 11194 39910 11250
rect 40222 11194 40278 11250
rect 40590 11194 40646 11250
rect 40958 11194 41014 11250
rect 41326 11194 41382 11250
rect 41694 11194 41750 11250
rect 42062 11194 42118 11250
rect 42430 11194 42486 11250
rect 42798 11194 42854 11250
rect 43166 11194 43222 11250
rect 43534 11194 43590 11250
rect 43902 11194 43958 11250
rect 44270 11194 44326 11250
rect 44638 11194 44694 11250
rect 45006 11194 45062 11250
rect 45374 11194 45430 11250
rect 45742 11194 45798 11250
rect 45848 11206 46060 11234
rect 39488 11154 39540 11160
rect 39120 9036 39172 9042
rect 39120 8978 39172 8984
rect 39010 8732 39318 8741
rect 39010 8730 39016 8732
rect 39072 8730 39096 8732
rect 39152 8730 39176 8732
rect 39232 8730 39256 8732
rect 39312 8730 39318 8732
rect 39072 8678 39074 8730
rect 39254 8678 39256 8730
rect 39010 8676 39016 8678
rect 39072 8676 39096 8678
rect 39152 8676 39176 8678
rect 39232 8676 39256 8678
rect 39312 8676 39318 8678
rect 39010 8667 39318 8676
rect 39868 8634 39896 11194
rect 40236 8634 40264 11194
rect 40500 8832 40552 8838
rect 40500 8774 40552 8780
rect 39856 8628 39908 8634
rect 39856 8570 39908 8576
rect 40224 8628 40276 8634
rect 40224 8570 40276 8576
rect 38752 8492 38804 8498
rect 38752 8434 38804 8440
rect 38568 8356 38620 8362
rect 38568 8298 38620 8304
rect 37950 8188 38258 8197
rect 37950 8186 37956 8188
rect 38012 8186 38036 8188
rect 38092 8186 38116 8188
rect 38172 8186 38196 8188
rect 38252 8186 38258 8188
rect 38012 8134 38014 8186
rect 38194 8134 38196 8186
rect 37950 8132 37956 8134
rect 38012 8132 38036 8134
rect 38092 8132 38116 8134
rect 38172 8132 38196 8134
rect 38252 8132 38258 8134
rect 37950 8123 38258 8132
rect 38292 7880 38344 7886
rect 38292 7822 38344 7828
rect 37830 7440 37886 7449
rect 37830 7375 37886 7384
rect 37950 7100 38258 7109
rect 37950 7098 37956 7100
rect 38012 7098 38036 7100
rect 38092 7098 38116 7100
rect 38172 7098 38196 7100
rect 38252 7098 38258 7100
rect 38012 7046 38014 7098
rect 38194 7046 38196 7098
rect 37950 7044 37956 7046
rect 38012 7044 38036 7046
rect 38092 7044 38116 7046
rect 38172 7044 38196 7046
rect 38252 7044 38258 7046
rect 37950 7035 38258 7044
rect 37950 6012 38258 6021
rect 37950 6010 37956 6012
rect 38012 6010 38036 6012
rect 38092 6010 38116 6012
rect 38172 6010 38196 6012
rect 38252 6010 38258 6012
rect 38012 5958 38014 6010
rect 38194 5958 38196 6010
rect 37950 5956 37956 5958
rect 38012 5956 38036 5958
rect 38092 5956 38116 5958
rect 38172 5956 38196 5958
rect 38252 5956 38258 5958
rect 37950 5947 38258 5956
rect 37556 5160 37608 5166
rect 37554 5128 37556 5137
rect 37608 5128 37610 5137
rect 37554 5063 37610 5072
rect 37950 4924 38258 4933
rect 37950 4922 37956 4924
rect 38012 4922 38036 4924
rect 38092 4922 38116 4924
rect 38172 4922 38196 4924
rect 38252 4922 38258 4924
rect 38012 4870 38014 4922
rect 38194 4870 38196 4922
rect 37950 4868 37956 4870
rect 38012 4868 38036 4870
rect 38092 4868 38116 4870
rect 38172 4868 38196 4870
rect 38252 4868 38258 4870
rect 37950 4859 38258 4868
rect 37648 3936 37700 3942
rect 37648 3878 37700 3884
rect 37280 3052 37332 3058
rect 37280 2994 37332 3000
rect 37660 2854 37688 3878
rect 37950 3836 38258 3845
rect 37950 3834 37956 3836
rect 38012 3834 38036 3836
rect 38092 3834 38116 3836
rect 38172 3834 38196 3836
rect 38252 3834 38258 3836
rect 38012 3782 38014 3834
rect 38194 3782 38196 3834
rect 37950 3780 37956 3782
rect 38012 3780 38036 3782
rect 38092 3780 38116 3782
rect 38172 3780 38196 3782
rect 38252 3780 38258 3782
rect 37950 3771 38258 3780
rect 37740 3188 37792 3194
rect 37740 3130 37792 3136
rect 37752 2854 37780 3130
rect 36912 2848 36964 2854
rect 36912 2790 36964 2796
rect 37648 2848 37700 2854
rect 37648 2790 37700 2796
rect 37740 2848 37792 2854
rect 37740 2790 37792 2796
rect 37950 2748 38258 2757
rect 37950 2746 37956 2748
rect 38012 2746 38036 2748
rect 38092 2746 38116 2748
rect 38172 2746 38196 2748
rect 38252 2746 38258 2748
rect 38012 2694 38014 2746
rect 38194 2694 38196 2746
rect 37950 2692 37956 2694
rect 38012 2692 38036 2694
rect 38092 2692 38116 2694
rect 38172 2692 38196 2694
rect 38252 2692 38258 2694
rect 37950 2683 38258 2692
rect 36268 2440 36320 2446
rect 36452 2440 36504 2446
rect 36320 2388 36452 2394
rect 36268 2382 36504 2388
rect 36280 2366 36492 2382
rect 38304 1442 38332 7822
rect 38580 6458 38608 8298
rect 38568 6452 38620 6458
rect 38568 6394 38620 6400
rect 38764 3194 38792 8434
rect 39672 8424 39724 8430
rect 39672 8366 39724 8372
rect 39580 7812 39632 7818
rect 39580 7754 39632 7760
rect 39010 7644 39318 7653
rect 39010 7642 39016 7644
rect 39072 7642 39096 7644
rect 39152 7642 39176 7644
rect 39232 7642 39256 7644
rect 39312 7642 39318 7644
rect 39072 7590 39074 7642
rect 39254 7590 39256 7642
rect 39010 7588 39016 7590
rect 39072 7588 39096 7590
rect 39152 7588 39176 7590
rect 39232 7588 39256 7590
rect 39312 7588 39318 7590
rect 39010 7579 39318 7588
rect 39592 7546 39620 7754
rect 39580 7540 39632 7546
rect 39580 7482 39632 7488
rect 39396 6860 39448 6866
rect 39396 6802 39448 6808
rect 39010 6556 39318 6565
rect 39010 6554 39016 6556
rect 39072 6554 39096 6556
rect 39152 6554 39176 6556
rect 39232 6554 39256 6556
rect 39312 6554 39318 6556
rect 39072 6502 39074 6554
rect 39254 6502 39256 6554
rect 39010 6500 39016 6502
rect 39072 6500 39096 6502
rect 39152 6500 39176 6502
rect 39232 6500 39256 6502
rect 39312 6500 39318 6502
rect 39010 6491 39318 6500
rect 39408 5710 39436 6802
rect 39396 5704 39448 5710
rect 39396 5646 39448 5652
rect 39010 5468 39318 5477
rect 39010 5466 39016 5468
rect 39072 5466 39096 5468
rect 39152 5466 39176 5468
rect 39232 5466 39256 5468
rect 39312 5466 39318 5468
rect 39072 5414 39074 5466
rect 39254 5414 39256 5466
rect 39010 5412 39016 5414
rect 39072 5412 39096 5414
rect 39152 5412 39176 5414
rect 39232 5412 39256 5414
rect 39312 5412 39318 5414
rect 39010 5403 39318 5412
rect 39010 4380 39318 4389
rect 39010 4378 39016 4380
rect 39072 4378 39096 4380
rect 39152 4378 39176 4380
rect 39232 4378 39256 4380
rect 39312 4378 39318 4380
rect 39072 4326 39074 4378
rect 39254 4326 39256 4378
rect 39010 4324 39016 4326
rect 39072 4324 39096 4326
rect 39152 4324 39176 4326
rect 39232 4324 39256 4326
rect 39312 4324 39318 4326
rect 39010 4315 39318 4324
rect 39010 3292 39318 3301
rect 39010 3290 39016 3292
rect 39072 3290 39096 3292
rect 39152 3290 39176 3292
rect 39232 3290 39256 3292
rect 39312 3290 39318 3292
rect 39072 3238 39074 3290
rect 39254 3238 39256 3290
rect 39010 3236 39016 3238
rect 39072 3236 39096 3238
rect 39152 3236 39176 3238
rect 39232 3236 39256 3238
rect 39312 3236 39318 3238
rect 39010 3227 39318 3236
rect 39684 3194 39712 8366
rect 39948 8288 40000 8294
rect 39948 8230 40000 8236
rect 39960 8022 39988 8230
rect 40512 8090 40540 8774
rect 40604 8634 40632 11194
rect 40776 8832 40828 8838
rect 40776 8774 40828 8780
rect 40592 8628 40644 8634
rect 40592 8570 40644 8576
rect 40684 8492 40736 8498
rect 40684 8434 40736 8440
rect 40500 8084 40552 8090
rect 40500 8026 40552 8032
rect 39948 8016 40000 8022
rect 39948 7958 40000 7964
rect 40500 7336 40552 7342
rect 40500 7278 40552 7284
rect 40040 6384 40092 6390
rect 40040 6326 40092 6332
rect 40052 4622 40080 6326
rect 40040 4616 40092 4622
rect 40040 4558 40092 4564
rect 38752 3188 38804 3194
rect 38752 3130 38804 3136
rect 39672 3188 39724 3194
rect 39672 3130 39724 3136
rect 38568 3052 38620 3058
rect 38568 2994 38620 3000
rect 39488 3052 39540 3058
rect 39488 2994 39540 3000
rect 40316 3052 40368 3058
rect 40316 2994 40368 3000
rect 38212 1414 38332 1442
rect 38212 56 38240 1414
rect 38580 66 38608 2994
rect 39010 2204 39318 2213
rect 39010 2202 39016 2204
rect 39072 2202 39096 2204
rect 39152 2202 39176 2204
rect 39232 2202 39256 2204
rect 39312 2202 39318 2204
rect 39072 2150 39074 2202
rect 39254 2150 39256 2202
rect 39010 2148 39016 2150
rect 39072 2148 39096 2150
rect 39152 2148 39176 2150
rect 39232 2148 39256 2150
rect 39312 2148 39318 2150
rect 39010 2139 39318 2148
rect 39500 134 39528 2994
rect 40328 202 40356 2994
rect 40316 196 40368 202
rect 40316 138 40368 144
rect 39488 128 39540 134
rect 39488 70 39540 76
rect 38568 60 38620 66
rect 15304 14 15424 42
rect 17498 0 17554 56
rect 19798 0 19854 56
rect 22098 0 22154 56
rect 24398 0 24454 56
rect 26698 0 26754 56
rect 28998 0 29054 56
rect 31298 0 31354 56
rect 33598 0 33654 56
rect 35898 0 35954 56
rect 38198 0 38254 56
rect 40512 56 40540 7278
rect 40696 3194 40724 8434
rect 40788 3466 40816 8774
rect 40972 8634 41000 11194
rect 41340 8634 41368 11194
rect 41708 8634 41736 11194
rect 42076 8634 42104 11194
rect 40960 8628 41012 8634
rect 40960 8570 41012 8576
rect 41328 8628 41380 8634
rect 41328 8570 41380 8576
rect 41696 8628 41748 8634
rect 41696 8570 41748 8576
rect 42064 8628 42116 8634
rect 42064 8570 42116 8576
rect 41602 8528 41658 8537
rect 41420 8492 41472 8498
rect 41602 8463 41658 8472
rect 41788 8492 41840 8498
rect 41420 8434 41472 8440
rect 41432 4434 41460 8434
rect 41616 8090 41644 8463
rect 41788 8434 41840 8440
rect 41880 8492 41932 8498
rect 41880 8434 41932 8440
rect 41604 8084 41656 8090
rect 41604 8026 41656 8032
rect 41604 7200 41656 7206
rect 41604 7142 41656 7148
rect 41340 4406 41460 4434
rect 41340 3482 41368 4406
rect 41616 3641 41644 7142
rect 41800 3670 41828 8434
rect 41788 3664 41840 3670
rect 41602 3632 41658 3641
rect 41788 3606 41840 3612
rect 41602 3567 41658 3576
rect 40776 3460 40828 3466
rect 41340 3454 41460 3482
rect 40776 3402 40828 3408
rect 40684 3188 40736 3194
rect 40684 3130 40736 3136
rect 41432 2961 41460 3454
rect 41418 2952 41474 2961
rect 41892 2922 41920 8434
rect 42248 8424 42300 8430
rect 42248 8366 42300 8372
rect 42260 2990 42288 8366
rect 42444 8362 42472 11194
rect 42812 8634 42840 11194
rect 42892 8968 42944 8974
rect 42892 8910 42944 8916
rect 42800 8628 42852 8634
rect 42800 8570 42852 8576
rect 42432 8356 42484 8362
rect 42432 8298 42484 8304
rect 42800 7336 42852 7342
rect 42800 7278 42852 7284
rect 42708 4276 42760 4282
rect 42708 4218 42760 4224
rect 42720 3602 42748 4218
rect 42708 3596 42760 3602
rect 42708 3538 42760 3544
rect 42248 2984 42300 2990
rect 42248 2926 42300 2932
rect 41418 2887 41474 2896
rect 41880 2916 41932 2922
rect 41880 2858 41932 2864
rect 42156 2644 42208 2650
rect 42156 2586 42208 2592
rect 42168 2553 42196 2586
rect 42154 2544 42210 2553
rect 42154 2479 42210 2488
rect 42812 56 42840 7278
rect 42904 7274 42932 8910
rect 42984 8492 43036 8498
rect 42984 8434 43036 8440
rect 42892 7268 42944 7274
rect 42892 7210 42944 7216
rect 42996 2854 43024 8434
rect 43180 8362 43208 11194
rect 43260 8900 43312 8906
rect 43260 8842 43312 8848
rect 43168 8356 43220 8362
rect 43168 8298 43220 8304
rect 43272 3194 43300 8842
rect 43548 8514 43576 11194
rect 43720 8832 43772 8838
rect 43720 8774 43772 8780
rect 43352 8492 43404 8498
rect 43548 8486 43668 8514
rect 43732 8498 43760 8774
rect 43916 8634 43944 11194
rect 43904 8628 43956 8634
rect 43904 8570 43956 8576
rect 43352 8434 43404 8440
rect 43364 3738 43392 8434
rect 43640 8430 43668 8486
rect 43720 8492 43772 8498
rect 43720 8434 43772 8440
rect 43996 8492 44048 8498
rect 43996 8434 44048 8440
rect 43628 8424 43680 8430
rect 44008 8378 44036 8434
rect 43628 8366 43680 8372
rect 43824 8350 44036 8378
rect 44284 8362 44312 11194
rect 44652 8634 44680 11194
rect 44822 9616 44878 9625
rect 44822 9551 44878 9560
rect 44640 8628 44692 8634
rect 44640 8570 44692 8576
rect 44364 8492 44416 8498
rect 44364 8434 44416 8440
rect 44272 8356 44324 8362
rect 43720 7744 43772 7750
rect 43720 7686 43772 7692
rect 43628 7472 43680 7478
rect 43628 7414 43680 7420
rect 43640 5778 43668 7414
rect 43732 6866 43760 7686
rect 43720 6860 43772 6866
rect 43720 6802 43772 6808
rect 43628 5772 43680 5778
rect 43628 5714 43680 5720
rect 43352 3732 43404 3738
rect 43352 3674 43404 3680
rect 43824 3482 43852 8350
rect 44272 8298 44324 8304
rect 43950 8188 44258 8197
rect 43950 8186 43956 8188
rect 44012 8186 44036 8188
rect 44092 8186 44116 8188
rect 44172 8186 44196 8188
rect 44252 8186 44258 8188
rect 44012 8134 44014 8186
rect 44194 8134 44196 8186
rect 43950 8132 43956 8134
rect 44012 8132 44036 8134
rect 44092 8132 44116 8134
rect 44172 8132 44196 8134
rect 44252 8132 44258 8134
rect 43950 8123 44258 8132
rect 44376 7970 44404 8434
rect 44836 8090 44864 9551
rect 45020 8922 45048 11194
rect 44928 8894 45048 8922
rect 44928 8566 44956 8894
rect 45388 8838 45416 11194
rect 45756 11098 45784 11194
rect 45848 11098 45876 11206
rect 45756 11070 45876 11098
rect 45926 9344 45982 9353
rect 45926 9279 45982 9288
rect 45560 9172 45612 9178
rect 45560 9114 45612 9120
rect 45468 8900 45520 8906
rect 45468 8842 45520 8848
rect 45376 8832 45428 8838
rect 45376 8774 45428 8780
rect 45010 8732 45318 8741
rect 45010 8730 45016 8732
rect 45072 8730 45096 8732
rect 45152 8730 45176 8732
rect 45232 8730 45256 8732
rect 45312 8730 45318 8732
rect 45072 8678 45074 8730
rect 45254 8678 45256 8730
rect 45010 8676 45016 8678
rect 45072 8676 45096 8678
rect 45152 8676 45176 8678
rect 45232 8676 45256 8678
rect 45312 8676 45318 8678
rect 45010 8667 45318 8676
rect 44916 8560 44968 8566
rect 44916 8502 44968 8508
rect 45480 8498 45508 8842
rect 45468 8492 45520 8498
rect 45468 8434 45520 8440
rect 45468 8356 45520 8362
rect 45468 8298 45520 8304
rect 44824 8084 44876 8090
rect 44824 8026 44876 8032
rect 44100 7942 44404 7970
rect 45098 7984 45154 7993
rect 44548 7948 44600 7954
rect 44100 7546 44128 7942
rect 45098 7919 45154 7928
rect 44548 7890 44600 7896
rect 44560 7546 44588 7890
rect 45112 7886 45140 7919
rect 45100 7880 45152 7886
rect 45100 7822 45152 7828
rect 45010 7644 45318 7653
rect 45010 7642 45016 7644
rect 45072 7642 45096 7644
rect 45152 7642 45176 7644
rect 45232 7642 45256 7644
rect 45312 7642 45318 7644
rect 45072 7590 45074 7642
rect 45254 7590 45256 7642
rect 45010 7588 45016 7590
rect 45072 7588 45096 7590
rect 45152 7588 45176 7590
rect 45232 7588 45256 7590
rect 45312 7588 45318 7590
rect 45010 7579 45318 7588
rect 44088 7540 44140 7546
rect 44088 7482 44140 7488
rect 44548 7540 44600 7546
rect 44548 7482 44600 7488
rect 45376 7404 45428 7410
rect 45376 7346 45428 7352
rect 43950 7100 44258 7109
rect 43950 7098 43956 7100
rect 44012 7098 44036 7100
rect 44092 7098 44116 7100
rect 44172 7098 44196 7100
rect 44252 7098 44258 7100
rect 44012 7046 44014 7098
rect 44194 7046 44196 7098
rect 43950 7044 43956 7046
rect 44012 7044 44036 7046
rect 44092 7044 44116 7046
rect 44172 7044 44196 7046
rect 44252 7044 44258 7046
rect 43950 7035 44258 7044
rect 45010 6556 45318 6565
rect 45010 6554 45016 6556
rect 45072 6554 45096 6556
rect 45152 6554 45176 6556
rect 45232 6554 45256 6556
rect 45312 6554 45318 6556
rect 45072 6502 45074 6554
rect 45254 6502 45256 6554
rect 45010 6500 45016 6502
rect 45072 6500 45096 6502
rect 45152 6500 45176 6502
rect 45232 6500 45256 6502
rect 45312 6500 45318 6502
rect 45010 6491 45318 6500
rect 43950 6012 44258 6021
rect 43950 6010 43956 6012
rect 44012 6010 44036 6012
rect 44092 6010 44116 6012
rect 44172 6010 44196 6012
rect 44252 6010 44258 6012
rect 44012 5958 44014 6010
rect 44194 5958 44196 6010
rect 43950 5956 43956 5958
rect 44012 5956 44036 5958
rect 44092 5956 44116 5958
rect 44172 5956 44196 5958
rect 44252 5956 44258 5958
rect 43950 5947 44258 5956
rect 44456 5636 44508 5642
rect 44456 5578 44508 5584
rect 44364 5092 44416 5098
rect 44364 5034 44416 5040
rect 43950 4924 44258 4933
rect 43950 4922 43956 4924
rect 44012 4922 44036 4924
rect 44092 4922 44116 4924
rect 44172 4922 44196 4924
rect 44252 4922 44258 4924
rect 44012 4870 44014 4922
rect 44194 4870 44196 4922
rect 43950 4868 43956 4870
rect 44012 4868 44036 4870
rect 44092 4868 44116 4870
rect 44172 4868 44196 4870
rect 44252 4868 44258 4870
rect 43950 4859 44258 4868
rect 44376 4078 44404 5034
rect 44364 4072 44416 4078
rect 44364 4014 44416 4020
rect 43950 3836 44258 3845
rect 43950 3834 43956 3836
rect 44012 3834 44036 3836
rect 44092 3834 44116 3836
rect 44172 3834 44196 3836
rect 44252 3834 44258 3836
rect 44012 3782 44014 3834
rect 44194 3782 44196 3834
rect 43950 3780 43956 3782
rect 44012 3780 44036 3782
rect 44092 3780 44116 3782
rect 44172 3780 44196 3782
rect 44252 3780 44258 3782
rect 43950 3771 44258 3780
rect 44180 3528 44232 3534
rect 44178 3496 44180 3505
rect 44232 3496 44234 3505
rect 43824 3454 43944 3482
rect 43812 3392 43864 3398
rect 43812 3334 43864 3340
rect 43260 3188 43312 3194
rect 43260 3130 43312 3136
rect 43824 3058 43852 3334
rect 43916 3194 43944 3454
rect 44178 3431 44234 3440
rect 43904 3188 43956 3194
rect 43904 3130 43956 3136
rect 44468 3126 44496 5578
rect 45010 5468 45318 5477
rect 45010 5466 45016 5468
rect 45072 5466 45096 5468
rect 45152 5466 45176 5468
rect 45232 5466 45256 5468
rect 45312 5466 45318 5468
rect 45072 5414 45074 5466
rect 45254 5414 45256 5466
rect 45010 5412 45016 5414
rect 45072 5412 45096 5414
rect 45152 5412 45176 5414
rect 45232 5412 45256 5414
rect 45312 5412 45318 5414
rect 45010 5403 45318 5412
rect 45010 4380 45318 4389
rect 45010 4378 45016 4380
rect 45072 4378 45096 4380
rect 45152 4378 45176 4380
rect 45232 4378 45256 4380
rect 45312 4378 45318 4380
rect 45072 4326 45074 4378
rect 45254 4326 45256 4378
rect 45010 4324 45016 4326
rect 45072 4324 45096 4326
rect 45152 4324 45176 4326
rect 45232 4324 45256 4326
rect 45312 4324 45318 4326
rect 45010 4315 45318 4324
rect 45010 3292 45318 3301
rect 45010 3290 45016 3292
rect 45072 3290 45096 3292
rect 45152 3290 45176 3292
rect 45232 3290 45256 3292
rect 45312 3290 45318 3292
rect 45072 3238 45074 3290
rect 45254 3238 45256 3290
rect 45010 3236 45016 3238
rect 45072 3236 45096 3238
rect 45152 3236 45176 3238
rect 45232 3236 45256 3238
rect 45312 3236 45318 3238
rect 45010 3227 45318 3236
rect 44456 3120 44508 3126
rect 44456 3062 44508 3068
rect 43076 3052 43128 3058
rect 43076 2994 43128 3000
rect 43812 3052 43864 3058
rect 43812 2994 43864 3000
rect 42984 2848 43036 2854
rect 42984 2790 43036 2796
rect 43088 2106 43116 2994
rect 43950 2748 44258 2757
rect 43950 2746 43956 2748
rect 44012 2746 44036 2748
rect 44092 2746 44116 2748
rect 44172 2746 44196 2748
rect 44252 2746 44258 2748
rect 44012 2694 44014 2746
rect 44194 2694 44196 2746
rect 43950 2692 43956 2694
rect 44012 2692 44036 2694
rect 44092 2692 44116 2694
rect 44172 2692 44196 2694
rect 44252 2692 44258 2694
rect 43950 2683 44258 2692
rect 45010 2204 45318 2213
rect 45010 2202 45016 2204
rect 45072 2202 45096 2204
rect 45152 2202 45176 2204
rect 45232 2202 45256 2204
rect 45312 2202 45318 2204
rect 45072 2150 45074 2202
rect 45254 2150 45256 2202
rect 45010 2148 45016 2150
rect 45072 2148 45096 2150
rect 45152 2148 45176 2150
rect 45232 2148 45256 2150
rect 45312 2148 45318 2150
rect 45010 2139 45318 2148
rect 43076 2100 43128 2106
rect 43076 2042 43128 2048
rect 45112 56 45232 82
rect 38568 2 38620 8
rect 40498 0 40554 56
rect 42798 0 42854 56
rect 45098 54 45232 56
rect 45098 0 45154 54
rect 45204 42 45232 54
rect 45388 42 45416 7346
rect 45480 7274 45508 8298
rect 45468 7268 45520 7274
rect 45468 7210 45520 7216
rect 45572 6798 45600 9114
rect 45650 9072 45706 9081
rect 45650 9007 45706 9016
rect 45664 8090 45692 9007
rect 45742 8392 45798 8401
rect 45742 8327 45798 8336
rect 45652 8084 45704 8090
rect 45652 8026 45704 8032
rect 45650 7848 45706 7857
rect 45650 7783 45706 7792
rect 45664 7410 45692 7783
rect 45756 7410 45784 8327
rect 45836 7880 45888 7886
rect 45836 7822 45888 7828
rect 45652 7404 45704 7410
rect 45652 7346 45704 7352
rect 45744 7404 45796 7410
rect 45744 7346 45796 7352
rect 45848 7002 45876 7822
rect 45940 7206 45968 9279
rect 46032 8634 46060 11206
rect 46110 11194 46166 11250
rect 46478 11194 46534 11250
rect 46846 11194 46902 11250
rect 47214 11194 47270 11250
rect 46020 8628 46072 8634
rect 46020 8570 46072 8576
rect 46124 8514 46152 11194
rect 46388 8832 46440 8838
rect 46294 8800 46350 8809
rect 46388 8774 46440 8780
rect 46294 8735 46350 8744
rect 46020 8492 46072 8498
rect 46124 8486 46244 8514
rect 46020 8434 46072 8440
rect 46032 8294 46060 8434
rect 46216 8430 46244 8486
rect 46204 8424 46256 8430
rect 46204 8366 46256 8372
rect 46020 8288 46072 8294
rect 46020 8230 46072 8236
rect 46020 8016 46072 8022
rect 46018 7984 46020 7993
rect 46072 7984 46074 7993
rect 46018 7919 46074 7928
rect 46204 7880 46256 7886
rect 46204 7822 46256 7828
rect 46216 7546 46244 7822
rect 46204 7540 46256 7546
rect 46204 7482 46256 7488
rect 46308 7206 46336 8735
rect 46400 8362 46428 8774
rect 46388 8356 46440 8362
rect 46388 8298 46440 8304
rect 46492 8090 46520 11194
rect 46572 8968 46624 8974
rect 46572 8910 46624 8916
rect 46584 8498 46612 8910
rect 46572 8492 46624 8498
rect 46572 8434 46624 8440
rect 46570 8256 46626 8265
rect 46570 8191 46626 8200
rect 46480 8084 46532 8090
rect 46480 8026 46532 8032
rect 46584 7546 46612 8191
rect 46860 8090 46888 11194
rect 47030 8528 47086 8537
rect 47030 8463 47086 8472
rect 46848 8084 46900 8090
rect 46848 8026 46900 8032
rect 46664 7880 46716 7886
rect 46664 7822 46716 7828
rect 46572 7540 46624 7546
rect 46572 7482 46624 7488
rect 46676 7274 46704 7822
rect 46940 7540 46992 7546
rect 46940 7482 46992 7488
rect 46952 7449 46980 7482
rect 46938 7440 46994 7449
rect 46756 7404 46808 7410
rect 46938 7375 46994 7384
rect 46756 7346 46808 7352
rect 46664 7268 46716 7274
rect 46664 7210 46716 7216
rect 45928 7200 45980 7206
rect 45928 7142 45980 7148
rect 46296 7200 46348 7206
rect 46296 7142 46348 7148
rect 45836 6996 45888 7002
rect 45836 6938 45888 6944
rect 46662 6896 46718 6905
rect 46662 6831 46718 6840
rect 45560 6792 45612 6798
rect 45560 6734 45612 6740
rect 46112 6792 46164 6798
rect 46112 6734 46164 6740
rect 46204 6792 46256 6798
rect 46204 6734 46256 6740
rect 46020 6656 46072 6662
rect 46020 6598 46072 6604
rect 46032 6390 46060 6598
rect 46020 6384 46072 6390
rect 46020 6326 46072 6332
rect 46124 5681 46152 6734
rect 46216 6186 46244 6734
rect 46676 6662 46704 6831
rect 46296 6656 46348 6662
rect 46296 6598 46348 6604
rect 46664 6656 46716 6662
rect 46664 6598 46716 6604
rect 46308 6361 46336 6598
rect 46294 6352 46350 6361
rect 46294 6287 46350 6296
rect 46388 6316 46440 6322
rect 46388 6258 46440 6264
rect 46204 6180 46256 6186
rect 46204 6122 46256 6128
rect 46400 5914 46428 6258
rect 46572 6112 46624 6118
rect 46572 6054 46624 6060
rect 46388 5908 46440 5914
rect 46388 5850 46440 5856
rect 46584 5817 46612 6054
rect 46570 5808 46626 5817
rect 46570 5743 46626 5752
rect 46110 5672 46166 5681
rect 46110 5607 46166 5616
rect 46768 3942 46796 7346
rect 47044 6662 47072 8463
rect 47228 8022 47256 11194
rect 47490 9888 47546 9897
rect 47490 9823 47546 9832
rect 47216 8016 47268 8022
rect 47216 7958 47268 7964
rect 47306 7712 47362 7721
rect 47306 7647 47362 7656
rect 47320 7546 47348 7647
rect 47308 7540 47360 7546
rect 47308 7482 47360 7488
rect 47124 7404 47176 7410
rect 47124 7346 47176 7352
rect 47032 6656 47084 6662
rect 46938 6624 46994 6633
rect 47032 6598 47084 6604
rect 46938 6559 46994 6568
rect 46952 6458 46980 6559
rect 46940 6452 46992 6458
rect 46940 6394 46992 6400
rect 47032 5568 47084 5574
rect 47030 5536 47032 5545
rect 47084 5536 47086 5545
rect 47030 5471 47086 5480
rect 46940 5024 46992 5030
rect 46938 4992 46940 5001
rect 46992 4992 46994 5001
rect 46938 4927 46994 4936
rect 47136 4826 47164 7346
rect 47216 7336 47268 7342
rect 47216 7278 47268 7284
rect 47124 4820 47176 4826
rect 47124 4762 47176 4768
rect 47124 4548 47176 4554
rect 47124 4490 47176 4496
rect 47032 4480 47084 4486
rect 47030 4448 47032 4457
rect 47084 4448 47086 4457
rect 47030 4383 47086 4392
rect 46756 3936 46808 3942
rect 46940 3936 46992 3942
rect 46756 3878 46808 3884
rect 46938 3904 46940 3913
rect 46992 3904 46994 3913
rect 46938 3839 46994 3848
rect 47032 3392 47084 3398
rect 47030 3360 47032 3369
rect 47084 3360 47086 3369
rect 47030 3295 47086 3304
rect 46754 3088 46810 3097
rect 47136 3058 47164 4490
rect 46754 3023 46756 3032
rect 46808 3023 46810 3032
rect 47124 3052 47176 3058
rect 46756 2994 46808 3000
rect 47124 2994 47176 3000
rect 46940 2848 46992 2854
rect 46938 2816 46940 2825
rect 46992 2816 46994 2825
rect 46938 2751 46994 2760
rect 45836 2644 45888 2650
rect 45836 2586 45888 2592
rect 45650 2544 45706 2553
rect 45650 2479 45706 2488
rect 45664 2446 45692 2479
rect 45652 2440 45704 2446
rect 45652 2382 45704 2388
rect 45848 2009 45876 2586
rect 46204 2304 46256 2310
rect 46204 2246 46256 2252
rect 46572 2304 46624 2310
rect 46940 2304 46992 2310
rect 46572 2246 46624 2252
rect 46938 2272 46940 2281
rect 46992 2272 46994 2281
rect 45834 2000 45890 2009
rect 45834 1935 45890 1944
rect 46216 1737 46244 2246
rect 46202 1728 46258 1737
rect 46202 1663 46258 1672
rect 46584 1465 46612 2246
rect 46938 2207 46994 2216
rect 46570 1456 46626 1465
rect 46570 1391 46626 1400
rect 45204 14 45416 42
rect 47228 42 47256 7278
rect 47398 7168 47454 7177
rect 47398 7103 47454 7112
rect 47412 6662 47440 7103
rect 47400 6656 47452 6662
rect 47400 6598 47452 6604
rect 47504 6458 47532 9823
rect 47492 6452 47544 6458
rect 47492 6394 47544 6400
rect 47398 6080 47454 6089
rect 47398 6015 47454 6024
rect 47412 5914 47440 6015
rect 47400 5908 47452 5914
rect 47400 5850 47452 5856
rect 47308 5364 47360 5370
rect 47308 5306 47360 5312
rect 47320 5273 47348 5306
rect 47306 5264 47362 5273
rect 47306 5199 47362 5208
rect 47400 4752 47452 4758
rect 47398 4720 47400 4729
rect 47452 4720 47454 4729
rect 47398 4655 47454 4664
rect 47306 4176 47362 4185
rect 47306 4111 47362 4120
rect 47320 4010 47348 4111
rect 47308 4004 47360 4010
rect 47308 3946 47360 3952
rect 47400 3664 47452 3670
rect 47398 3632 47400 3641
rect 47452 3632 47454 3641
rect 47398 3567 47454 3576
rect 47308 3188 47360 3194
rect 47308 3130 47360 3136
rect 47320 3097 47348 3130
rect 47306 3088 47362 3097
rect 47306 3023 47362 3032
rect 47308 2576 47360 2582
rect 47306 2544 47308 2553
rect 47360 2544 47362 2553
rect 47306 2479 47362 2488
rect 47320 56 47440 82
rect 47320 54 47454 56
rect 47320 42 47348 54
rect 47228 14 47348 42
rect 47398 0 47454 54
<< via2 >>
rect 1122 9424 1178 9480
rect 202 9288 258 9344
rect 1306 8200 1362 8256
rect 3016 8730 3072 8732
rect 3096 8730 3152 8732
rect 3176 8730 3232 8732
rect 3256 8730 3312 8732
rect 3016 8678 3062 8730
rect 3062 8678 3072 8730
rect 3096 8678 3126 8730
rect 3126 8678 3138 8730
rect 3138 8678 3152 8730
rect 3176 8678 3190 8730
rect 3190 8678 3202 8730
rect 3202 8678 3232 8730
rect 3256 8678 3266 8730
rect 3266 8678 3312 8730
rect 3016 8676 3072 8678
rect 3096 8676 3152 8678
rect 3176 8676 3232 8678
rect 3256 8676 3312 8678
rect 1956 8186 2012 8188
rect 2036 8186 2092 8188
rect 2116 8186 2172 8188
rect 2196 8186 2252 8188
rect 1956 8134 2002 8186
rect 2002 8134 2012 8186
rect 2036 8134 2066 8186
rect 2066 8134 2078 8186
rect 2078 8134 2092 8186
rect 2116 8134 2130 8186
rect 2130 8134 2142 8186
rect 2142 8134 2172 8186
rect 2196 8134 2206 8186
rect 2206 8134 2252 8186
rect 1956 8132 2012 8134
rect 2036 8132 2092 8134
rect 2116 8132 2172 8134
rect 2196 8132 2252 8134
rect 1122 7384 1178 7440
rect 1956 7098 2012 7100
rect 2036 7098 2092 7100
rect 2116 7098 2172 7100
rect 2196 7098 2252 7100
rect 1956 7046 2002 7098
rect 2002 7046 2012 7098
rect 2036 7046 2066 7098
rect 2066 7046 2078 7098
rect 2078 7046 2092 7098
rect 2116 7046 2130 7098
rect 2130 7046 2142 7098
rect 2142 7046 2172 7098
rect 2196 7046 2206 7098
rect 2206 7046 2252 7098
rect 1956 7044 2012 7046
rect 2036 7044 2092 7046
rect 2116 7044 2172 7046
rect 2196 7044 2252 7046
rect 1956 6010 2012 6012
rect 2036 6010 2092 6012
rect 2116 6010 2172 6012
rect 2196 6010 2252 6012
rect 1956 5958 2002 6010
rect 2002 5958 2012 6010
rect 2036 5958 2066 6010
rect 2066 5958 2078 6010
rect 2078 5958 2092 6010
rect 2116 5958 2130 6010
rect 2130 5958 2142 6010
rect 2142 5958 2172 6010
rect 2196 5958 2206 6010
rect 2206 5958 2252 6010
rect 1956 5956 2012 5958
rect 2036 5956 2092 5958
rect 2116 5956 2172 5958
rect 2196 5956 2252 5958
rect 1956 4922 2012 4924
rect 2036 4922 2092 4924
rect 2116 4922 2172 4924
rect 2196 4922 2252 4924
rect 1956 4870 2002 4922
rect 2002 4870 2012 4922
rect 2036 4870 2066 4922
rect 2066 4870 2078 4922
rect 2078 4870 2092 4922
rect 2116 4870 2130 4922
rect 2130 4870 2142 4922
rect 2142 4870 2172 4922
rect 2196 4870 2206 4922
rect 2206 4870 2252 4922
rect 1956 4868 2012 4870
rect 2036 4868 2092 4870
rect 2116 4868 2172 4870
rect 2196 4868 2252 4870
rect 1956 3834 2012 3836
rect 2036 3834 2092 3836
rect 2116 3834 2172 3836
rect 2196 3834 2252 3836
rect 1956 3782 2002 3834
rect 2002 3782 2012 3834
rect 2036 3782 2066 3834
rect 2066 3782 2078 3834
rect 2078 3782 2092 3834
rect 2116 3782 2130 3834
rect 2130 3782 2142 3834
rect 2142 3782 2172 3834
rect 2196 3782 2206 3834
rect 2206 3782 2252 3834
rect 1956 3780 2012 3782
rect 2036 3780 2092 3782
rect 2116 3780 2172 3782
rect 2196 3780 2252 3782
rect 2410 7828 2412 7848
rect 2412 7828 2464 7848
rect 2464 7828 2466 7848
rect 2410 7792 2466 7828
rect 4618 8744 4674 8800
rect 5170 9560 5226 9616
rect 4618 7928 4674 7984
rect 5354 7964 5356 7984
rect 5356 7964 5408 7984
rect 5408 7964 5410 7984
rect 5354 7928 5410 7964
rect 3016 7642 3072 7644
rect 3096 7642 3152 7644
rect 3176 7642 3232 7644
rect 3256 7642 3312 7644
rect 3016 7590 3062 7642
rect 3062 7590 3072 7642
rect 3096 7590 3126 7642
rect 3126 7590 3138 7642
rect 3138 7590 3152 7642
rect 3176 7590 3190 7642
rect 3190 7590 3202 7642
rect 3202 7590 3232 7642
rect 3256 7590 3266 7642
rect 3266 7590 3312 7642
rect 3016 7588 3072 7590
rect 3096 7588 3152 7590
rect 3176 7588 3232 7590
rect 3256 7588 3312 7590
rect 5998 7248 6054 7304
rect 2778 6568 2834 6624
rect 2686 5208 2742 5264
rect 2686 4936 2742 4992
rect 3016 6554 3072 6556
rect 3096 6554 3152 6556
rect 3176 6554 3232 6556
rect 3256 6554 3312 6556
rect 3016 6502 3062 6554
rect 3062 6502 3072 6554
rect 3096 6502 3126 6554
rect 3126 6502 3138 6554
rect 3138 6502 3152 6554
rect 3176 6502 3190 6554
rect 3190 6502 3202 6554
rect 3202 6502 3232 6554
rect 3256 6502 3266 6554
rect 3266 6502 3312 6554
rect 3016 6500 3072 6502
rect 3096 6500 3152 6502
rect 3176 6500 3232 6502
rect 3256 6500 3312 6502
rect 5630 6160 5686 6216
rect 3016 5466 3072 5468
rect 3096 5466 3152 5468
rect 3176 5466 3232 5468
rect 3256 5466 3312 5468
rect 3016 5414 3062 5466
rect 3062 5414 3072 5466
rect 3096 5414 3126 5466
rect 3126 5414 3138 5466
rect 3138 5414 3152 5466
rect 3176 5414 3190 5466
rect 3190 5414 3202 5466
rect 3202 5414 3232 5466
rect 3256 5414 3266 5466
rect 3266 5414 3312 5466
rect 3016 5412 3072 5414
rect 3096 5412 3152 5414
rect 3176 5412 3232 5414
rect 3256 5412 3312 5414
rect 3146 5208 3202 5264
rect 2870 5072 2926 5128
rect 3016 4378 3072 4380
rect 3096 4378 3152 4380
rect 3176 4378 3232 4380
rect 3256 4378 3312 4380
rect 3016 4326 3062 4378
rect 3062 4326 3072 4378
rect 3096 4326 3126 4378
rect 3126 4326 3138 4378
rect 3138 4326 3152 4378
rect 3176 4326 3190 4378
rect 3190 4326 3202 4378
rect 3202 4326 3232 4378
rect 3256 4326 3266 4378
rect 3266 4326 3312 4378
rect 3016 4324 3072 4326
rect 3096 4324 3152 4326
rect 3176 4324 3232 4326
rect 3256 4324 3312 4326
rect 3016 3290 3072 3292
rect 3096 3290 3152 3292
rect 3176 3290 3232 3292
rect 3256 3290 3312 3292
rect 3016 3238 3062 3290
rect 3062 3238 3072 3290
rect 3096 3238 3126 3290
rect 3126 3238 3138 3290
rect 3138 3238 3152 3290
rect 3176 3238 3190 3290
rect 3190 3238 3202 3290
rect 3202 3238 3232 3290
rect 3256 3238 3266 3290
rect 3266 3238 3312 3290
rect 3016 3236 3072 3238
rect 3096 3236 3152 3238
rect 3176 3236 3232 3238
rect 3256 3236 3312 3238
rect 1956 2746 2012 2748
rect 2036 2746 2092 2748
rect 2116 2746 2172 2748
rect 2196 2746 2252 2748
rect 1956 2694 2002 2746
rect 2002 2694 2012 2746
rect 2036 2694 2066 2746
rect 2066 2694 2078 2746
rect 2078 2694 2092 2746
rect 2116 2694 2130 2746
rect 2130 2694 2142 2746
rect 2142 2694 2172 2746
rect 2196 2694 2206 2746
rect 2206 2694 2252 2746
rect 1956 2692 2012 2694
rect 2036 2692 2092 2694
rect 2116 2692 2172 2694
rect 2196 2692 2252 2694
rect 7746 8880 7802 8936
rect 8298 8336 8354 8392
rect 7956 8186 8012 8188
rect 8036 8186 8092 8188
rect 8116 8186 8172 8188
rect 8196 8186 8252 8188
rect 7956 8134 8002 8186
rect 8002 8134 8012 8186
rect 8036 8134 8066 8186
rect 8066 8134 8078 8186
rect 8078 8134 8092 8186
rect 8116 8134 8130 8186
rect 8130 8134 8142 8186
rect 8142 8134 8172 8186
rect 8196 8134 8206 8186
rect 8206 8134 8252 8186
rect 7956 8132 8012 8134
rect 8036 8132 8092 8134
rect 8116 8132 8172 8134
rect 8196 8132 8252 8134
rect 7956 7098 8012 7100
rect 8036 7098 8092 7100
rect 8116 7098 8172 7100
rect 8196 7098 8252 7100
rect 7956 7046 8002 7098
rect 8002 7046 8012 7098
rect 8036 7046 8066 7098
rect 8066 7046 8078 7098
rect 8078 7046 8092 7098
rect 8116 7046 8130 7098
rect 8130 7046 8142 7098
rect 8142 7046 8172 7098
rect 8196 7046 8206 7098
rect 8206 7046 8252 7098
rect 7956 7044 8012 7046
rect 8036 7044 8092 7046
rect 8116 7044 8172 7046
rect 8196 7044 8252 7046
rect 7956 6010 8012 6012
rect 8036 6010 8092 6012
rect 8116 6010 8172 6012
rect 8196 6010 8252 6012
rect 7956 5958 8002 6010
rect 8002 5958 8012 6010
rect 8036 5958 8066 6010
rect 8066 5958 8078 6010
rect 8078 5958 8092 6010
rect 8116 5958 8130 6010
rect 8130 5958 8142 6010
rect 8142 5958 8172 6010
rect 8196 5958 8206 6010
rect 8206 5958 8252 6010
rect 7956 5956 8012 5958
rect 8036 5956 8092 5958
rect 8116 5956 8172 5958
rect 8196 5956 8252 5958
rect 7470 5208 7526 5264
rect 7956 4922 8012 4924
rect 8036 4922 8092 4924
rect 8116 4922 8172 4924
rect 8196 4922 8252 4924
rect 7956 4870 8002 4922
rect 8002 4870 8012 4922
rect 8036 4870 8066 4922
rect 8066 4870 8078 4922
rect 8078 4870 8092 4922
rect 8116 4870 8130 4922
rect 8130 4870 8142 4922
rect 8142 4870 8172 4922
rect 8196 4870 8206 4922
rect 8206 4870 8252 4922
rect 7956 4868 8012 4870
rect 8036 4868 8092 4870
rect 8116 4868 8172 4870
rect 8196 4868 8252 4870
rect 7470 4664 7526 4720
rect 9016 8730 9072 8732
rect 9096 8730 9152 8732
rect 9176 8730 9232 8732
rect 9256 8730 9312 8732
rect 9016 8678 9062 8730
rect 9062 8678 9072 8730
rect 9096 8678 9126 8730
rect 9126 8678 9138 8730
rect 9138 8678 9152 8730
rect 9176 8678 9190 8730
rect 9190 8678 9202 8730
rect 9202 8678 9232 8730
rect 9256 8678 9266 8730
rect 9266 8678 9312 8730
rect 9016 8676 9072 8678
rect 9096 8676 9152 8678
rect 9176 8676 9232 8678
rect 9256 8676 9312 8678
rect 10874 10920 10930 10976
rect 9016 7642 9072 7644
rect 9096 7642 9152 7644
rect 9176 7642 9232 7644
rect 9256 7642 9312 7644
rect 9016 7590 9062 7642
rect 9062 7590 9072 7642
rect 9096 7590 9126 7642
rect 9126 7590 9138 7642
rect 9138 7590 9152 7642
rect 9176 7590 9190 7642
rect 9190 7590 9202 7642
rect 9202 7590 9232 7642
rect 9256 7590 9266 7642
rect 9266 7590 9312 7642
rect 9016 7588 9072 7590
rect 9096 7588 9152 7590
rect 9176 7588 9232 7590
rect 9256 7588 9312 7590
rect 9016 6554 9072 6556
rect 9096 6554 9152 6556
rect 9176 6554 9232 6556
rect 9256 6554 9312 6556
rect 9016 6502 9062 6554
rect 9062 6502 9072 6554
rect 9096 6502 9126 6554
rect 9126 6502 9138 6554
rect 9138 6502 9152 6554
rect 9176 6502 9190 6554
rect 9190 6502 9202 6554
rect 9202 6502 9232 6554
rect 9256 6502 9266 6554
rect 9266 6502 9312 6554
rect 9016 6500 9072 6502
rect 9096 6500 9152 6502
rect 9176 6500 9232 6502
rect 9256 6500 9312 6502
rect 9494 6024 9550 6080
rect 9862 6704 9918 6760
rect 11150 7656 11206 7712
rect 11978 10784 12034 10840
rect 12438 8200 12494 8256
rect 11058 6296 11114 6352
rect 12806 8200 12862 8256
rect 9016 5466 9072 5468
rect 9096 5466 9152 5468
rect 9176 5466 9232 5468
rect 9256 5466 9312 5468
rect 9016 5414 9062 5466
rect 9062 5414 9072 5466
rect 9096 5414 9126 5466
rect 9126 5414 9138 5466
rect 9138 5414 9152 5466
rect 9176 5414 9190 5466
rect 9190 5414 9202 5466
rect 9202 5414 9232 5466
rect 9256 5414 9266 5466
rect 9266 5414 9312 5466
rect 9016 5412 9072 5414
rect 9096 5412 9152 5414
rect 9176 5412 9232 5414
rect 9256 5412 9312 5414
rect 9678 5344 9734 5400
rect 9586 5228 9642 5264
rect 9586 5208 9588 5228
rect 9588 5208 9640 5228
rect 9640 5208 9642 5228
rect 9016 4378 9072 4380
rect 9096 4378 9152 4380
rect 9176 4378 9232 4380
rect 9256 4378 9312 4380
rect 9016 4326 9062 4378
rect 9062 4326 9072 4378
rect 9096 4326 9126 4378
rect 9126 4326 9138 4378
rect 9138 4326 9152 4378
rect 9176 4326 9190 4378
rect 9190 4326 9202 4378
rect 9202 4326 9232 4378
rect 9256 4326 9266 4378
rect 9266 4326 9312 4378
rect 9016 4324 9072 4326
rect 9096 4324 9152 4326
rect 9176 4324 9232 4326
rect 9256 4324 9312 4326
rect 13956 8186 14012 8188
rect 14036 8186 14092 8188
rect 14116 8186 14172 8188
rect 14196 8186 14252 8188
rect 13956 8134 14002 8186
rect 14002 8134 14012 8186
rect 14036 8134 14066 8186
rect 14066 8134 14078 8186
rect 14078 8134 14092 8186
rect 14116 8134 14130 8186
rect 14130 8134 14142 8186
rect 14142 8134 14172 8186
rect 14196 8134 14206 8186
rect 14206 8134 14252 8186
rect 13956 8132 14012 8134
rect 14036 8132 14092 8134
rect 14116 8132 14172 8134
rect 14196 8132 14252 8134
rect 14278 7656 14334 7712
rect 13542 6840 13598 6896
rect 7956 3834 8012 3836
rect 8036 3834 8092 3836
rect 8116 3834 8172 3836
rect 8196 3834 8252 3836
rect 7956 3782 8002 3834
rect 8002 3782 8012 3834
rect 8036 3782 8066 3834
rect 8066 3782 8078 3834
rect 8078 3782 8092 3834
rect 8116 3782 8130 3834
rect 8130 3782 8142 3834
rect 8142 3782 8172 3834
rect 8196 3782 8206 3834
rect 8206 3782 8252 3834
rect 7956 3780 8012 3782
rect 8036 3780 8092 3782
rect 8116 3780 8172 3782
rect 8196 3780 8252 3782
rect 9016 3290 9072 3292
rect 9096 3290 9152 3292
rect 9176 3290 9232 3292
rect 9256 3290 9312 3292
rect 9016 3238 9062 3290
rect 9062 3238 9072 3290
rect 9096 3238 9126 3290
rect 9126 3238 9138 3290
rect 9138 3238 9152 3290
rect 9176 3238 9190 3290
rect 9190 3238 9202 3290
rect 9202 3238 9232 3290
rect 9256 3238 9266 3290
rect 9266 3238 9312 3290
rect 9016 3236 9072 3238
rect 9096 3236 9152 3238
rect 9176 3236 9232 3238
rect 9256 3236 9312 3238
rect 9402 3168 9458 3224
rect 15016 8730 15072 8732
rect 15096 8730 15152 8732
rect 15176 8730 15232 8732
rect 15256 8730 15312 8732
rect 15016 8678 15062 8730
rect 15062 8678 15072 8730
rect 15096 8678 15126 8730
rect 15126 8678 15138 8730
rect 15138 8678 15152 8730
rect 15176 8678 15190 8730
rect 15190 8678 15202 8730
rect 15202 8678 15232 8730
rect 15256 8678 15266 8730
rect 15266 8678 15312 8730
rect 15016 8676 15072 8678
rect 15096 8676 15152 8678
rect 15176 8676 15232 8678
rect 15256 8676 15312 8678
rect 15016 7642 15072 7644
rect 15096 7642 15152 7644
rect 15176 7642 15232 7644
rect 15256 7642 15312 7644
rect 15016 7590 15062 7642
rect 15062 7590 15072 7642
rect 15096 7590 15126 7642
rect 15126 7590 15138 7642
rect 15138 7590 15152 7642
rect 15176 7590 15190 7642
rect 15190 7590 15202 7642
rect 15202 7590 15232 7642
rect 15256 7590 15266 7642
rect 15266 7590 15312 7642
rect 15016 7588 15072 7590
rect 15096 7588 15152 7590
rect 15176 7588 15232 7590
rect 15256 7588 15312 7590
rect 15566 7692 15568 7712
rect 15568 7692 15620 7712
rect 15620 7692 15622 7712
rect 15566 7656 15622 7692
rect 13956 7098 14012 7100
rect 14036 7098 14092 7100
rect 14116 7098 14172 7100
rect 14196 7098 14252 7100
rect 13956 7046 14002 7098
rect 14002 7046 14012 7098
rect 14036 7046 14066 7098
rect 14066 7046 14078 7098
rect 14078 7046 14092 7098
rect 14116 7046 14130 7098
rect 14130 7046 14142 7098
rect 14142 7046 14172 7098
rect 14196 7046 14206 7098
rect 14206 7046 14252 7098
rect 13956 7044 14012 7046
rect 14036 7044 14092 7046
rect 14116 7044 14172 7046
rect 14196 7044 14252 7046
rect 15016 6554 15072 6556
rect 15096 6554 15152 6556
rect 15176 6554 15232 6556
rect 15256 6554 15312 6556
rect 15016 6502 15062 6554
rect 15062 6502 15072 6554
rect 15096 6502 15126 6554
rect 15126 6502 15138 6554
rect 15138 6502 15152 6554
rect 15176 6502 15190 6554
rect 15190 6502 15202 6554
rect 15202 6502 15232 6554
rect 15256 6502 15266 6554
rect 15266 6502 15312 6554
rect 15016 6500 15072 6502
rect 15096 6500 15152 6502
rect 15176 6500 15232 6502
rect 15256 6500 15312 6502
rect 13956 6010 14012 6012
rect 14036 6010 14092 6012
rect 14116 6010 14172 6012
rect 14196 6010 14252 6012
rect 13956 5958 14002 6010
rect 14002 5958 14012 6010
rect 14036 5958 14066 6010
rect 14066 5958 14078 6010
rect 14078 5958 14092 6010
rect 14116 5958 14130 6010
rect 14130 5958 14142 6010
rect 14142 5958 14172 6010
rect 14196 5958 14206 6010
rect 14206 5958 14252 6010
rect 13956 5956 14012 5958
rect 14036 5956 14092 5958
rect 14116 5956 14172 5958
rect 14196 5956 14252 5958
rect 14922 5652 14924 5672
rect 14924 5652 14976 5672
rect 14976 5652 14978 5672
rect 14922 5616 14978 5652
rect 15016 5466 15072 5468
rect 15096 5466 15152 5468
rect 15176 5466 15232 5468
rect 15256 5466 15312 5468
rect 15016 5414 15062 5466
rect 15062 5414 15072 5466
rect 15096 5414 15126 5466
rect 15126 5414 15138 5466
rect 15138 5414 15152 5466
rect 15176 5414 15190 5466
rect 15190 5414 15202 5466
rect 15202 5414 15232 5466
rect 15256 5414 15266 5466
rect 15266 5414 15312 5466
rect 15016 5412 15072 5414
rect 15096 5412 15152 5414
rect 15176 5412 15232 5414
rect 15256 5412 15312 5414
rect 14830 5344 14886 5400
rect 14830 5072 14886 5128
rect 13956 4922 14012 4924
rect 14036 4922 14092 4924
rect 14116 4922 14172 4924
rect 14196 4922 14252 4924
rect 13956 4870 14002 4922
rect 14002 4870 14012 4922
rect 14036 4870 14066 4922
rect 14066 4870 14078 4922
rect 14078 4870 14092 4922
rect 14116 4870 14130 4922
rect 14130 4870 14142 4922
rect 14142 4870 14172 4922
rect 14196 4870 14206 4922
rect 14206 4870 14252 4922
rect 13956 4868 14012 4870
rect 14036 4868 14092 4870
rect 14116 4868 14172 4870
rect 14196 4868 14252 4870
rect 13634 4528 13690 4584
rect 15016 4378 15072 4380
rect 15096 4378 15152 4380
rect 15176 4378 15232 4380
rect 15256 4378 15312 4380
rect 15016 4326 15062 4378
rect 15062 4326 15072 4378
rect 15096 4326 15126 4378
rect 15126 4326 15138 4378
rect 15138 4326 15152 4378
rect 15176 4326 15190 4378
rect 15190 4326 15202 4378
rect 15202 4326 15232 4378
rect 15256 4326 15266 4378
rect 15266 4326 15312 4378
rect 15016 4324 15072 4326
rect 15096 4324 15152 4326
rect 15176 4324 15232 4326
rect 15256 4324 15312 4326
rect 16026 10648 16082 10704
rect 16394 11056 16450 11112
rect 16578 7404 16634 7440
rect 16578 7384 16580 7404
rect 16580 7384 16632 7404
rect 16632 7384 16634 7404
rect 17406 4936 17462 4992
rect 18234 6296 18290 6352
rect 17866 4664 17922 4720
rect 14830 3848 14886 3904
rect 13956 3834 14012 3836
rect 14036 3834 14092 3836
rect 14116 3834 14172 3836
rect 14196 3834 14252 3836
rect 13956 3782 14002 3834
rect 14002 3782 14012 3834
rect 14036 3782 14066 3834
rect 14066 3782 14078 3834
rect 14078 3782 14092 3834
rect 14116 3782 14130 3834
rect 14130 3782 14142 3834
rect 14142 3782 14172 3834
rect 14196 3782 14206 3834
rect 14206 3782 14252 3834
rect 13956 3780 14012 3782
rect 14036 3780 14092 3782
rect 14116 3780 14172 3782
rect 14196 3780 14252 3782
rect 15016 3290 15072 3292
rect 15096 3290 15152 3292
rect 15176 3290 15232 3292
rect 15256 3290 15312 3292
rect 15016 3238 15062 3290
rect 15062 3238 15072 3290
rect 15096 3238 15126 3290
rect 15126 3238 15138 3290
rect 15138 3238 15152 3290
rect 15176 3238 15190 3290
rect 15190 3238 15202 3290
rect 15202 3238 15232 3290
rect 15256 3238 15266 3290
rect 15266 3238 15312 3290
rect 15016 3236 15072 3238
rect 15096 3236 15152 3238
rect 15176 3236 15232 3238
rect 15256 3236 15312 3238
rect 7956 2746 8012 2748
rect 8036 2746 8092 2748
rect 8116 2746 8172 2748
rect 8196 2746 8252 2748
rect 7956 2694 8002 2746
rect 8002 2694 8012 2746
rect 8036 2694 8066 2746
rect 8066 2694 8078 2746
rect 8078 2694 8092 2746
rect 8116 2694 8130 2746
rect 8130 2694 8142 2746
rect 8142 2694 8172 2746
rect 8196 2694 8206 2746
rect 8206 2694 8252 2746
rect 7956 2692 8012 2694
rect 8036 2692 8092 2694
rect 8116 2692 8172 2694
rect 8196 2692 8252 2694
rect 3016 2202 3072 2204
rect 3096 2202 3152 2204
rect 3176 2202 3232 2204
rect 3256 2202 3312 2204
rect 3016 2150 3062 2202
rect 3062 2150 3072 2202
rect 3096 2150 3126 2202
rect 3126 2150 3138 2202
rect 3138 2150 3152 2202
rect 3176 2150 3190 2202
rect 3190 2150 3202 2202
rect 3202 2150 3232 2202
rect 3256 2150 3266 2202
rect 3266 2150 3312 2202
rect 3016 2148 3072 2150
rect 3096 2148 3152 2150
rect 3176 2148 3232 2150
rect 3256 2148 3312 2150
rect 1306 1400 1362 1456
rect 14830 3168 14886 3224
rect 17958 4004 18014 4040
rect 17958 3984 17960 4004
rect 17960 3984 18012 4004
rect 18012 3984 18014 4004
rect 19522 9696 19578 9752
rect 19798 9152 19854 9208
rect 20718 9696 20774 9752
rect 20442 9288 20498 9344
rect 19956 8186 20012 8188
rect 20036 8186 20092 8188
rect 20116 8186 20172 8188
rect 20196 8186 20252 8188
rect 19956 8134 20002 8186
rect 20002 8134 20012 8186
rect 20036 8134 20066 8186
rect 20066 8134 20078 8186
rect 20078 8134 20092 8186
rect 20116 8134 20130 8186
rect 20130 8134 20142 8186
rect 20142 8134 20172 8186
rect 20196 8134 20206 8186
rect 20206 8134 20252 8186
rect 19956 8132 20012 8134
rect 20036 8132 20092 8134
rect 20116 8132 20172 8134
rect 20196 8132 20252 8134
rect 19956 7098 20012 7100
rect 20036 7098 20092 7100
rect 20116 7098 20172 7100
rect 20196 7098 20252 7100
rect 19956 7046 20002 7098
rect 20002 7046 20012 7098
rect 20036 7046 20066 7098
rect 20066 7046 20078 7098
rect 20078 7046 20092 7098
rect 20116 7046 20130 7098
rect 20130 7046 20142 7098
rect 20142 7046 20172 7098
rect 20196 7046 20206 7098
rect 20206 7046 20252 7098
rect 19956 7044 20012 7046
rect 20036 7044 20092 7046
rect 20116 7044 20172 7046
rect 20196 7044 20252 7046
rect 19956 6010 20012 6012
rect 20036 6010 20092 6012
rect 20116 6010 20172 6012
rect 20196 6010 20252 6012
rect 19956 5958 20002 6010
rect 20002 5958 20012 6010
rect 20036 5958 20066 6010
rect 20066 5958 20078 6010
rect 20078 5958 20092 6010
rect 20116 5958 20130 6010
rect 20130 5958 20142 6010
rect 20142 5958 20172 6010
rect 20196 5958 20206 6010
rect 20206 5958 20252 6010
rect 19956 5956 20012 5958
rect 20036 5956 20092 5958
rect 20116 5956 20172 5958
rect 20196 5956 20252 5958
rect 19798 5752 19854 5808
rect 20626 7656 20682 7712
rect 20718 7520 20774 7576
rect 20626 7112 20682 7168
rect 20534 6432 20590 6488
rect 19956 4922 20012 4924
rect 20036 4922 20092 4924
rect 20116 4922 20172 4924
rect 20196 4922 20252 4924
rect 19956 4870 20002 4922
rect 20002 4870 20012 4922
rect 20036 4870 20066 4922
rect 20066 4870 20078 4922
rect 20078 4870 20092 4922
rect 20116 4870 20130 4922
rect 20130 4870 20142 4922
rect 20142 4870 20172 4922
rect 20196 4870 20206 4922
rect 20206 4870 20252 4922
rect 19956 4868 20012 4870
rect 20036 4868 20092 4870
rect 20116 4868 20172 4870
rect 20196 4868 20252 4870
rect 19956 3834 20012 3836
rect 20036 3834 20092 3836
rect 20116 3834 20172 3836
rect 20196 3834 20252 3836
rect 19956 3782 20002 3834
rect 20002 3782 20012 3834
rect 20036 3782 20066 3834
rect 20066 3782 20078 3834
rect 20078 3782 20092 3834
rect 20116 3782 20130 3834
rect 20130 3782 20142 3834
rect 20142 3782 20172 3834
rect 20196 3782 20206 3834
rect 20206 3782 20252 3834
rect 19956 3780 20012 3782
rect 20036 3780 20092 3782
rect 20116 3780 20172 3782
rect 20196 3780 20252 3782
rect 20718 3440 20774 3496
rect 21016 8730 21072 8732
rect 21096 8730 21152 8732
rect 21176 8730 21232 8732
rect 21256 8730 21312 8732
rect 21016 8678 21062 8730
rect 21062 8678 21072 8730
rect 21096 8678 21126 8730
rect 21126 8678 21138 8730
rect 21138 8678 21152 8730
rect 21176 8678 21190 8730
rect 21190 8678 21202 8730
rect 21202 8678 21232 8730
rect 21256 8678 21266 8730
rect 21266 8678 21312 8730
rect 21016 8676 21072 8678
rect 21096 8676 21152 8678
rect 21176 8676 21232 8678
rect 21256 8676 21312 8678
rect 21016 7642 21072 7644
rect 21096 7642 21152 7644
rect 21176 7642 21232 7644
rect 21256 7642 21312 7644
rect 21016 7590 21062 7642
rect 21062 7590 21072 7642
rect 21096 7590 21126 7642
rect 21126 7590 21138 7642
rect 21138 7590 21152 7642
rect 21176 7590 21190 7642
rect 21190 7590 21202 7642
rect 21202 7590 21232 7642
rect 21256 7590 21266 7642
rect 21266 7590 21312 7642
rect 21016 7588 21072 7590
rect 21096 7588 21152 7590
rect 21176 7588 21232 7590
rect 21256 7588 21312 7590
rect 21016 6554 21072 6556
rect 21096 6554 21152 6556
rect 21176 6554 21232 6556
rect 21256 6554 21312 6556
rect 21016 6502 21062 6554
rect 21062 6502 21072 6554
rect 21096 6502 21126 6554
rect 21126 6502 21138 6554
rect 21138 6502 21152 6554
rect 21176 6502 21190 6554
rect 21190 6502 21202 6554
rect 21202 6502 21232 6554
rect 21256 6502 21266 6554
rect 21266 6502 21312 6554
rect 21016 6500 21072 6502
rect 21096 6500 21152 6502
rect 21176 6500 21232 6502
rect 21256 6500 21312 6502
rect 21016 5466 21072 5468
rect 21096 5466 21152 5468
rect 21176 5466 21232 5468
rect 21256 5466 21312 5468
rect 21016 5414 21062 5466
rect 21062 5414 21072 5466
rect 21096 5414 21126 5466
rect 21126 5414 21138 5466
rect 21138 5414 21152 5466
rect 21176 5414 21190 5466
rect 21190 5414 21202 5466
rect 21202 5414 21232 5466
rect 21256 5414 21266 5466
rect 21266 5414 21312 5466
rect 21016 5412 21072 5414
rect 21096 5412 21152 5414
rect 21176 5412 21232 5414
rect 21256 5412 21312 5414
rect 21016 4378 21072 4380
rect 21096 4378 21152 4380
rect 21176 4378 21232 4380
rect 21256 4378 21312 4380
rect 21016 4326 21062 4378
rect 21062 4326 21072 4378
rect 21096 4326 21126 4378
rect 21126 4326 21138 4378
rect 21138 4326 21152 4378
rect 21176 4326 21190 4378
rect 21190 4326 21202 4378
rect 21202 4326 21232 4378
rect 21256 4326 21266 4378
rect 21266 4326 21312 4378
rect 21016 4324 21072 4326
rect 21096 4324 21152 4326
rect 21176 4324 21232 4326
rect 21256 4324 21312 4326
rect 22190 6296 22246 6352
rect 21016 3290 21072 3292
rect 21096 3290 21152 3292
rect 21176 3290 21232 3292
rect 21256 3290 21312 3292
rect 21016 3238 21062 3290
rect 21062 3238 21072 3290
rect 21096 3238 21126 3290
rect 21126 3238 21138 3290
rect 21138 3238 21152 3290
rect 21176 3238 21190 3290
rect 21190 3238 21202 3290
rect 21202 3238 21232 3290
rect 21256 3238 21266 3290
rect 21266 3238 21312 3290
rect 21016 3236 21072 3238
rect 21096 3236 21152 3238
rect 21176 3236 21232 3238
rect 21256 3236 21312 3238
rect 9402 2896 9458 2952
rect 9494 2488 9550 2544
rect 9016 2202 9072 2204
rect 9096 2202 9152 2204
rect 9176 2202 9232 2204
rect 9256 2202 9312 2204
rect 9016 2150 9062 2202
rect 9062 2150 9072 2202
rect 9096 2150 9126 2202
rect 9126 2150 9138 2202
rect 9138 2150 9152 2202
rect 9176 2150 9190 2202
rect 9190 2150 9202 2202
rect 9202 2150 9232 2202
rect 9256 2150 9266 2202
rect 9266 2150 9312 2202
rect 9016 2148 9072 2150
rect 9096 2148 9152 2150
rect 9176 2148 9232 2150
rect 9256 2148 9312 2150
rect 17222 3032 17278 3088
rect 9586 1672 9642 1728
rect 11058 2932 11060 2952
rect 11060 2932 11112 2952
rect 11112 2932 11114 2952
rect 11058 2896 11114 2932
rect 13956 2746 14012 2748
rect 14036 2746 14092 2748
rect 14116 2746 14172 2748
rect 14196 2746 14252 2748
rect 13956 2694 14002 2746
rect 14002 2694 14012 2746
rect 14036 2694 14066 2746
rect 14066 2694 14078 2746
rect 14078 2694 14092 2746
rect 14116 2694 14130 2746
rect 14130 2694 14142 2746
rect 14142 2694 14172 2746
rect 14196 2694 14206 2746
rect 14206 2694 14252 2746
rect 13956 2692 14012 2694
rect 14036 2692 14092 2694
rect 14116 2692 14172 2694
rect 14196 2692 14252 2694
rect 15016 2202 15072 2204
rect 15096 2202 15152 2204
rect 15176 2202 15232 2204
rect 15256 2202 15312 2204
rect 15016 2150 15062 2202
rect 15062 2150 15072 2202
rect 15096 2150 15126 2202
rect 15126 2150 15138 2202
rect 15138 2150 15152 2202
rect 15176 2150 15190 2202
rect 15190 2150 15202 2202
rect 15202 2150 15232 2202
rect 15256 2150 15266 2202
rect 15266 2150 15312 2202
rect 15016 2148 15072 2150
rect 15096 2148 15152 2150
rect 15176 2148 15232 2150
rect 15256 2148 15312 2150
rect 19706 1944 19762 2000
rect 19956 2746 20012 2748
rect 20036 2746 20092 2748
rect 20116 2746 20172 2748
rect 20196 2746 20252 2748
rect 19956 2694 20002 2746
rect 20002 2694 20012 2746
rect 20036 2694 20066 2746
rect 20066 2694 20078 2746
rect 20078 2694 20092 2746
rect 20116 2694 20130 2746
rect 20130 2694 20142 2746
rect 20142 2694 20172 2746
rect 20196 2694 20206 2746
rect 20206 2694 20252 2746
rect 19956 2692 20012 2694
rect 20036 2692 20092 2694
rect 20116 2692 20172 2694
rect 20196 2692 20252 2694
rect 20718 2352 20774 2408
rect 21016 2202 21072 2204
rect 21096 2202 21152 2204
rect 21176 2202 21232 2204
rect 21256 2202 21312 2204
rect 21016 2150 21062 2202
rect 21062 2150 21072 2202
rect 21096 2150 21126 2202
rect 21126 2150 21138 2202
rect 21138 2150 21152 2202
rect 21176 2150 21190 2202
rect 21190 2150 21202 2202
rect 21202 2150 21232 2202
rect 21256 2150 21266 2202
rect 21266 2150 21312 2202
rect 21016 2148 21072 2150
rect 21096 2148 21152 2150
rect 21176 2148 21232 2150
rect 21256 2148 21312 2150
rect 22742 6976 22798 7032
rect 25956 8186 26012 8188
rect 26036 8186 26092 8188
rect 26116 8186 26172 8188
rect 26196 8186 26252 8188
rect 25956 8134 26002 8186
rect 26002 8134 26012 8186
rect 26036 8134 26066 8186
rect 26066 8134 26078 8186
rect 26078 8134 26092 8186
rect 26116 8134 26130 8186
rect 26130 8134 26142 8186
rect 26142 8134 26172 8186
rect 26196 8134 26206 8186
rect 26206 8134 26252 8186
rect 25956 8132 26012 8134
rect 26036 8132 26092 8134
rect 26116 8132 26172 8134
rect 26196 8132 26252 8134
rect 27016 8730 27072 8732
rect 27096 8730 27152 8732
rect 27176 8730 27232 8732
rect 27256 8730 27312 8732
rect 27016 8678 27062 8730
rect 27062 8678 27072 8730
rect 27096 8678 27126 8730
rect 27126 8678 27138 8730
rect 27138 8678 27152 8730
rect 27176 8678 27190 8730
rect 27190 8678 27202 8730
rect 27202 8678 27232 8730
rect 27256 8678 27266 8730
rect 27266 8678 27312 8730
rect 27016 8676 27072 8678
rect 27096 8676 27152 8678
rect 27176 8676 27232 8678
rect 27256 8676 27312 8678
rect 27016 7642 27072 7644
rect 27096 7642 27152 7644
rect 27176 7642 27232 7644
rect 27256 7642 27312 7644
rect 27016 7590 27062 7642
rect 27062 7590 27072 7642
rect 27096 7590 27126 7642
rect 27126 7590 27138 7642
rect 27138 7590 27152 7642
rect 27176 7590 27190 7642
rect 27190 7590 27202 7642
rect 27202 7590 27232 7642
rect 27256 7590 27266 7642
rect 27266 7590 27312 7642
rect 27016 7588 27072 7590
rect 27096 7588 27152 7590
rect 27176 7588 27232 7590
rect 27256 7588 27312 7590
rect 28814 10920 28870 10976
rect 28446 10784 28502 10840
rect 28078 7248 28134 7304
rect 25956 7098 26012 7100
rect 26036 7098 26092 7100
rect 26116 7098 26172 7100
rect 26196 7098 26252 7100
rect 25956 7046 26002 7098
rect 26002 7046 26012 7098
rect 26036 7046 26066 7098
rect 26066 7046 26078 7098
rect 26078 7046 26092 7098
rect 26116 7046 26130 7098
rect 26130 7046 26142 7098
rect 26142 7046 26172 7098
rect 26196 7046 26206 7098
rect 26206 7046 26252 7098
rect 25956 7044 26012 7046
rect 26036 7044 26092 7046
rect 26116 7044 26172 7046
rect 26196 7044 26252 7046
rect 27016 6554 27072 6556
rect 27096 6554 27152 6556
rect 27176 6554 27232 6556
rect 27256 6554 27312 6556
rect 27016 6502 27062 6554
rect 27062 6502 27072 6554
rect 27096 6502 27126 6554
rect 27126 6502 27138 6554
rect 27138 6502 27152 6554
rect 27176 6502 27190 6554
rect 27190 6502 27202 6554
rect 27202 6502 27232 6554
rect 27256 6502 27266 6554
rect 27266 6502 27312 6554
rect 27016 6500 27072 6502
rect 27096 6500 27152 6502
rect 27176 6500 27232 6502
rect 27256 6500 27312 6502
rect 25956 6010 26012 6012
rect 26036 6010 26092 6012
rect 26116 6010 26172 6012
rect 26196 6010 26252 6012
rect 25956 5958 26002 6010
rect 26002 5958 26012 6010
rect 26036 5958 26066 6010
rect 26066 5958 26078 6010
rect 26078 5958 26092 6010
rect 26116 5958 26130 6010
rect 26130 5958 26142 6010
rect 26142 5958 26172 6010
rect 26196 5958 26206 6010
rect 26206 5958 26252 6010
rect 25956 5956 26012 5958
rect 26036 5956 26092 5958
rect 26116 5956 26172 5958
rect 26196 5956 26252 5958
rect 25956 4922 26012 4924
rect 26036 4922 26092 4924
rect 26116 4922 26172 4924
rect 26196 4922 26252 4924
rect 25956 4870 26002 4922
rect 26002 4870 26012 4922
rect 26036 4870 26066 4922
rect 26066 4870 26078 4922
rect 26078 4870 26092 4922
rect 26116 4870 26130 4922
rect 26130 4870 26142 4922
rect 26142 4870 26172 4922
rect 26196 4870 26206 4922
rect 26206 4870 26252 4922
rect 25956 4868 26012 4870
rect 26036 4868 26092 4870
rect 26116 4868 26172 4870
rect 26196 4868 26252 4870
rect 24674 4120 24730 4176
rect 24766 3984 24822 4040
rect 24858 3576 24914 3632
rect 25956 3834 26012 3836
rect 26036 3834 26092 3836
rect 26116 3834 26172 3836
rect 26196 3834 26252 3836
rect 25956 3782 26002 3834
rect 26002 3782 26012 3834
rect 26036 3782 26066 3834
rect 26066 3782 26078 3834
rect 26078 3782 26092 3834
rect 26116 3782 26130 3834
rect 26130 3782 26142 3834
rect 26142 3782 26172 3834
rect 26196 3782 26206 3834
rect 26206 3782 26252 3834
rect 25956 3780 26012 3782
rect 26036 3780 26092 3782
rect 26116 3780 26172 3782
rect 26196 3780 26252 3782
rect 25870 3440 25926 3496
rect 27016 5466 27072 5468
rect 27096 5466 27152 5468
rect 27176 5466 27232 5468
rect 27256 5466 27312 5468
rect 27016 5414 27062 5466
rect 27062 5414 27072 5466
rect 27096 5414 27126 5466
rect 27126 5414 27138 5466
rect 27138 5414 27152 5466
rect 27176 5414 27190 5466
rect 27190 5414 27202 5466
rect 27202 5414 27232 5466
rect 27256 5414 27266 5466
rect 27266 5414 27312 5466
rect 27016 5412 27072 5414
rect 27096 5412 27152 5414
rect 27176 5412 27232 5414
rect 27256 5412 27312 5414
rect 27016 4378 27072 4380
rect 27096 4378 27152 4380
rect 27176 4378 27232 4380
rect 27256 4378 27312 4380
rect 27016 4326 27062 4378
rect 27062 4326 27072 4378
rect 27096 4326 27126 4378
rect 27126 4326 27138 4378
rect 27138 4326 27152 4378
rect 27176 4326 27190 4378
rect 27190 4326 27202 4378
rect 27202 4326 27232 4378
rect 27256 4326 27266 4378
rect 27266 4326 27312 4378
rect 27016 4324 27072 4326
rect 27096 4324 27152 4326
rect 27176 4324 27232 4326
rect 27256 4324 27312 4326
rect 28998 3576 29054 3632
rect 30194 9016 30250 9072
rect 31956 8186 32012 8188
rect 32036 8186 32092 8188
rect 32116 8186 32172 8188
rect 32196 8186 32252 8188
rect 31956 8134 32002 8186
rect 32002 8134 32012 8186
rect 32036 8134 32066 8186
rect 32066 8134 32078 8186
rect 32078 8134 32092 8186
rect 32116 8134 32130 8186
rect 32130 8134 32142 8186
rect 32142 8134 32172 8186
rect 32196 8134 32206 8186
rect 32206 8134 32252 8186
rect 31956 8132 32012 8134
rect 32036 8132 32092 8134
rect 32116 8132 32172 8134
rect 32196 8132 32252 8134
rect 31956 7098 32012 7100
rect 32036 7098 32092 7100
rect 32116 7098 32172 7100
rect 32196 7098 32252 7100
rect 31956 7046 32002 7098
rect 32002 7046 32012 7098
rect 32036 7046 32066 7098
rect 32066 7046 32078 7098
rect 32078 7046 32092 7098
rect 32116 7046 32130 7098
rect 32130 7046 32142 7098
rect 32142 7046 32172 7098
rect 32196 7046 32206 7098
rect 32206 7046 32252 7098
rect 31956 7044 32012 7046
rect 32036 7044 32092 7046
rect 32116 7044 32172 7046
rect 32196 7044 32252 7046
rect 33016 8730 33072 8732
rect 33096 8730 33152 8732
rect 33176 8730 33232 8732
rect 33256 8730 33312 8732
rect 33016 8678 33062 8730
rect 33062 8678 33072 8730
rect 33096 8678 33126 8730
rect 33126 8678 33138 8730
rect 33138 8678 33152 8730
rect 33176 8678 33190 8730
rect 33190 8678 33202 8730
rect 33202 8678 33232 8730
rect 33256 8678 33266 8730
rect 33266 8678 33312 8730
rect 33016 8676 33072 8678
rect 33096 8676 33152 8678
rect 33176 8676 33232 8678
rect 33256 8676 33312 8678
rect 33016 7642 33072 7644
rect 33096 7642 33152 7644
rect 33176 7642 33232 7644
rect 33256 7642 33312 7644
rect 33016 7590 33062 7642
rect 33062 7590 33072 7642
rect 33096 7590 33126 7642
rect 33126 7590 33138 7642
rect 33138 7590 33152 7642
rect 33176 7590 33190 7642
rect 33190 7590 33202 7642
rect 33202 7590 33232 7642
rect 33256 7590 33266 7642
rect 33266 7590 33312 7642
rect 33016 7588 33072 7590
rect 33096 7588 33152 7590
rect 33176 7588 33232 7590
rect 33256 7588 33312 7590
rect 31956 6010 32012 6012
rect 32036 6010 32092 6012
rect 32116 6010 32172 6012
rect 32196 6010 32252 6012
rect 31956 5958 32002 6010
rect 32002 5958 32012 6010
rect 32036 5958 32066 6010
rect 32066 5958 32078 6010
rect 32078 5958 32092 6010
rect 32116 5958 32130 6010
rect 32130 5958 32142 6010
rect 32142 5958 32172 6010
rect 32196 5958 32206 6010
rect 32206 5958 32252 6010
rect 31956 5956 32012 5958
rect 32036 5956 32092 5958
rect 32116 5956 32172 5958
rect 32196 5956 32252 5958
rect 33016 6554 33072 6556
rect 33096 6554 33152 6556
rect 33176 6554 33232 6556
rect 33256 6554 33312 6556
rect 33016 6502 33062 6554
rect 33062 6502 33072 6554
rect 33096 6502 33126 6554
rect 33126 6502 33138 6554
rect 33138 6502 33152 6554
rect 33176 6502 33190 6554
rect 33190 6502 33202 6554
rect 33202 6502 33232 6554
rect 33256 6502 33266 6554
rect 33266 6502 33312 6554
rect 33016 6500 33072 6502
rect 33096 6500 33152 6502
rect 33176 6500 33232 6502
rect 33256 6500 33312 6502
rect 33016 5466 33072 5468
rect 33096 5466 33152 5468
rect 33176 5466 33232 5468
rect 33256 5466 33312 5468
rect 33016 5414 33062 5466
rect 33062 5414 33072 5466
rect 33096 5414 33126 5466
rect 33126 5414 33138 5466
rect 33138 5414 33152 5466
rect 33176 5414 33190 5466
rect 33190 5414 33202 5466
rect 33202 5414 33232 5466
rect 33256 5414 33266 5466
rect 33266 5414 33312 5466
rect 33016 5412 33072 5414
rect 33096 5412 33152 5414
rect 33176 5412 33232 5414
rect 33256 5412 33312 5414
rect 32770 5208 32826 5264
rect 34426 9832 34482 9888
rect 35438 9288 35494 9344
rect 35806 9152 35862 9208
rect 37278 11056 37334 11112
rect 37646 10648 37702 10704
rect 37278 9424 37334 9480
rect 36450 8880 36506 8936
rect 35346 6704 35402 6760
rect 31956 4922 32012 4924
rect 32036 4922 32092 4924
rect 32116 4922 32172 4924
rect 32196 4922 32252 4924
rect 31956 4870 32002 4922
rect 32002 4870 32012 4922
rect 32036 4870 32066 4922
rect 32066 4870 32078 4922
rect 32078 4870 32092 4922
rect 32116 4870 32130 4922
rect 32130 4870 32142 4922
rect 32142 4870 32172 4922
rect 32196 4870 32206 4922
rect 32206 4870 32252 4922
rect 31956 4868 32012 4870
rect 32036 4868 32092 4870
rect 32116 4868 32172 4870
rect 32196 4868 32252 4870
rect 33016 4378 33072 4380
rect 33096 4378 33152 4380
rect 33176 4378 33232 4380
rect 33256 4378 33312 4380
rect 33016 4326 33062 4378
rect 33062 4326 33072 4378
rect 33096 4326 33126 4378
rect 33126 4326 33138 4378
rect 33138 4326 33152 4378
rect 33176 4326 33190 4378
rect 33190 4326 33202 4378
rect 33202 4326 33232 4378
rect 33256 4326 33266 4378
rect 33266 4326 33312 4378
rect 33016 4324 33072 4326
rect 33096 4324 33152 4326
rect 33176 4324 33232 4326
rect 33256 4324 33312 4326
rect 31956 3834 32012 3836
rect 32036 3834 32092 3836
rect 32116 3834 32172 3836
rect 32196 3834 32252 3836
rect 31956 3782 32002 3834
rect 32002 3782 32012 3834
rect 32036 3782 32066 3834
rect 32066 3782 32078 3834
rect 32078 3782 32092 3834
rect 32116 3782 32130 3834
rect 32130 3782 32142 3834
rect 32142 3782 32172 3834
rect 32196 3782 32206 3834
rect 32206 3782 32252 3834
rect 31956 3780 32012 3782
rect 32036 3780 32092 3782
rect 32116 3780 32172 3782
rect 32196 3780 32252 3782
rect 27016 3290 27072 3292
rect 27096 3290 27152 3292
rect 27176 3290 27232 3292
rect 27256 3290 27312 3292
rect 27016 3238 27062 3290
rect 27062 3238 27072 3290
rect 27096 3238 27126 3290
rect 27126 3238 27138 3290
rect 27138 3238 27152 3290
rect 27176 3238 27190 3290
rect 27190 3238 27202 3290
rect 27202 3238 27232 3290
rect 27256 3238 27266 3290
rect 27266 3238 27312 3290
rect 27016 3236 27072 3238
rect 27096 3236 27152 3238
rect 27176 3236 27232 3238
rect 27256 3236 27312 3238
rect 25956 2746 26012 2748
rect 26036 2746 26092 2748
rect 26116 2746 26172 2748
rect 26196 2746 26252 2748
rect 25956 2694 26002 2746
rect 26002 2694 26012 2746
rect 26036 2694 26066 2746
rect 26066 2694 26078 2746
rect 26078 2694 26092 2746
rect 26116 2694 26130 2746
rect 26130 2694 26142 2746
rect 26142 2694 26172 2746
rect 26196 2694 26206 2746
rect 26206 2694 26252 2746
rect 25956 2692 26012 2694
rect 26036 2692 26092 2694
rect 26116 2692 26172 2694
rect 26196 2692 26252 2694
rect 28538 3032 28594 3088
rect 27016 2202 27072 2204
rect 27096 2202 27152 2204
rect 27176 2202 27232 2204
rect 27256 2202 27312 2204
rect 27016 2150 27062 2202
rect 27062 2150 27072 2202
rect 27096 2150 27126 2202
rect 27126 2150 27138 2202
rect 27138 2150 27152 2202
rect 27176 2150 27190 2202
rect 27190 2150 27202 2202
rect 27202 2150 27232 2202
rect 27256 2150 27266 2202
rect 27266 2150 27312 2202
rect 27016 2148 27072 2150
rect 27096 2148 27152 2150
rect 27176 2148 27232 2150
rect 27256 2148 27312 2150
rect 33016 3290 33072 3292
rect 33096 3290 33152 3292
rect 33176 3290 33232 3292
rect 33256 3290 33312 3292
rect 33016 3238 33062 3290
rect 33062 3238 33072 3290
rect 33096 3238 33126 3290
rect 33126 3238 33138 3290
rect 33138 3238 33152 3290
rect 33176 3238 33190 3290
rect 33190 3238 33202 3290
rect 33202 3238 33232 3290
rect 33256 3238 33266 3290
rect 33266 3238 33312 3290
rect 33016 3236 33072 3238
rect 33096 3236 33152 3238
rect 33176 3236 33232 3238
rect 33256 3236 33312 3238
rect 31956 2746 32012 2748
rect 32036 2746 32092 2748
rect 32116 2746 32172 2748
rect 32196 2746 32252 2748
rect 31956 2694 32002 2746
rect 32002 2694 32012 2746
rect 32036 2694 32066 2746
rect 32066 2694 32078 2746
rect 32078 2694 32092 2746
rect 32116 2694 32130 2746
rect 32130 2694 32142 2746
rect 32142 2694 32172 2746
rect 32196 2694 32206 2746
rect 32206 2694 32252 2746
rect 31956 2692 32012 2694
rect 32036 2692 32092 2694
rect 32116 2692 32172 2694
rect 32196 2692 32252 2694
rect 33016 2202 33072 2204
rect 33096 2202 33152 2204
rect 33176 2202 33232 2204
rect 33256 2202 33312 2204
rect 33016 2150 33062 2202
rect 33062 2150 33072 2202
rect 33096 2150 33126 2202
rect 33126 2150 33138 2202
rect 33138 2150 33152 2202
rect 33176 2150 33190 2202
rect 33190 2150 33202 2202
rect 33202 2150 33232 2202
rect 33256 2150 33266 2202
rect 33266 2150 33312 2202
rect 33016 2148 33072 2150
rect 33096 2148 33152 2150
rect 33176 2148 33232 2150
rect 33256 2148 33312 2150
rect 36174 6180 36230 6216
rect 36174 6160 36176 6180
rect 36176 6160 36228 6180
rect 36228 6160 36230 6180
rect 39016 8730 39072 8732
rect 39096 8730 39152 8732
rect 39176 8730 39232 8732
rect 39256 8730 39312 8732
rect 39016 8678 39062 8730
rect 39062 8678 39072 8730
rect 39096 8678 39126 8730
rect 39126 8678 39138 8730
rect 39138 8678 39152 8730
rect 39176 8678 39190 8730
rect 39190 8678 39202 8730
rect 39202 8678 39232 8730
rect 39256 8678 39266 8730
rect 39266 8678 39312 8730
rect 39016 8676 39072 8678
rect 39096 8676 39152 8678
rect 39176 8676 39232 8678
rect 39256 8676 39312 8678
rect 37956 8186 38012 8188
rect 38036 8186 38092 8188
rect 38116 8186 38172 8188
rect 38196 8186 38252 8188
rect 37956 8134 38002 8186
rect 38002 8134 38012 8186
rect 38036 8134 38066 8186
rect 38066 8134 38078 8186
rect 38078 8134 38092 8186
rect 38116 8134 38130 8186
rect 38130 8134 38142 8186
rect 38142 8134 38172 8186
rect 38196 8134 38206 8186
rect 38206 8134 38252 8186
rect 37956 8132 38012 8134
rect 38036 8132 38092 8134
rect 38116 8132 38172 8134
rect 38196 8132 38252 8134
rect 37830 7384 37886 7440
rect 37956 7098 38012 7100
rect 38036 7098 38092 7100
rect 38116 7098 38172 7100
rect 38196 7098 38252 7100
rect 37956 7046 38002 7098
rect 38002 7046 38012 7098
rect 38036 7046 38066 7098
rect 38066 7046 38078 7098
rect 38078 7046 38092 7098
rect 38116 7046 38130 7098
rect 38130 7046 38142 7098
rect 38142 7046 38172 7098
rect 38196 7046 38206 7098
rect 38206 7046 38252 7098
rect 37956 7044 38012 7046
rect 38036 7044 38092 7046
rect 38116 7044 38172 7046
rect 38196 7044 38252 7046
rect 37956 6010 38012 6012
rect 38036 6010 38092 6012
rect 38116 6010 38172 6012
rect 38196 6010 38252 6012
rect 37956 5958 38002 6010
rect 38002 5958 38012 6010
rect 38036 5958 38066 6010
rect 38066 5958 38078 6010
rect 38078 5958 38092 6010
rect 38116 5958 38130 6010
rect 38130 5958 38142 6010
rect 38142 5958 38172 6010
rect 38196 5958 38206 6010
rect 38206 5958 38252 6010
rect 37956 5956 38012 5958
rect 38036 5956 38092 5958
rect 38116 5956 38172 5958
rect 38196 5956 38252 5958
rect 37554 5108 37556 5128
rect 37556 5108 37608 5128
rect 37608 5108 37610 5128
rect 37554 5072 37610 5108
rect 37956 4922 38012 4924
rect 38036 4922 38092 4924
rect 38116 4922 38172 4924
rect 38196 4922 38252 4924
rect 37956 4870 38002 4922
rect 38002 4870 38012 4922
rect 38036 4870 38066 4922
rect 38066 4870 38078 4922
rect 38078 4870 38092 4922
rect 38116 4870 38130 4922
rect 38130 4870 38142 4922
rect 38142 4870 38172 4922
rect 38196 4870 38206 4922
rect 38206 4870 38252 4922
rect 37956 4868 38012 4870
rect 38036 4868 38092 4870
rect 38116 4868 38172 4870
rect 38196 4868 38252 4870
rect 37956 3834 38012 3836
rect 38036 3834 38092 3836
rect 38116 3834 38172 3836
rect 38196 3834 38252 3836
rect 37956 3782 38002 3834
rect 38002 3782 38012 3834
rect 38036 3782 38066 3834
rect 38066 3782 38078 3834
rect 38078 3782 38092 3834
rect 38116 3782 38130 3834
rect 38130 3782 38142 3834
rect 38142 3782 38172 3834
rect 38196 3782 38206 3834
rect 38206 3782 38252 3834
rect 37956 3780 38012 3782
rect 38036 3780 38092 3782
rect 38116 3780 38172 3782
rect 38196 3780 38252 3782
rect 37956 2746 38012 2748
rect 38036 2746 38092 2748
rect 38116 2746 38172 2748
rect 38196 2746 38252 2748
rect 37956 2694 38002 2746
rect 38002 2694 38012 2746
rect 38036 2694 38066 2746
rect 38066 2694 38078 2746
rect 38078 2694 38092 2746
rect 38116 2694 38130 2746
rect 38130 2694 38142 2746
rect 38142 2694 38172 2746
rect 38196 2694 38206 2746
rect 38206 2694 38252 2746
rect 37956 2692 38012 2694
rect 38036 2692 38092 2694
rect 38116 2692 38172 2694
rect 38196 2692 38252 2694
rect 39016 7642 39072 7644
rect 39096 7642 39152 7644
rect 39176 7642 39232 7644
rect 39256 7642 39312 7644
rect 39016 7590 39062 7642
rect 39062 7590 39072 7642
rect 39096 7590 39126 7642
rect 39126 7590 39138 7642
rect 39138 7590 39152 7642
rect 39176 7590 39190 7642
rect 39190 7590 39202 7642
rect 39202 7590 39232 7642
rect 39256 7590 39266 7642
rect 39266 7590 39312 7642
rect 39016 7588 39072 7590
rect 39096 7588 39152 7590
rect 39176 7588 39232 7590
rect 39256 7588 39312 7590
rect 39016 6554 39072 6556
rect 39096 6554 39152 6556
rect 39176 6554 39232 6556
rect 39256 6554 39312 6556
rect 39016 6502 39062 6554
rect 39062 6502 39072 6554
rect 39096 6502 39126 6554
rect 39126 6502 39138 6554
rect 39138 6502 39152 6554
rect 39176 6502 39190 6554
rect 39190 6502 39202 6554
rect 39202 6502 39232 6554
rect 39256 6502 39266 6554
rect 39266 6502 39312 6554
rect 39016 6500 39072 6502
rect 39096 6500 39152 6502
rect 39176 6500 39232 6502
rect 39256 6500 39312 6502
rect 39016 5466 39072 5468
rect 39096 5466 39152 5468
rect 39176 5466 39232 5468
rect 39256 5466 39312 5468
rect 39016 5414 39062 5466
rect 39062 5414 39072 5466
rect 39096 5414 39126 5466
rect 39126 5414 39138 5466
rect 39138 5414 39152 5466
rect 39176 5414 39190 5466
rect 39190 5414 39202 5466
rect 39202 5414 39232 5466
rect 39256 5414 39266 5466
rect 39266 5414 39312 5466
rect 39016 5412 39072 5414
rect 39096 5412 39152 5414
rect 39176 5412 39232 5414
rect 39256 5412 39312 5414
rect 39016 4378 39072 4380
rect 39096 4378 39152 4380
rect 39176 4378 39232 4380
rect 39256 4378 39312 4380
rect 39016 4326 39062 4378
rect 39062 4326 39072 4378
rect 39096 4326 39126 4378
rect 39126 4326 39138 4378
rect 39138 4326 39152 4378
rect 39176 4326 39190 4378
rect 39190 4326 39202 4378
rect 39202 4326 39232 4378
rect 39256 4326 39266 4378
rect 39266 4326 39312 4378
rect 39016 4324 39072 4326
rect 39096 4324 39152 4326
rect 39176 4324 39232 4326
rect 39256 4324 39312 4326
rect 39016 3290 39072 3292
rect 39096 3290 39152 3292
rect 39176 3290 39232 3292
rect 39256 3290 39312 3292
rect 39016 3238 39062 3290
rect 39062 3238 39072 3290
rect 39096 3238 39126 3290
rect 39126 3238 39138 3290
rect 39138 3238 39152 3290
rect 39176 3238 39190 3290
rect 39190 3238 39202 3290
rect 39202 3238 39232 3290
rect 39256 3238 39266 3290
rect 39266 3238 39312 3290
rect 39016 3236 39072 3238
rect 39096 3236 39152 3238
rect 39176 3236 39232 3238
rect 39256 3236 39312 3238
rect 39016 2202 39072 2204
rect 39096 2202 39152 2204
rect 39176 2202 39232 2204
rect 39256 2202 39312 2204
rect 39016 2150 39062 2202
rect 39062 2150 39072 2202
rect 39096 2150 39126 2202
rect 39126 2150 39138 2202
rect 39138 2150 39152 2202
rect 39176 2150 39190 2202
rect 39190 2150 39202 2202
rect 39202 2150 39232 2202
rect 39256 2150 39266 2202
rect 39266 2150 39312 2202
rect 39016 2148 39072 2150
rect 39096 2148 39152 2150
rect 39176 2148 39232 2150
rect 39256 2148 39312 2150
rect 41602 8472 41658 8528
rect 41602 3576 41658 3632
rect 41418 2896 41474 2952
rect 42154 2488 42210 2544
rect 44822 9560 44878 9616
rect 43956 8186 44012 8188
rect 44036 8186 44092 8188
rect 44116 8186 44172 8188
rect 44196 8186 44252 8188
rect 43956 8134 44002 8186
rect 44002 8134 44012 8186
rect 44036 8134 44066 8186
rect 44066 8134 44078 8186
rect 44078 8134 44092 8186
rect 44116 8134 44130 8186
rect 44130 8134 44142 8186
rect 44142 8134 44172 8186
rect 44196 8134 44206 8186
rect 44206 8134 44252 8186
rect 43956 8132 44012 8134
rect 44036 8132 44092 8134
rect 44116 8132 44172 8134
rect 44196 8132 44252 8134
rect 45926 9288 45982 9344
rect 45016 8730 45072 8732
rect 45096 8730 45152 8732
rect 45176 8730 45232 8732
rect 45256 8730 45312 8732
rect 45016 8678 45062 8730
rect 45062 8678 45072 8730
rect 45096 8678 45126 8730
rect 45126 8678 45138 8730
rect 45138 8678 45152 8730
rect 45176 8678 45190 8730
rect 45190 8678 45202 8730
rect 45202 8678 45232 8730
rect 45256 8678 45266 8730
rect 45266 8678 45312 8730
rect 45016 8676 45072 8678
rect 45096 8676 45152 8678
rect 45176 8676 45232 8678
rect 45256 8676 45312 8678
rect 45098 7928 45154 7984
rect 45016 7642 45072 7644
rect 45096 7642 45152 7644
rect 45176 7642 45232 7644
rect 45256 7642 45312 7644
rect 45016 7590 45062 7642
rect 45062 7590 45072 7642
rect 45096 7590 45126 7642
rect 45126 7590 45138 7642
rect 45138 7590 45152 7642
rect 45176 7590 45190 7642
rect 45190 7590 45202 7642
rect 45202 7590 45232 7642
rect 45256 7590 45266 7642
rect 45266 7590 45312 7642
rect 45016 7588 45072 7590
rect 45096 7588 45152 7590
rect 45176 7588 45232 7590
rect 45256 7588 45312 7590
rect 43956 7098 44012 7100
rect 44036 7098 44092 7100
rect 44116 7098 44172 7100
rect 44196 7098 44252 7100
rect 43956 7046 44002 7098
rect 44002 7046 44012 7098
rect 44036 7046 44066 7098
rect 44066 7046 44078 7098
rect 44078 7046 44092 7098
rect 44116 7046 44130 7098
rect 44130 7046 44142 7098
rect 44142 7046 44172 7098
rect 44196 7046 44206 7098
rect 44206 7046 44252 7098
rect 43956 7044 44012 7046
rect 44036 7044 44092 7046
rect 44116 7044 44172 7046
rect 44196 7044 44252 7046
rect 45016 6554 45072 6556
rect 45096 6554 45152 6556
rect 45176 6554 45232 6556
rect 45256 6554 45312 6556
rect 45016 6502 45062 6554
rect 45062 6502 45072 6554
rect 45096 6502 45126 6554
rect 45126 6502 45138 6554
rect 45138 6502 45152 6554
rect 45176 6502 45190 6554
rect 45190 6502 45202 6554
rect 45202 6502 45232 6554
rect 45256 6502 45266 6554
rect 45266 6502 45312 6554
rect 45016 6500 45072 6502
rect 45096 6500 45152 6502
rect 45176 6500 45232 6502
rect 45256 6500 45312 6502
rect 43956 6010 44012 6012
rect 44036 6010 44092 6012
rect 44116 6010 44172 6012
rect 44196 6010 44252 6012
rect 43956 5958 44002 6010
rect 44002 5958 44012 6010
rect 44036 5958 44066 6010
rect 44066 5958 44078 6010
rect 44078 5958 44092 6010
rect 44116 5958 44130 6010
rect 44130 5958 44142 6010
rect 44142 5958 44172 6010
rect 44196 5958 44206 6010
rect 44206 5958 44252 6010
rect 43956 5956 44012 5958
rect 44036 5956 44092 5958
rect 44116 5956 44172 5958
rect 44196 5956 44252 5958
rect 43956 4922 44012 4924
rect 44036 4922 44092 4924
rect 44116 4922 44172 4924
rect 44196 4922 44252 4924
rect 43956 4870 44002 4922
rect 44002 4870 44012 4922
rect 44036 4870 44066 4922
rect 44066 4870 44078 4922
rect 44078 4870 44092 4922
rect 44116 4870 44130 4922
rect 44130 4870 44142 4922
rect 44142 4870 44172 4922
rect 44196 4870 44206 4922
rect 44206 4870 44252 4922
rect 43956 4868 44012 4870
rect 44036 4868 44092 4870
rect 44116 4868 44172 4870
rect 44196 4868 44252 4870
rect 43956 3834 44012 3836
rect 44036 3834 44092 3836
rect 44116 3834 44172 3836
rect 44196 3834 44252 3836
rect 43956 3782 44002 3834
rect 44002 3782 44012 3834
rect 44036 3782 44066 3834
rect 44066 3782 44078 3834
rect 44078 3782 44092 3834
rect 44116 3782 44130 3834
rect 44130 3782 44142 3834
rect 44142 3782 44172 3834
rect 44196 3782 44206 3834
rect 44206 3782 44252 3834
rect 43956 3780 44012 3782
rect 44036 3780 44092 3782
rect 44116 3780 44172 3782
rect 44196 3780 44252 3782
rect 44178 3476 44180 3496
rect 44180 3476 44232 3496
rect 44232 3476 44234 3496
rect 44178 3440 44234 3476
rect 45016 5466 45072 5468
rect 45096 5466 45152 5468
rect 45176 5466 45232 5468
rect 45256 5466 45312 5468
rect 45016 5414 45062 5466
rect 45062 5414 45072 5466
rect 45096 5414 45126 5466
rect 45126 5414 45138 5466
rect 45138 5414 45152 5466
rect 45176 5414 45190 5466
rect 45190 5414 45202 5466
rect 45202 5414 45232 5466
rect 45256 5414 45266 5466
rect 45266 5414 45312 5466
rect 45016 5412 45072 5414
rect 45096 5412 45152 5414
rect 45176 5412 45232 5414
rect 45256 5412 45312 5414
rect 45016 4378 45072 4380
rect 45096 4378 45152 4380
rect 45176 4378 45232 4380
rect 45256 4378 45312 4380
rect 45016 4326 45062 4378
rect 45062 4326 45072 4378
rect 45096 4326 45126 4378
rect 45126 4326 45138 4378
rect 45138 4326 45152 4378
rect 45176 4326 45190 4378
rect 45190 4326 45202 4378
rect 45202 4326 45232 4378
rect 45256 4326 45266 4378
rect 45266 4326 45312 4378
rect 45016 4324 45072 4326
rect 45096 4324 45152 4326
rect 45176 4324 45232 4326
rect 45256 4324 45312 4326
rect 45016 3290 45072 3292
rect 45096 3290 45152 3292
rect 45176 3290 45232 3292
rect 45256 3290 45312 3292
rect 45016 3238 45062 3290
rect 45062 3238 45072 3290
rect 45096 3238 45126 3290
rect 45126 3238 45138 3290
rect 45138 3238 45152 3290
rect 45176 3238 45190 3290
rect 45190 3238 45202 3290
rect 45202 3238 45232 3290
rect 45256 3238 45266 3290
rect 45266 3238 45312 3290
rect 45016 3236 45072 3238
rect 45096 3236 45152 3238
rect 45176 3236 45232 3238
rect 45256 3236 45312 3238
rect 43956 2746 44012 2748
rect 44036 2746 44092 2748
rect 44116 2746 44172 2748
rect 44196 2746 44252 2748
rect 43956 2694 44002 2746
rect 44002 2694 44012 2746
rect 44036 2694 44066 2746
rect 44066 2694 44078 2746
rect 44078 2694 44092 2746
rect 44116 2694 44130 2746
rect 44130 2694 44142 2746
rect 44142 2694 44172 2746
rect 44196 2694 44206 2746
rect 44206 2694 44252 2746
rect 43956 2692 44012 2694
rect 44036 2692 44092 2694
rect 44116 2692 44172 2694
rect 44196 2692 44252 2694
rect 45016 2202 45072 2204
rect 45096 2202 45152 2204
rect 45176 2202 45232 2204
rect 45256 2202 45312 2204
rect 45016 2150 45062 2202
rect 45062 2150 45072 2202
rect 45096 2150 45126 2202
rect 45126 2150 45138 2202
rect 45138 2150 45152 2202
rect 45176 2150 45190 2202
rect 45190 2150 45202 2202
rect 45202 2150 45232 2202
rect 45256 2150 45266 2202
rect 45266 2150 45312 2202
rect 45016 2148 45072 2150
rect 45096 2148 45152 2150
rect 45176 2148 45232 2150
rect 45256 2148 45312 2150
rect 45650 9016 45706 9072
rect 45742 8336 45798 8392
rect 45650 7792 45706 7848
rect 46294 8744 46350 8800
rect 46018 7964 46020 7984
rect 46020 7964 46072 7984
rect 46072 7964 46074 7984
rect 46018 7928 46074 7964
rect 46570 8200 46626 8256
rect 47030 8472 47086 8528
rect 46938 7384 46994 7440
rect 46662 6840 46718 6896
rect 46294 6296 46350 6352
rect 46570 5752 46626 5808
rect 46110 5616 46166 5672
rect 47490 9832 47546 9888
rect 47306 7656 47362 7712
rect 46938 6568 46994 6624
rect 47030 5516 47032 5536
rect 47032 5516 47084 5536
rect 47084 5516 47086 5536
rect 47030 5480 47086 5516
rect 46938 4972 46940 4992
rect 46940 4972 46992 4992
rect 46992 4972 46994 4992
rect 46938 4936 46994 4972
rect 47030 4428 47032 4448
rect 47032 4428 47084 4448
rect 47084 4428 47086 4448
rect 47030 4392 47086 4428
rect 46938 3884 46940 3904
rect 46940 3884 46992 3904
rect 46992 3884 46994 3904
rect 46938 3848 46994 3884
rect 47030 3340 47032 3360
rect 47032 3340 47084 3360
rect 47084 3340 47086 3360
rect 47030 3304 47086 3340
rect 46754 3052 46810 3088
rect 46754 3032 46756 3052
rect 46756 3032 46808 3052
rect 46808 3032 46810 3052
rect 46938 2796 46940 2816
rect 46940 2796 46992 2816
rect 46992 2796 46994 2816
rect 46938 2760 46994 2796
rect 45650 2488 45706 2544
rect 46938 2252 46940 2272
rect 46940 2252 46992 2272
rect 46992 2252 46994 2272
rect 45834 1944 45890 2000
rect 46202 1672 46258 1728
rect 46938 2216 46994 2252
rect 46570 1400 46626 1456
rect 47398 7112 47454 7168
rect 47398 6024 47454 6080
rect 47306 5208 47362 5264
rect 47398 4700 47400 4720
rect 47400 4700 47452 4720
rect 47452 4700 47454 4720
rect 47398 4664 47454 4700
rect 47306 4120 47362 4176
rect 47398 3612 47400 3632
rect 47400 3612 47452 3632
rect 47452 3612 47454 3632
rect 47398 3576 47454 3612
rect 47306 3032 47362 3088
rect 47306 2524 47308 2544
rect 47308 2524 47360 2544
rect 47360 2524 47362 2544
rect 47306 2488 47362 2524
<< metal3 >>
rect 16389 11114 16455 11117
rect 37273 11114 37339 11117
rect 16389 11112 37339 11114
rect 16389 11056 16394 11112
rect 16450 11056 37278 11112
rect 37334 11056 37339 11112
rect 16389 11054 37339 11056
rect 16389 11051 16455 11054
rect 37273 11051 37339 11054
rect 10869 10978 10935 10981
rect 28809 10978 28875 10981
rect 10869 10976 28875 10978
rect 10869 10920 10874 10976
rect 10930 10920 28814 10976
rect 28870 10920 28875 10976
rect 10869 10918 28875 10920
rect 10869 10915 10935 10918
rect 28809 10915 28875 10918
rect 11973 10842 12039 10845
rect 28441 10842 28507 10845
rect 11973 10840 28507 10842
rect 11973 10784 11978 10840
rect 12034 10784 28446 10840
rect 28502 10784 28507 10840
rect 11973 10782 28507 10784
rect 11973 10779 12039 10782
rect 28441 10779 28507 10782
rect 16021 10706 16087 10709
rect 37641 10706 37707 10709
rect 16021 10704 37707 10706
rect 16021 10648 16026 10704
rect 16082 10648 37646 10704
rect 37702 10648 37707 10704
rect 16021 10646 37707 10648
rect 16021 10643 16087 10646
rect 37641 10643 37707 10646
rect 0 9890 120 9920
rect 34421 9890 34487 9893
rect 0 9888 34487 9890
rect 0 9832 34426 9888
rect 34482 9832 34487 9888
rect 0 9830 34487 9832
rect 0 9800 120 9830
rect 34421 9827 34487 9830
rect 47485 9890 47551 9893
rect 48880 9890 49000 9920
rect 47485 9888 49000 9890
rect 47485 9832 47490 9888
rect 47546 9832 49000 9888
rect 47485 9830 49000 9832
rect 47485 9827 47551 9830
rect 48880 9800 49000 9830
rect 19517 9754 19583 9757
rect 20713 9754 20779 9757
rect 19517 9752 20779 9754
rect 19517 9696 19522 9752
rect 19578 9696 20718 9752
rect 20774 9696 20779 9752
rect 19517 9694 20779 9696
rect 19517 9691 19583 9694
rect 20713 9691 20779 9694
rect 0 9618 120 9648
rect 5165 9618 5231 9621
rect 0 9616 5231 9618
rect 0 9560 5170 9616
rect 5226 9560 5231 9616
rect 0 9558 5231 9560
rect 0 9528 120 9558
rect 5165 9555 5231 9558
rect 44817 9618 44883 9621
rect 48880 9618 49000 9648
rect 44817 9616 49000 9618
rect 44817 9560 44822 9616
rect 44878 9560 49000 9616
rect 44817 9558 49000 9560
rect 44817 9555 44883 9558
rect 48880 9528 49000 9558
rect 1117 9482 1183 9485
rect 37273 9482 37339 9485
rect 1117 9480 37339 9482
rect 1117 9424 1122 9480
rect 1178 9424 37278 9480
rect 37334 9424 37339 9480
rect 1117 9422 37339 9424
rect 1117 9419 1183 9422
rect 37273 9419 37339 9422
rect 0 9346 120 9376
rect 197 9346 263 9349
rect 0 9344 263 9346
rect 0 9288 202 9344
rect 258 9288 263 9344
rect 0 9286 263 9288
rect 0 9256 120 9286
rect 197 9283 263 9286
rect 20437 9346 20503 9349
rect 35433 9346 35499 9349
rect 20437 9344 35499 9346
rect 20437 9288 20442 9344
rect 20498 9288 35438 9344
rect 35494 9288 35499 9344
rect 20437 9286 35499 9288
rect 20437 9283 20503 9286
rect 35433 9283 35499 9286
rect 45921 9346 45987 9349
rect 48880 9346 49000 9376
rect 45921 9344 49000 9346
rect 45921 9288 45926 9344
rect 45982 9288 49000 9344
rect 45921 9286 49000 9288
rect 45921 9283 45987 9286
rect 48880 9256 49000 9286
rect 19793 9210 19859 9213
rect 35801 9210 35867 9213
rect 19793 9208 35867 9210
rect 19793 9152 19798 9208
rect 19854 9152 35806 9208
rect 35862 9152 35867 9208
rect 19793 9150 35867 9152
rect 19793 9147 19859 9150
rect 35801 9147 35867 9150
rect 0 9074 120 9104
rect 30189 9074 30255 9077
rect 0 9072 30255 9074
rect 0 9016 30194 9072
rect 30250 9016 30255 9072
rect 0 9014 30255 9016
rect 0 8984 120 9014
rect 30189 9011 30255 9014
rect 45645 9074 45711 9077
rect 48880 9074 49000 9104
rect 45645 9072 49000 9074
rect 45645 9016 45650 9072
rect 45706 9016 49000 9072
rect 45645 9014 49000 9016
rect 45645 9011 45711 9014
rect 48880 8984 49000 9014
rect 7741 8938 7807 8941
rect 36445 8938 36511 8941
rect 2730 8936 7807 8938
rect 2730 8880 7746 8936
rect 7802 8880 7807 8936
rect 2730 8878 7807 8880
rect 0 8802 120 8832
rect 2730 8802 2790 8878
rect 7741 8875 7807 8878
rect 7974 8936 36511 8938
rect 7974 8880 36450 8936
rect 36506 8880 36511 8936
rect 7974 8878 36511 8880
rect 0 8742 2790 8802
rect 4613 8802 4679 8805
rect 7974 8802 8034 8878
rect 36445 8875 36511 8878
rect 4613 8800 8034 8802
rect 4613 8744 4618 8800
rect 4674 8744 8034 8800
rect 4613 8742 8034 8744
rect 46289 8802 46355 8805
rect 48880 8802 49000 8832
rect 46289 8800 49000 8802
rect 46289 8744 46294 8800
rect 46350 8744 49000 8800
rect 46289 8742 49000 8744
rect 0 8712 120 8742
rect 4613 8739 4679 8742
rect 46289 8739 46355 8742
rect 3006 8736 3322 8737
rect 3006 8672 3012 8736
rect 3076 8672 3092 8736
rect 3156 8672 3172 8736
rect 3236 8672 3252 8736
rect 3316 8672 3322 8736
rect 3006 8671 3322 8672
rect 9006 8736 9322 8737
rect 9006 8672 9012 8736
rect 9076 8672 9092 8736
rect 9156 8672 9172 8736
rect 9236 8672 9252 8736
rect 9316 8672 9322 8736
rect 9006 8671 9322 8672
rect 15006 8736 15322 8737
rect 15006 8672 15012 8736
rect 15076 8672 15092 8736
rect 15156 8672 15172 8736
rect 15236 8672 15252 8736
rect 15316 8672 15322 8736
rect 15006 8671 15322 8672
rect 21006 8736 21322 8737
rect 21006 8672 21012 8736
rect 21076 8672 21092 8736
rect 21156 8672 21172 8736
rect 21236 8672 21252 8736
rect 21316 8672 21322 8736
rect 21006 8671 21322 8672
rect 27006 8736 27322 8737
rect 27006 8672 27012 8736
rect 27076 8672 27092 8736
rect 27156 8672 27172 8736
rect 27236 8672 27252 8736
rect 27316 8672 27322 8736
rect 27006 8671 27322 8672
rect 33006 8736 33322 8737
rect 33006 8672 33012 8736
rect 33076 8672 33092 8736
rect 33156 8672 33172 8736
rect 33236 8672 33252 8736
rect 33316 8672 33322 8736
rect 33006 8671 33322 8672
rect 39006 8736 39322 8737
rect 39006 8672 39012 8736
rect 39076 8672 39092 8736
rect 39156 8672 39172 8736
rect 39236 8672 39252 8736
rect 39316 8672 39322 8736
rect 39006 8671 39322 8672
rect 45006 8736 45322 8737
rect 45006 8672 45012 8736
rect 45076 8672 45092 8736
rect 45156 8672 45172 8736
rect 45236 8672 45252 8736
rect 45316 8672 45322 8736
rect 48880 8712 49000 8742
rect 45006 8671 45322 8672
rect 0 8530 120 8560
rect 41597 8530 41663 8533
rect 0 8528 41663 8530
rect 0 8472 41602 8528
rect 41658 8472 41663 8528
rect 0 8470 41663 8472
rect 0 8440 120 8470
rect 41597 8467 41663 8470
rect 47025 8530 47091 8533
rect 48880 8530 49000 8560
rect 47025 8528 49000 8530
rect 47025 8472 47030 8528
rect 47086 8472 49000 8528
rect 47025 8470 49000 8472
rect 47025 8467 47091 8470
rect 48880 8440 49000 8470
rect 8293 8394 8359 8397
rect 45737 8394 45803 8397
rect 8293 8392 45803 8394
rect 8293 8336 8298 8392
rect 8354 8336 45742 8392
rect 45798 8336 45803 8392
rect 8293 8334 45803 8336
rect 8293 8331 8359 8334
rect 45737 8331 45803 8334
rect 0 8258 120 8288
rect 1301 8258 1367 8261
rect 0 8256 1367 8258
rect 0 8200 1306 8256
rect 1362 8200 1367 8256
rect 0 8198 1367 8200
rect 0 8168 120 8198
rect 1301 8195 1367 8198
rect 12433 8258 12499 8261
rect 12801 8258 12867 8261
rect 12433 8256 12867 8258
rect 12433 8200 12438 8256
rect 12494 8200 12806 8256
rect 12862 8200 12867 8256
rect 12433 8198 12867 8200
rect 12433 8195 12499 8198
rect 12801 8195 12867 8198
rect 46565 8258 46631 8261
rect 48880 8258 49000 8288
rect 46565 8256 49000 8258
rect 46565 8200 46570 8256
rect 46626 8200 49000 8256
rect 46565 8198 49000 8200
rect 46565 8195 46631 8198
rect 1946 8192 2262 8193
rect 1946 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2262 8192
rect 1946 8127 2262 8128
rect 7946 8192 8262 8193
rect 7946 8128 7952 8192
rect 8016 8128 8032 8192
rect 8096 8128 8112 8192
rect 8176 8128 8192 8192
rect 8256 8128 8262 8192
rect 7946 8127 8262 8128
rect 13946 8192 14262 8193
rect 13946 8128 13952 8192
rect 14016 8128 14032 8192
rect 14096 8128 14112 8192
rect 14176 8128 14192 8192
rect 14256 8128 14262 8192
rect 13946 8127 14262 8128
rect 19946 8192 20262 8193
rect 19946 8128 19952 8192
rect 20016 8128 20032 8192
rect 20096 8128 20112 8192
rect 20176 8128 20192 8192
rect 20256 8128 20262 8192
rect 19946 8127 20262 8128
rect 25946 8192 26262 8193
rect 25946 8128 25952 8192
rect 26016 8128 26032 8192
rect 26096 8128 26112 8192
rect 26176 8128 26192 8192
rect 26256 8128 26262 8192
rect 25946 8127 26262 8128
rect 31946 8192 32262 8193
rect 31946 8128 31952 8192
rect 32016 8128 32032 8192
rect 32096 8128 32112 8192
rect 32176 8128 32192 8192
rect 32256 8128 32262 8192
rect 31946 8127 32262 8128
rect 37946 8192 38262 8193
rect 37946 8128 37952 8192
rect 38016 8128 38032 8192
rect 38096 8128 38112 8192
rect 38176 8128 38192 8192
rect 38256 8128 38262 8192
rect 37946 8127 38262 8128
rect 43946 8192 44262 8193
rect 43946 8128 43952 8192
rect 44016 8128 44032 8192
rect 44096 8128 44112 8192
rect 44176 8128 44192 8192
rect 44256 8128 44262 8192
rect 48880 8168 49000 8198
rect 43946 8127 44262 8128
rect 0 7986 120 8016
rect 4613 7986 4679 7989
rect 0 7984 4679 7986
rect 0 7928 4618 7984
rect 4674 7928 4679 7984
rect 0 7926 4679 7928
rect 0 7896 120 7926
rect 4613 7923 4679 7926
rect 5349 7986 5415 7989
rect 45093 7986 45159 7989
rect 5349 7984 45159 7986
rect 5349 7928 5354 7984
rect 5410 7928 45098 7984
rect 45154 7928 45159 7984
rect 5349 7926 45159 7928
rect 5349 7923 5415 7926
rect 45093 7923 45159 7926
rect 46013 7986 46079 7989
rect 48880 7986 49000 8016
rect 46013 7984 49000 7986
rect 46013 7928 46018 7984
rect 46074 7928 49000 7984
rect 46013 7926 49000 7928
rect 46013 7923 46079 7926
rect 48880 7896 49000 7926
rect 2405 7850 2471 7853
rect 45645 7850 45711 7853
rect 2405 7848 45711 7850
rect 2405 7792 2410 7848
rect 2466 7792 45650 7848
rect 45706 7792 45711 7848
rect 2405 7790 45711 7792
rect 2405 7787 2471 7790
rect 45645 7787 45711 7790
rect 0 7714 120 7744
rect 11145 7714 11211 7717
rect 14273 7714 14339 7717
rect 0 7654 2790 7714
rect 0 7624 120 7654
rect 0 7442 120 7472
rect 1117 7442 1183 7445
rect 0 7440 1183 7442
rect 0 7384 1122 7440
rect 1178 7384 1183 7440
rect 0 7382 1183 7384
rect 2730 7442 2790 7654
rect 11145 7712 14339 7714
rect 11145 7656 11150 7712
rect 11206 7656 14278 7712
rect 14334 7656 14339 7712
rect 11145 7654 14339 7656
rect 11145 7651 11211 7654
rect 14273 7651 14339 7654
rect 15561 7714 15627 7717
rect 20621 7714 20687 7717
rect 15561 7712 20687 7714
rect 15561 7656 15566 7712
rect 15622 7656 20626 7712
rect 20682 7656 20687 7712
rect 15561 7654 20687 7656
rect 15561 7651 15627 7654
rect 20621 7651 20687 7654
rect 47301 7714 47367 7717
rect 48880 7714 49000 7744
rect 47301 7712 49000 7714
rect 47301 7656 47306 7712
rect 47362 7656 49000 7712
rect 47301 7654 49000 7656
rect 47301 7651 47367 7654
rect 3006 7648 3322 7649
rect 3006 7584 3012 7648
rect 3076 7584 3092 7648
rect 3156 7584 3172 7648
rect 3236 7584 3252 7648
rect 3316 7584 3322 7648
rect 3006 7583 3322 7584
rect 9006 7648 9322 7649
rect 9006 7584 9012 7648
rect 9076 7584 9092 7648
rect 9156 7584 9172 7648
rect 9236 7584 9252 7648
rect 9316 7584 9322 7648
rect 9006 7583 9322 7584
rect 15006 7648 15322 7649
rect 15006 7584 15012 7648
rect 15076 7584 15092 7648
rect 15156 7584 15172 7648
rect 15236 7584 15252 7648
rect 15316 7584 15322 7648
rect 15006 7583 15322 7584
rect 21006 7648 21322 7649
rect 21006 7584 21012 7648
rect 21076 7584 21092 7648
rect 21156 7584 21172 7648
rect 21236 7584 21252 7648
rect 21316 7584 21322 7648
rect 21006 7583 21322 7584
rect 27006 7648 27322 7649
rect 27006 7584 27012 7648
rect 27076 7584 27092 7648
rect 27156 7584 27172 7648
rect 27236 7584 27252 7648
rect 27316 7584 27322 7648
rect 27006 7583 27322 7584
rect 33006 7648 33322 7649
rect 33006 7584 33012 7648
rect 33076 7584 33092 7648
rect 33156 7584 33172 7648
rect 33236 7584 33252 7648
rect 33316 7584 33322 7648
rect 33006 7583 33322 7584
rect 39006 7648 39322 7649
rect 39006 7584 39012 7648
rect 39076 7584 39092 7648
rect 39156 7584 39172 7648
rect 39236 7584 39252 7648
rect 39316 7584 39322 7648
rect 39006 7583 39322 7584
rect 45006 7648 45322 7649
rect 45006 7584 45012 7648
rect 45076 7584 45092 7648
rect 45156 7584 45172 7648
rect 45236 7584 45252 7648
rect 45316 7584 45322 7648
rect 48880 7624 49000 7654
rect 45006 7583 45322 7584
rect 20713 7578 20779 7581
rect 15518 7576 20779 7578
rect 15518 7520 20718 7576
rect 20774 7520 20779 7576
rect 15518 7518 20779 7520
rect 2730 7382 12450 7442
rect 0 7352 120 7382
rect 1117 7379 1183 7382
rect 5993 7306 6059 7309
rect 1718 7304 6059 7306
rect 1718 7248 5998 7304
rect 6054 7248 6059 7304
rect 1718 7246 6059 7248
rect 12390 7306 12450 7382
rect 14774 7380 14780 7444
rect 14844 7442 14850 7444
rect 15518 7442 15578 7518
rect 20713 7515 20779 7518
rect 14844 7382 15578 7442
rect 16573 7442 16639 7445
rect 37825 7442 37891 7445
rect 16573 7440 37891 7442
rect 16573 7384 16578 7440
rect 16634 7384 37830 7440
rect 37886 7384 37891 7440
rect 16573 7382 37891 7384
rect 14844 7380 14850 7382
rect 16573 7379 16639 7382
rect 37825 7379 37891 7382
rect 46933 7442 46999 7445
rect 48880 7442 49000 7472
rect 46933 7440 49000 7442
rect 46933 7384 46938 7440
rect 46994 7384 49000 7440
rect 46933 7382 49000 7384
rect 46933 7379 46999 7382
rect 48880 7352 49000 7382
rect 28073 7306 28139 7309
rect 12390 7246 20546 7306
rect 0 7170 120 7200
rect 1718 7170 1778 7246
rect 5993 7243 6059 7246
rect 0 7110 1778 7170
rect 0 7080 120 7110
rect 1946 7104 2262 7105
rect 1946 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2262 7104
rect 1946 7039 2262 7040
rect 7946 7104 8262 7105
rect 7946 7040 7952 7104
rect 8016 7040 8032 7104
rect 8096 7040 8112 7104
rect 8176 7040 8192 7104
rect 8256 7040 8262 7104
rect 7946 7039 8262 7040
rect 13946 7104 14262 7105
rect 13946 7040 13952 7104
rect 14016 7040 14032 7104
rect 14096 7040 14112 7104
rect 14176 7040 14192 7104
rect 14256 7040 14262 7104
rect 13946 7039 14262 7040
rect 19946 7104 20262 7105
rect 19946 7040 19952 7104
rect 20016 7040 20032 7104
rect 20096 7040 20112 7104
rect 20176 7040 20192 7104
rect 20256 7040 20262 7104
rect 19946 7039 20262 7040
rect 20486 7034 20546 7246
rect 22050 7304 28139 7306
rect 22050 7248 28078 7304
rect 28134 7248 28139 7304
rect 22050 7246 28139 7248
rect 20621 7170 20687 7173
rect 22050 7170 22110 7246
rect 28073 7243 28139 7246
rect 20621 7168 22110 7170
rect 20621 7112 20626 7168
rect 20682 7112 22110 7168
rect 20621 7110 22110 7112
rect 47393 7170 47459 7173
rect 48880 7170 49000 7200
rect 47393 7168 49000 7170
rect 47393 7112 47398 7168
rect 47454 7112 49000 7168
rect 47393 7110 49000 7112
rect 20621 7107 20687 7110
rect 47393 7107 47459 7110
rect 25946 7104 26262 7105
rect 25946 7040 25952 7104
rect 26016 7040 26032 7104
rect 26096 7040 26112 7104
rect 26176 7040 26192 7104
rect 26256 7040 26262 7104
rect 25946 7039 26262 7040
rect 31946 7104 32262 7105
rect 31946 7040 31952 7104
rect 32016 7040 32032 7104
rect 32096 7040 32112 7104
rect 32176 7040 32192 7104
rect 32256 7040 32262 7104
rect 31946 7039 32262 7040
rect 37946 7104 38262 7105
rect 37946 7040 37952 7104
rect 38016 7040 38032 7104
rect 38096 7040 38112 7104
rect 38176 7040 38192 7104
rect 38256 7040 38262 7104
rect 37946 7039 38262 7040
rect 43946 7104 44262 7105
rect 43946 7040 43952 7104
rect 44016 7040 44032 7104
rect 44096 7040 44112 7104
rect 44176 7040 44192 7104
rect 44256 7040 44262 7104
rect 48880 7080 49000 7110
rect 43946 7039 44262 7040
rect 22737 7034 22803 7037
rect 20486 7032 22803 7034
rect 20486 6976 22742 7032
rect 22798 6976 22803 7032
rect 20486 6974 22803 6976
rect 22737 6971 22803 6974
rect 0 6898 120 6928
rect 13537 6898 13603 6901
rect 0 6896 13603 6898
rect 0 6840 13542 6896
rect 13598 6840 13603 6896
rect 0 6838 13603 6840
rect 0 6808 120 6838
rect 13537 6835 13603 6838
rect 46657 6898 46723 6901
rect 48880 6898 49000 6928
rect 46657 6896 49000 6898
rect 46657 6840 46662 6896
rect 46718 6840 49000 6896
rect 46657 6838 49000 6840
rect 46657 6835 46723 6838
rect 48880 6808 49000 6838
rect 9857 6762 9923 6765
rect 35341 6762 35407 6765
rect 9857 6760 35407 6762
rect 9857 6704 9862 6760
rect 9918 6704 35346 6760
rect 35402 6704 35407 6760
rect 9857 6702 35407 6704
rect 9857 6699 9923 6702
rect 35341 6699 35407 6702
rect 0 6626 120 6656
rect 2773 6626 2839 6629
rect 0 6624 2839 6626
rect 0 6568 2778 6624
rect 2834 6568 2839 6624
rect 0 6566 2839 6568
rect 0 6536 120 6566
rect 2773 6563 2839 6566
rect 46933 6626 46999 6629
rect 48880 6626 49000 6656
rect 46933 6624 49000 6626
rect 46933 6568 46938 6624
rect 46994 6568 49000 6624
rect 46933 6566 49000 6568
rect 46933 6563 46999 6566
rect 3006 6560 3322 6561
rect 3006 6496 3012 6560
rect 3076 6496 3092 6560
rect 3156 6496 3172 6560
rect 3236 6496 3252 6560
rect 3316 6496 3322 6560
rect 3006 6495 3322 6496
rect 9006 6560 9322 6561
rect 9006 6496 9012 6560
rect 9076 6496 9092 6560
rect 9156 6496 9172 6560
rect 9236 6496 9252 6560
rect 9316 6496 9322 6560
rect 9006 6495 9322 6496
rect 15006 6560 15322 6561
rect 15006 6496 15012 6560
rect 15076 6496 15092 6560
rect 15156 6496 15172 6560
rect 15236 6496 15252 6560
rect 15316 6496 15322 6560
rect 15006 6495 15322 6496
rect 21006 6560 21322 6561
rect 21006 6496 21012 6560
rect 21076 6496 21092 6560
rect 21156 6496 21172 6560
rect 21236 6496 21252 6560
rect 21316 6496 21322 6560
rect 21006 6495 21322 6496
rect 27006 6560 27322 6561
rect 27006 6496 27012 6560
rect 27076 6496 27092 6560
rect 27156 6496 27172 6560
rect 27236 6496 27252 6560
rect 27316 6496 27322 6560
rect 27006 6495 27322 6496
rect 33006 6560 33322 6561
rect 33006 6496 33012 6560
rect 33076 6496 33092 6560
rect 33156 6496 33172 6560
rect 33236 6496 33252 6560
rect 33316 6496 33322 6560
rect 33006 6495 33322 6496
rect 39006 6560 39322 6561
rect 39006 6496 39012 6560
rect 39076 6496 39092 6560
rect 39156 6496 39172 6560
rect 39236 6496 39252 6560
rect 39316 6496 39322 6560
rect 39006 6495 39322 6496
rect 45006 6560 45322 6561
rect 45006 6496 45012 6560
rect 45076 6496 45092 6560
rect 45156 6496 45172 6560
rect 45236 6496 45252 6560
rect 45316 6496 45322 6560
rect 48880 6536 49000 6566
rect 45006 6495 45322 6496
rect 20529 6490 20595 6493
rect 15518 6488 20595 6490
rect 15518 6432 20534 6488
rect 20590 6432 20595 6488
rect 15518 6430 20595 6432
rect 0 6354 120 6384
rect 11053 6354 11119 6357
rect 15518 6354 15578 6430
rect 20529 6427 20595 6430
rect 0 6352 11119 6354
rect 0 6296 11058 6352
rect 11114 6296 11119 6352
rect 0 6294 11119 6296
rect 0 6264 120 6294
rect 11053 6291 11119 6294
rect 13494 6294 15578 6354
rect 18229 6354 18295 6357
rect 22185 6354 22251 6357
rect 18229 6352 22251 6354
rect 18229 6296 18234 6352
rect 18290 6296 22190 6352
rect 22246 6296 22251 6352
rect 18229 6294 22251 6296
rect 5625 6218 5691 6221
rect 1718 6216 5691 6218
rect 1718 6160 5630 6216
rect 5686 6160 5691 6216
rect 1718 6158 5691 6160
rect 0 6082 120 6112
rect 1718 6082 1778 6158
rect 5625 6155 5691 6158
rect 9806 6156 9812 6220
rect 9876 6218 9882 6220
rect 13494 6218 13554 6294
rect 18229 6291 18295 6294
rect 22185 6291 22251 6294
rect 46289 6354 46355 6357
rect 48880 6354 49000 6384
rect 46289 6352 49000 6354
rect 46289 6296 46294 6352
rect 46350 6296 49000 6352
rect 46289 6294 49000 6296
rect 46289 6291 46355 6294
rect 48880 6264 49000 6294
rect 36169 6218 36235 6221
rect 9876 6158 13554 6218
rect 13678 6216 36235 6218
rect 13678 6160 36174 6216
rect 36230 6160 36235 6216
rect 13678 6158 36235 6160
rect 9876 6156 9882 6158
rect 0 6022 1778 6082
rect 9489 6082 9555 6085
rect 13678 6082 13738 6158
rect 36169 6155 36235 6158
rect 9489 6080 13738 6082
rect 9489 6024 9494 6080
rect 9550 6024 13738 6080
rect 9489 6022 13738 6024
rect 47393 6082 47459 6085
rect 48880 6082 49000 6112
rect 47393 6080 49000 6082
rect 47393 6024 47398 6080
rect 47454 6024 49000 6080
rect 47393 6022 49000 6024
rect 0 5992 120 6022
rect 9489 6019 9555 6022
rect 47393 6019 47459 6022
rect 1946 6016 2262 6017
rect 1946 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2262 6016
rect 1946 5951 2262 5952
rect 7946 6016 8262 6017
rect 7946 5952 7952 6016
rect 8016 5952 8032 6016
rect 8096 5952 8112 6016
rect 8176 5952 8192 6016
rect 8256 5952 8262 6016
rect 7946 5951 8262 5952
rect 13946 6016 14262 6017
rect 13946 5952 13952 6016
rect 14016 5952 14032 6016
rect 14096 5952 14112 6016
rect 14176 5952 14192 6016
rect 14256 5952 14262 6016
rect 13946 5951 14262 5952
rect 19946 6016 20262 6017
rect 19946 5952 19952 6016
rect 20016 5952 20032 6016
rect 20096 5952 20112 6016
rect 20176 5952 20192 6016
rect 20256 5952 20262 6016
rect 19946 5951 20262 5952
rect 25946 6016 26262 6017
rect 25946 5952 25952 6016
rect 26016 5952 26032 6016
rect 26096 5952 26112 6016
rect 26176 5952 26192 6016
rect 26256 5952 26262 6016
rect 25946 5951 26262 5952
rect 31946 6016 32262 6017
rect 31946 5952 31952 6016
rect 32016 5952 32032 6016
rect 32096 5952 32112 6016
rect 32176 5952 32192 6016
rect 32256 5952 32262 6016
rect 31946 5951 32262 5952
rect 37946 6016 38262 6017
rect 37946 5952 37952 6016
rect 38016 5952 38032 6016
rect 38096 5952 38112 6016
rect 38176 5952 38192 6016
rect 38256 5952 38262 6016
rect 37946 5951 38262 5952
rect 43946 6016 44262 6017
rect 43946 5952 43952 6016
rect 44016 5952 44032 6016
rect 44096 5952 44112 6016
rect 44176 5952 44192 6016
rect 44256 5952 44262 6016
rect 48880 5992 49000 6022
rect 43946 5951 44262 5952
rect 0 5810 120 5840
rect 19793 5810 19859 5813
rect 0 5808 19859 5810
rect 0 5752 19798 5808
rect 19854 5752 19859 5808
rect 0 5750 19859 5752
rect 0 5720 120 5750
rect 19793 5747 19859 5750
rect 46565 5810 46631 5813
rect 48880 5810 49000 5840
rect 46565 5808 49000 5810
rect 46565 5752 46570 5808
rect 46626 5752 49000 5808
rect 46565 5750 49000 5752
rect 46565 5747 46631 5750
rect 48880 5720 49000 5750
rect 9806 5674 9812 5676
rect 8710 5614 9812 5674
rect 0 5538 120 5568
rect 0 5478 2882 5538
rect 0 5448 120 5478
rect 0 5266 120 5296
rect 2681 5266 2747 5269
rect 0 5264 2747 5266
rect 0 5208 2686 5264
rect 2742 5208 2747 5264
rect 0 5206 2747 5208
rect 2822 5266 2882 5478
rect 3006 5472 3322 5473
rect 3006 5408 3012 5472
rect 3076 5408 3092 5472
rect 3156 5408 3172 5472
rect 3236 5408 3252 5472
rect 3316 5408 3322 5472
rect 3006 5407 3322 5408
rect 8710 5402 8770 5614
rect 9806 5612 9812 5614
rect 9876 5612 9882 5676
rect 14917 5674 14983 5677
rect 46105 5674 46171 5677
rect 14917 5672 46171 5674
rect 14917 5616 14922 5672
rect 14978 5616 46110 5672
rect 46166 5616 46171 5672
rect 14917 5614 46171 5616
rect 14917 5611 14983 5614
rect 46105 5611 46171 5614
rect 14774 5538 14780 5540
rect 9446 5478 14780 5538
rect 9006 5472 9322 5473
rect 9006 5408 9012 5472
rect 9076 5408 9092 5472
rect 9156 5408 9172 5472
rect 9236 5408 9252 5472
rect 9316 5408 9322 5472
rect 9006 5407 9322 5408
rect 3558 5342 8770 5402
rect 3141 5266 3207 5269
rect 3558 5266 3618 5342
rect 2822 5206 3066 5266
rect 0 5176 120 5206
rect 2681 5203 2747 5206
rect 2865 5130 2931 5133
rect 1718 5128 2931 5130
rect 1718 5072 2870 5128
rect 2926 5072 2931 5128
rect 1718 5070 2931 5072
rect 3006 5130 3066 5206
rect 3141 5264 3618 5266
rect 3141 5208 3146 5264
rect 3202 5208 3618 5264
rect 3141 5206 3618 5208
rect 7465 5266 7531 5269
rect 9446 5266 9506 5478
rect 14774 5476 14780 5478
rect 14844 5476 14850 5540
rect 47025 5538 47091 5541
rect 48880 5538 49000 5568
rect 47025 5536 49000 5538
rect 47025 5480 47030 5536
rect 47086 5480 49000 5536
rect 47025 5478 49000 5480
rect 47025 5475 47091 5478
rect 15006 5472 15322 5473
rect 15006 5408 15012 5472
rect 15076 5408 15092 5472
rect 15156 5408 15172 5472
rect 15236 5408 15252 5472
rect 15316 5408 15322 5472
rect 15006 5407 15322 5408
rect 21006 5472 21322 5473
rect 21006 5408 21012 5472
rect 21076 5408 21092 5472
rect 21156 5408 21172 5472
rect 21236 5408 21252 5472
rect 21316 5408 21322 5472
rect 21006 5407 21322 5408
rect 27006 5472 27322 5473
rect 27006 5408 27012 5472
rect 27076 5408 27092 5472
rect 27156 5408 27172 5472
rect 27236 5408 27252 5472
rect 27316 5408 27322 5472
rect 27006 5407 27322 5408
rect 33006 5472 33322 5473
rect 33006 5408 33012 5472
rect 33076 5408 33092 5472
rect 33156 5408 33172 5472
rect 33236 5408 33252 5472
rect 33316 5408 33322 5472
rect 33006 5407 33322 5408
rect 39006 5472 39322 5473
rect 39006 5408 39012 5472
rect 39076 5408 39092 5472
rect 39156 5408 39172 5472
rect 39236 5408 39252 5472
rect 39316 5408 39322 5472
rect 39006 5407 39322 5408
rect 45006 5472 45322 5473
rect 45006 5408 45012 5472
rect 45076 5408 45092 5472
rect 45156 5408 45172 5472
rect 45236 5408 45252 5472
rect 45316 5408 45322 5472
rect 48880 5448 49000 5478
rect 45006 5407 45322 5408
rect 9673 5402 9739 5405
rect 14825 5402 14891 5405
rect 9673 5400 14891 5402
rect 9673 5344 9678 5400
rect 9734 5344 14830 5400
rect 14886 5344 14891 5400
rect 9673 5342 14891 5344
rect 9673 5339 9739 5342
rect 14825 5339 14891 5342
rect 7465 5264 9506 5266
rect 7465 5208 7470 5264
rect 7526 5208 9506 5264
rect 7465 5206 9506 5208
rect 9581 5266 9647 5269
rect 32765 5266 32831 5269
rect 9581 5264 32831 5266
rect 9581 5208 9586 5264
rect 9642 5208 32770 5264
rect 32826 5208 32831 5264
rect 9581 5206 32831 5208
rect 3141 5203 3207 5206
rect 7465 5203 7531 5206
rect 9581 5203 9647 5206
rect 32765 5203 32831 5206
rect 47301 5266 47367 5269
rect 48880 5266 49000 5296
rect 47301 5264 49000 5266
rect 47301 5208 47306 5264
rect 47362 5208 49000 5264
rect 47301 5206 49000 5208
rect 47301 5203 47367 5206
rect 48880 5176 49000 5206
rect 14825 5130 14891 5133
rect 37549 5130 37615 5133
rect 3006 5070 14658 5130
rect 0 4994 120 5024
rect 1718 4994 1778 5070
rect 2865 5067 2931 5070
rect 0 4934 1778 4994
rect 2681 4994 2747 4997
rect 14598 4994 14658 5070
rect 14825 5128 37615 5130
rect 14825 5072 14830 5128
rect 14886 5072 37554 5128
rect 37610 5072 37615 5128
rect 14825 5070 37615 5072
rect 14825 5067 14891 5070
rect 37549 5067 37615 5070
rect 17401 4994 17467 4997
rect 2681 4992 7666 4994
rect 2681 4936 2686 4992
rect 2742 4936 7666 4992
rect 2681 4934 7666 4936
rect 14598 4992 17467 4994
rect 14598 4936 17406 4992
rect 17462 4936 17467 4992
rect 14598 4934 17467 4936
rect 0 4904 120 4934
rect 2681 4931 2747 4934
rect 1946 4928 2262 4929
rect 1946 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2262 4928
rect 1946 4863 2262 4864
rect 0 4722 120 4752
rect 7465 4722 7531 4725
rect 0 4720 7531 4722
rect 0 4664 7470 4720
rect 7526 4664 7531 4720
rect 0 4662 7531 4664
rect 7606 4722 7666 4934
rect 17401 4931 17467 4934
rect 46933 4994 46999 4997
rect 48880 4994 49000 5024
rect 46933 4992 49000 4994
rect 46933 4936 46938 4992
rect 46994 4936 49000 4992
rect 46933 4934 49000 4936
rect 46933 4931 46999 4934
rect 7946 4928 8262 4929
rect 7946 4864 7952 4928
rect 8016 4864 8032 4928
rect 8096 4864 8112 4928
rect 8176 4864 8192 4928
rect 8256 4864 8262 4928
rect 7946 4863 8262 4864
rect 13946 4928 14262 4929
rect 13946 4864 13952 4928
rect 14016 4864 14032 4928
rect 14096 4864 14112 4928
rect 14176 4864 14192 4928
rect 14256 4864 14262 4928
rect 13946 4863 14262 4864
rect 19946 4928 20262 4929
rect 19946 4864 19952 4928
rect 20016 4864 20032 4928
rect 20096 4864 20112 4928
rect 20176 4864 20192 4928
rect 20256 4864 20262 4928
rect 19946 4863 20262 4864
rect 25946 4928 26262 4929
rect 25946 4864 25952 4928
rect 26016 4864 26032 4928
rect 26096 4864 26112 4928
rect 26176 4864 26192 4928
rect 26256 4864 26262 4928
rect 25946 4863 26262 4864
rect 31946 4928 32262 4929
rect 31946 4864 31952 4928
rect 32016 4864 32032 4928
rect 32096 4864 32112 4928
rect 32176 4864 32192 4928
rect 32256 4864 32262 4928
rect 31946 4863 32262 4864
rect 37946 4928 38262 4929
rect 37946 4864 37952 4928
rect 38016 4864 38032 4928
rect 38096 4864 38112 4928
rect 38176 4864 38192 4928
rect 38256 4864 38262 4928
rect 37946 4863 38262 4864
rect 43946 4928 44262 4929
rect 43946 4864 43952 4928
rect 44016 4864 44032 4928
rect 44096 4864 44112 4928
rect 44176 4864 44192 4928
rect 44256 4864 44262 4928
rect 48880 4904 49000 4934
rect 43946 4863 44262 4864
rect 17861 4722 17927 4725
rect 7606 4720 17927 4722
rect 7606 4664 17866 4720
rect 17922 4664 17927 4720
rect 7606 4662 17927 4664
rect 0 4632 120 4662
rect 7465 4659 7531 4662
rect 17861 4659 17927 4662
rect 47393 4722 47459 4725
rect 48880 4722 49000 4752
rect 47393 4720 49000 4722
rect 47393 4664 47398 4720
rect 47454 4664 49000 4720
rect 47393 4662 49000 4664
rect 47393 4659 47459 4662
rect 48880 4632 49000 4662
rect 13629 4586 13695 4589
rect 2730 4584 13695 4586
rect 2730 4528 13634 4584
rect 13690 4528 13695 4584
rect 2730 4526 13695 4528
rect 0 4450 120 4480
rect 2730 4450 2790 4526
rect 13629 4523 13695 4526
rect 0 4390 2790 4450
rect 47025 4450 47091 4453
rect 48880 4450 49000 4480
rect 47025 4448 49000 4450
rect 47025 4392 47030 4448
rect 47086 4392 49000 4448
rect 47025 4390 49000 4392
rect 0 4360 120 4390
rect 47025 4387 47091 4390
rect 3006 4384 3322 4385
rect 3006 4320 3012 4384
rect 3076 4320 3092 4384
rect 3156 4320 3172 4384
rect 3236 4320 3252 4384
rect 3316 4320 3322 4384
rect 3006 4319 3322 4320
rect 9006 4384 9322 4385
rect 9006 4320 9012 4384
rect 9076 4320 9092 4384
rect 9156 4320 9172 4384
rect 9236 4320 9252 4384
rect 9316 4320 9322 4384
rect 9006 4319 9322 4320
rect 15006 4384 15322 4385
rect 15006 4320 15012 4384
rect 15076 4320 15092 4384
rect 15156 4320 15172 4384
rect 15236 4320 15252 4384
rect 15316 4320 15322 4384
rect 15006 4319 15322 4320
rect 21006 4384 21322 4385
rect 21006 4320 21012 4384
rect 21076 4320 21092 4384
rect 21156 4320 21172 4384
rect 21236 4320 21252 4384
rect 21316 4320 21322 4384
rect 21006 4319 21322 4320
rect 27006 4384 27322 4385
rect 27006 4320 27012 4384
rect 27076 4320 27092 4384
rect 27156 4320 27172 4384
rect 27236 4320 27252 4384
rect 27316 4320 27322 4384
rect 27006 4319 27322 4320
rect 33006 4384 33322 4385
rect 33006 4320 33012 4384
rect 33076 4320 33092 4384
rect 33156 4320 33172 4384
rect 33236 4320 33252 4384
rect 33316 4320 33322 4384
rect 33006 4319 33322 4320
rect 39006 4384 39322 4385
rect 39006 4320 39012 4384
rect 39076 4320 39092 4384
rect 39156 4320 39172 4384
rect 39236 4320 39252 4384
rect 39316 4320 39322 4384
rect 39006 4319 39322 4320
rect 45006 4384 45322 4385
rect 45006 4320 45012 4384
rect 45076 4320 45092 4384
rect 45156 4320 45172 4384
rect 45236 4320 45252 4384
rect 45316 4320 45322 4384
rect 48880 4360 49000 4390
rect 45006 4319 45322 4320
rect 0 4178 120 4208
rect 24669 4178 24735 4181
rect 0 4176 24735 4178
rect 0 4120 24674 4176
rect 24730 4120 24735 4176
rect 0 4118 24735 4120
rect 0 4088 120 4118
rect 24669 4115 24735 4118
rect 47301 4178 47367 4181
rect 48880 4178 49000 4208
rect 47301 4176 49000 4178
rect 47301 4120 47306 4176
rect 47362 4120 49000 4176
rect 47301 4118 49000 4120
rect 47301 4115 47367 4118
rect 48880 4088 49000 4118
rect 17953 4042 18019 4045
rect 24761 4042 24827 4045
rect 1718 4040 18019 4042
rect 1718 3984 17958 4040
rect 18014 3984 18019 4040
rect 1718 3982 18019 3984
rect 0 3906 120 3936
rect 1718 3906 1778 3982
rect 17953 3979 18019 3982
rect 18094 4040 24827 4042
rect 18094 3984 24766 4040
rect 24822 3984 24827 4040
rect 18094 3982 24827 3984
rect 0 3846 1778 3906
rect 14825 3906 14891 3909
rect 18094 3906 18154 3982
rect 24761 3979 24827 3982
rect 14825 3904 18154 3906
rect 14825 3848 14830 3904
rect 14886 3848 18154 3904
rect 14825 3846 18154 3848
rect 46933 3906 46999 3909
rect 48880 3906 49000 3936
rect 46933 3904 49000 3906
rect 46933 3848 46938 3904
rect 46994 3848 49000 3904
rect 46933 3846 49000 3848
rect 0 3816 120 3846
rect 14825 3843 14891 3846
rect 46933 3843 46999 3846
rect 1946 3840 2262 3841
rect 1946 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2262 3840
rect 1946 3775 2262 3776
rect 7946 3840 8262 3841
rect 7946 3776 7952 3840
rect 8016 3776 8032 3840
rect 8096 3776 8112 3840
rect 8176 3776 8192 3840
rect 8256 3776 8262 3840
rect 7946 3775 8262 3776
rect 13946 3840 14262 3841
rect 13946 3776 13952 3840
rect 14016 3776 14032 3840
rect 14096 3776 14112 3840
rect 14176 3776 14192 3840
rect 14256 3776 14262 3840
rect 13946 3775 14262 3776
rect 19946 3840 20262 3841
rect 19946 3776 19952 3840
rect 20016 3776 20032 3840
rect 20096 3776 20112 3840
rect 20176 3776 20192 3840
rect 20256 3776 20262 3840
rect 19946 3775 20262 3776
rect 25946 3840 26262 3841
rect 25946 3776 25952 3840
rect 26016 3776 26032 3840
rect 26096 3776 26112 3840
rect 26176 3776 26192 3840
rect 26256 3776 26262 3840
rect 25946 3775 26262 3776
rect 31946 3840 32262 3841
rect 31946 3776 31952 3840
rect 32016 3776 32032 3840
rect 32096 3776 32112 3840
rect 32176 3776 32192 3840
rect 32256 3776 32262 3840
rect 31946 3775 32262 3776
rect 37946 3840 38262 3841
rect 37946 3776 37952 3840
rect 38016 3776 38032 3840
rect 38096 3776 38112 3840
rect 38176 3776 38192 3840
rect 38256 3776 38262 3840
rect 37946 3775 38262 3776
rect 43946 3840 44262 3841
rect 43946 3776 43952 3840
rect 44016 3776 44032 3840
rect 44096 3776 44112 3840
rect 44176 3776 44192 3840
rect 44256 3776 44262 3840
rect 48880 3816 49000 3846
rect 43946 3775 44262 3776
rect 0 3634 120 3664
rect 24853 3634 24919 3637
rect 0 3632 24919 3634
rect 0 3576 24858 3632
rect 24914 3576 24919 3632
rect 0 3574 24919 3576
rect 0 3544 120 3574
rect 24853 3571 24919 3574
rect 28993 3634 29059 3637
rect 41597 3634 41663 3637
rect 28993 3632 41663 3634
rect 28993 3576 28998 3632
rect 29054 3576 41602 3632
rect 41658 3576 41663 3632
rect 28993 3574 41663 3576
rect 28993 3571 29059 3574
rect 41597 3571 41663 3574
rect 47393 3634 47459 3637
rect 48880 3634 49000 3664
rect 47393 3632 49000 3634
rect 47393 3576 47398 3632
rect 47454 3576 49000 3632
rect 47393 3574 49000 3576
rect 47393 3571 47459 3574
rect 48880 3544 49000 3574
rect 20713 3498 20779 3501
rect 2730 3496 20779 3498
rect 2730 3440 20718 3496
rect 20774 3440 20779 3496
rect 2730 3438 20779 3440
rect 0 3362 120 3392
rect 2730 3362 2790 3438
rect 20713 3435 20779 3438
rect 25865 3498 25931 3501
rect 44173 3498 44239 3501
rect 25865 3496 44239 3498
rect 25865 3440 25870 3496
rect 25926 3440 44178 3496
rect 44234 3440 44239 3496
rect 25865 3438 44239 3440
rect 25865 3435 25931 3438
rect 44173 3435 44239 3438
rect 0 3302 2790 3362
rect 47025 3362 47091 3365
rect 48880 3362 49000 3392
rect 47025 3360 49000 3362
rect 47025 3304 47030 3360
rect 47086 3304 49000 3360
rect 47025 3302 49000 3304
rect 0 3272 120 3302
rect 47025 3299 47091 3302
rect 3006 3296 3322 3297
rect 3006 3232 3012 3296
rect 3076 3232 3092 3296
rect 3156 3232 3172 3296
rect 3236 3232 3252 3296
rect 3316 3232 3322 3296
rect 3006 3231 3322 3232
rect 9006 3296 9322 3297
rect 9006 3232 9012 3296
rect 9076 3232 9092 3296
rect 9156 3232 9172 3296
rect 9236 3232 9252 3296
rect 9316 3232 9322 3296
rect 9006 3231 9322 3232
rect 15006 3296 15322 3297
rect 15006 3232 15012 3296
rect 15076 3232 15092 3296
rect 15156 3232 15172 3296
rect 15236 3232 15252 3296
rect 15316 3232 15322 3296
rect 15006 3231 15322 3232
rect 21006 3296 21322 3297
rect 21006 3232 21012 3296
rect 21076 3232 21092 3296
rect 21156 3232 21172 3296
rect 21236 3232 21252 3296
rect 21316 3232 21322 3296
rect 21006 3231 21322 3232
rect 27006 3296 27322 3297
rect 27006 3232 27012 3296
rect 27076 3232 27092 3296
rect 27156 3232 27172 3296
rect 27236 3232 27252 3296
rect 27316 3232 27322 3296
rect 27006 3231 27322 3232
rect 33006 3296 33322 3297
rect 33006 3232 33012 3296
rect 33076 3232 33092 3296
rect 33156 3232 33172 3296
rect 33236 3232 33252 3296
rect 33316 3232 33322 3296
rect 33006 3231 33322 3232
rect 39006 3296 39322 3297
rect 39006 3232 39012 3296
rect 39076 3232 39092 3296
rect 39156 3232 39172 3296
rect 39236 3232 39252 3296
rect 39316 3232 39322 3296
rect 39006 3231 39322 3232
rect 45006 3296 45322 3297
rect 45006 3232 45012 3296
rect 45076 3232 45092 3296
rect 45156 3232 45172 3296
rect 45236 3232 45252 3296
rect 45316 3232 45322 3296
rect 48880 3272 49000 3302
rect 45006 3231 45322 3232
rect 9397 3226 9463 3229
rect 14825 3226 14891 3229
rect 9397 3224 14891 3226
rect 9397 3168 9402 3224
rect 9458 3168 14830 3224
rect 14886 3168 14891 3224
rect 9397 3166 14891 3168
rect 9397 3163 9463 3166
rect 14825 3163 14891 3166
rect 0 3090 120 3120
rect 17217 3090 17283 3093
rect 0 3088 17283 3090
rect 0 3032 17222 3088
rect 17278 3032 17283 3088
rect 0 3030 17283 3032
rect 0 3000 120 3030
rect 17217 3027 17283 3030
rect 28533 3090 28599 3093
rect 46749 3090 46815 3093
rect 28533 3088 46815 3090
rect 28533 3032 28538 3088
rect 28594 3032 46754 3088
rect 46810 3032 46815 3088
rect 28533 3030 46815 3032
rect 28533 3027 28599 3030
rect 46749 3027 46815 3030
rect 47301 3090 47367 3093
rect 48880 3090 49000 3120
rect 47301 3088 49000 3090
rect 47301 3032 47306 3088
rect 47362 3032 49000 3088
rect 47301 3030 49000 3032
rect 47301 3027 47367 3030
rect 48880 3000 49000 3030
rect 9397 2954 9463 2957
rect 1718 2952 9463 2954
rect 1718 2896 9402 2952
rect 9458 2896 9463 2952
rect 1718 2894 9463 2896
rect 0 2818 120 2848
rect 1718 2818 1778 2894
rect 9397 2891 9463 2894
rect 11053 2954 11119 2957
rect 41413 2954 41479 2957
rect 11053 2952 41479 2954
rect 11053 2896 11058 2952
rect 11114 2896 41418 2952
rect 41474 2896 41479 2952
rect 11053 2894 41479 2896
rect 11053 2891 11119 2894
rect 41413 2891 41479 2894
rect 0 2758 1778 2818
rect 46933 2818 46999 2821
rect 48880 2818 49000 2848
rect 46933 2816 49000 2818
rect 46933 2760 46938 2816
rect 46994 2760 49000 2816
rect 46933 2758 49000 2760
rect 0 2728 120 2758
rect 46933 2755 46999 2758
rect 1946 2752 2262 2753
rect 1946 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2262 2752
rect 1946 2687 2262 2688
rect 7946 2752 8262 2753
rect 7946 2688 7952 2752
rect 8016 2688 8032 2752
rect 8096 2688 8112 2752
rect 8176 2688 8192 2752
rect 8256 2688 8262 2752
rect 7946 2687 8262 2688
rect 13946 2752 14262 2753
rect 13946 2688 13952 2752
rect 14016 2688 14032 2752
rect 14096 2688 14112 2752
rect 14176 2688 14192 2752
rect 14256 2688 14262 2752
rect 13946 2687 14262 2688
rect 19946 2752 20262 2753
rect 19946 2688 19952 2752
rect 20016 2688 20032 2752
rect 20096 2688 20112 2752
rect 20176 2688 20192 2752
rect 20256 2688 20262 2752
rect 19946 2687 20262 2688
rect 25946 2752 26262 2753
rect 25946 2688 25952 2752
rect 26016 2688 26032 2752
rect 26096 2688 26112 2752
rect 26176 2688 26192 2752
rect 26256 2688 26262 2752
rect 25946 2687 26262 2688
rect 31946 2752 32262 2753
rect 31946 2688 31952 2752
rect 32016 2688 32032 2752
rect 32096 2688 32112 2752
rect 32176 2688 32192 2752
rect 32256 2688 32262 2752
rect 31946 2687 32262 2688
rect 37946 2752 38262 2753
rect 37946 2688 37952 2752
rect 38016 2688 38032 2752
rect 38096 2688 38112 2752
rect 38176 2688 38192 2752
rect 38256 2688 38262 2752
rect 37946 2687 38262 2688
rect 43946 2752 44262 2753
rect 43946 2688 43952 2752
rect 44016 2688 44032 2752
rect 44096 2688 44112 2752
rect 44176 2688 44192 2752
rect 44256 2688 44262 2752
rect 48880 2728 49000 2758
rect 43946 2687 44262 2688
rect 0 2546 120 2576
rect 9489 2546 9555 2549
rect 0 2544 9555 2546
rect 0 2488 9494 2544
rect 9550 2488 9555 2544
rect 0 2486 9555 2488
rect 0 2456 120 2486
rect 9489 2483 9555 2486
rect 42149 2546 42215 2549
rect 45645 2546 45711 2549
rect 42149 2544 45711 2546
rect 42149 2488 42154 2544
rect 42210 2488 45650 2544
rect 45706 2488 45711 2544
rect 42149 2486 45711 2488
rect 42149 2483 42215 2486
rect 45645 2483 45711 2486
rect 47301 2546 47367 2549
rect 48880 2546 49000 2576
rect 47301 2544 49000 2546
rect 47301 2488 47306 2544
rect 47362 2488 49000 2544
rect 47301 2486 49000 2488
rect 47301 2483 47367 2486
rect 48880 2456 49000 2486
rect 20713 2410 20779 2413
rect 2822 2408 20779 2410
rect 2822 2352 20718 2408
rect 20774 2352 20779 2408
rect 2822 2350 20779 2352
rect 0 2274 120 2304
rect 2822 2274 2882 2350
rect 20713 2347 20779 2350
rect 0 2214 2882 2274
rect 46933 2274 46999 2277
rect 48880 2274 49000 2304
rect 46933 2272 49000 2274
rect 46933 2216 46938 2272
rect 46994 2216 49000 2272
rect 46933 2214 49000 2216
rect 0 2184 120 2214
rect 46933 2211 46999 2214
rect 3006 2208 3322 2209
rect 3006 2144 3012 2208
rect 3076 2144 3092 2208
rect 3156 2144 3172 2208
rect 3236 2144 3252 2208
rect 3316 2144 3322 2208
rect 3006 2143 3322 2144
rect 9006 2208 9322 2209
rect 9006 2144 9012 2208
rect 9076 2144 9092 2208
rect 9156 2144 9172 2208
rect 9236 2144 9252 2208
rect 9316 2144 9322 2208
rect 9006 2143 9322 2144
rect 15006 2208 15322 2209
rect 15006 2144 15012 2208
rect 15076 2144 15092 2208
rect 15156 2144 15172 2208
rect 15236 2144 15252 2208
rect 15316 2144 15322 2208
rect 15006 2143 15322 2144
rect 21006 2208 21322 2209
rect 21006 2144 21012 2208
rect 21076 2144 21092 2208
rect 21156 2144 21172 2208
rect 21236 2144 21252 2208
rect 21316 2144 21322 2208
rect 21006 2143 21322 2144
rect 27006 2208 27322 2209
rect 27006 2144 27012 2208
rect 27076 2144 27092 2208
rect 27156 2144 27172 2208
rect 27236 2144 27252 2208
rect 27316 2144 27322 2208
rect 27006 2143 27322 2144
rect 33006 2208 33322 2209
rect 33006 2144 33012 2208
rect 33076 2144 33092 2208
rect 33156 2144 33172 2208
rect 33236 2144 33252 2208
rect 33316 2144 33322 2208
rect 33006 2143 33322 2144
rect 39006 2208 39322 2209
rect 39006 2144 39012 2208
rect 39076 2144 39092 2208
rect 39156 2144 39172 2208
rect 39236 2144 39252 2208
rect 39316 2144 39322 2208
rect 39006 2143 39322 2144
rect 45006 2208 45322 2209
rect 45006 2144 45012 2208
rect 45076 2144 45092 2208
rect 45156 2144 45172 2208
rect 45236 2144 45252 2208
rect 45316 2144 45322 2208
rect 48880 2184 49000 2214
rect 45006 2143 45322 2144
rect 0 2002 120 2032
rect 19701 2002 19767 2005
rect 0 2000 19767 2002
rect 0 1944 19706 2000
rect 19762 1944 19767 2000
rect 0 1942 19767 1944
rect 0 1912 120 1942
rect 19701 1939 19767 1942
rect 45829 2002 45895 2005
rect 48880 2002 49000 2032
rect 45829 2000 49000 2002
rect 45829 1944 45834 2000
rect 45890 1944 49000 2000
rect 45829 1942 49000 1944
rect 45829 1939 45895 1942
rect 48880 1912 49000 1942
rect 0 1730 120 1760
rect 9581 1730 9647 1733
rect 0 1728 9647 1730
rect 0 1672 9586 1728
rect 9642 1672 9647 1728
rect 0 1670 9647 1672
rect 0 1640 120 1670
rect 9581 1667 9647 1670
rect 46197 1730 46263 1733
rect 48880 1730 49000 1760
rect 46197 1728 49000 1730
rect 46197 1672 46202 1728
rect 46258 1672 49000 1728
rect 46197 1670 49000 1672
rect 46197 1667 46263 1670
rect 48880 1640 49000 1670
rect 0 1458 120 1488
rect 1301 1458 1367 1461
rect 0 1456 1367 1458
rect 0 1400 1306 1456
rect 1362 1400 1367 1456
rect 0 1398 1367 1400
rect 0 1368 120 1398
rect 1301 1395 1367 1398
rect 46565 1458 46631 1461
rect 48880 1458 49000 1488
rect 46565 1456 49000 1458
rect 46565 1400 46570 1456
rect 46626 1400 49000 1456
rect 46565 1398 49000 1400
rect 46565 1395 46631 1398
rect 48880 1368 49000 1398
<< via3 >>
rect 3012 8732 3076 8736
rect 3012 8676 3016 8732
rect 3016 8676 3072 8732
rect 3072 8676 3076 8732
rect 3012 8672 3076 8676
rect 3092 8732 3156 8736
rect 3092 8676 3096 8732
rect 3096 8676 3152 8732
rect 3152 8676 3156 8732
rect 3092 8672 3156 8676
rect 3172 8732 3236 8736
rect 3172 8676 3176 8732
rect 3176 8676 3232 8732
rect 3232 8676 3236 8732
rect 3172 8672 3236 8676
rect 3252 8732 3316 8736
rect 3252 8676 3256 8732
rect 3256 8676 3312 8732
rect 3312 8676 3316 8732
rect 3252 8672 3316 8676
rect 9012 8732 9076 8736
rect 9012 8676 9016 8732
rect 9016 8676 9072 8732
rect 9072 8676 9076 8732
rect 9012 8672 9076 8676
rect 9092 8732 9156 8736
rect 9092 8676 9096 8732
rect 9096 8676 9152 8732
rect 9152 8676 9156 8732
rect 9092 8672 9156 8676
rect 9172 8732 9236 8736
rect 9172 8676 9176 8732
rect 9176 8676 9232 8732
rect 9232 8676 9236 8732
rect 9172 8672 9236 8676
rect 9252 8732 9316 8736
rect 9252 8676 9256 8732
rect 9256 8676 9312 8732
rect 9312 8676 9316 8732
rect 9252 8672 9316 8676
rect 15012 8732 15076 8736
rect 15012 8676 15016 8732
rect 15016 8676 15072 8732
rect 15072 8676 15076 8732
rect 15012 8672 15076 8676
rect 15092 8732 15156 8736
rect 15092 8676 15096 8732
rect 15096 8676 15152 8732
rect 15152 8676 15156 8732
rect 15092 8672 15156 8676
rect 15172 8732 15236 8736
rect 15172 8676 15176 8732
rect 15176 8676 15232 8732
rect 15232 8676 15236 8732
rect 15172 8672 15236 8676
rect 15252 8732 15316 8736
rect 15252 8676 15256 8732
rect 15256 8676 15312 8732
rect 15312 8676 15316 8732
rect 15252 8672 15316 8676
rect 21012 8732 21076 8736
rect 21012 8676 21016 8732
rect 21016 8676 21072 8732
rect 21072 8676 21076 8732
rect 21012 8672 21076 8676
rect 21092 8732 21156 8736
rect 21092 8676 21096 8732
rect 21096 8676 21152 8732
rect 21152 8676 21156 8732
rect 21092 8672 21156 8676
rect 21172 8732 21236 8736
rect 21172 8676 21176 8732
rect 21176 8676 21232 8732
rect 21232 8676 21236 8732
rect 21172 8672 21236 8676
rect 21252 8732 21316 8736
rect 21252 8676 21256 8732
rect 21256 8676 21312 8732
rect 21312 8676 21316 8732
rect 21252 8672 21316 8676
rect 27012 8732 27076 8736
rect 27012 8676 27016 8732
rect 27016 8676 27072 8732
rect 27072 8676 27076 8732
rect 27012 8672 27076 8676
rect 27092 8732 27156 8736
rect 27092 8676 27096 8732
rect 27096 8676 27152 8732
rect 27152 8676 27156 8732
rect 27092 8672 27156 8676
rect 27172 8732 27236 8736
rect 27172 8676 27176 8732
rect 27176 8676 27232 8732
rect 27232 8676 27236 8732
rect 27172 8672 27236 8676
rect 27252 8732 27316 8736
rect 27252 8676 27256 8732
rect 27256 8676 27312 8732
rect 27312 8676 27316 8732
rect 27252 8672 27316 8676
rect 33012 8732 33076 8736
rect 33012 8676 33016 8732
rect 33016 8676 33072 8732
rect 33072 8676 33076 8732
rect 33012 8672 33076 8676
rect 33092 8732 33156 8736
rect 33092 8676 33096 8732
rect 33096 8676 33152 8732
rect 33152 8676 33156 8732
rect 33092 8672 33156 8676
rect 33172 8732 33236 8736
rect 33172 8676 33176 8732
rect 33176 8676 33232 8732
rect 33232 8676 33236 8732
rect 33172 8672 33236 8676
rect 33252 8732 33316 8736
rect 33252 8676 33256 8732
rect 33256 8676 33312 8732
rect 33312 8676 33316 8732
rect 33252 8672 33316 8676
rect 39012 8732 39076 8736
rect 39012 8676 39016 8732
rect 39016 8676 39072 8732
rect 39072 8676 39076 8732
rect 39012 8672 39076 8676
rect 39092 8732 39156 8736
rect 39092 8676 39096 8732
rect 39096 8676 39152 8732
rect 39152 8676 39156 8732
rect 39092 8672 39156 8676
rect 39172 8732 39236 8736
rect 39172 8676 39176 8732
rect 39176 8676 39232 8732
rect 39232 8676 39236 8732
rect 39172 8672 39236 8676
rect 39252 8732 39316 8736
rect 39252 8676 39256 8732
rect 39256 8676 39312 8732
rect 39312 8676 39316 8732
rect 39252 8672 39316 8676
rect 45012 8732 45076 8736
rect 45012 8676 45016 8732
rect 45016 8676 45072 8732
rect 45072 8676 45076 8732
rect 45012 8672 45076 8676
rect 45092 8732 45156 8736
rect 45092 8676 45096 8732
rect 45096 8676 45152 8732
rect 45152 8676 45156 8732
rect 45092 8672 45156 8676
rect 45172 8732 45236 8736
rect 45172 8676 45176 8732
rect 45176 8676 45232 8732
rect 45232 8676 45236 8732
rect 45172 8672 45236 8676
rect 45252 8732 45316 8736
rect 45252 8676 45256 8732
rect 45256 8676 45312 8732
rect 45312 8676 45316 8732
rect 45252 8672 45316 8676
rect 1952 8188 2016 8192
rect 1952 8132 1956 8188
rect 1956 8132 2012 8188
rect 2012 8132 2016 8188
rect 1952 8128 2016 8132
rect 2032 8188 2096 8192
rect 2032 8132 2036 8188
rect 2036 8132 2092 8188
rect 2092 8132 2096 8188
rect 2032 8128 2096 8132
rect 2112 8188 2176 8192
rect 2112 8132 2116 8188
rect 2116 8132 2172 8188
rect 2172 8132 2176 8188
rect 2112 8128 2176 8132
rect 2192 8188 2256 8192
rect 2192 8132 2196 8188
rect 2196 8132 2252 8188
rect 2252 8132 2256 8188
rect 2192 8128 2256 8132
rect 7952 8188 8016 8192
rect 7952 8132 7956 8188
rect 7956 8132 8012 8188
rect 8012 8132 8016 8188
rect 7952 8128 8016 8132
rect 8032 8188 8096 8192
rect 8032 8132 8036 8188
rect 8036 8132 8092 8188
rect 8092 8132 8096 8188
rect 8032 8128 8096 8132
rect 8112 8188 8176 8192
rect 8112 8132 8116 8188
rect 8116 8132 8172 8188
rect 8172 8132 8176 8188
rect 8112 8128 8176 8132
rect 8192 8188 8256 8192
rect 8192 8132 8196 8188
rect 8196 8132 8252 8188
rect 8252 8132 8256 8188
rect 8192 8128 8256 8132
rect 13952 8188 14016 8192
rect 13952 8132 13956 8188
rect 13956 8132 14012 8188
rect 14012 8132 14016 8188
rect 13952 8128 14016 8132
rect 14032 8188 14096 8192
rect 14032 8132 14036 8188
rect 14036 8132 14092 8188
rect 14092 8132 14096 8188
rect 14032 8128 14096 8132
rect 14112 8188 14176 8192
rect 14112 8132 14116 8188
rect 14116 8132 14172 8188
rect 14172 8132 14176 8188
rect 14112 8128 14176 8132
rect 14192 8188 14256 8192
rect 14192 8132 14196 8188
rect 14196 8132 14252 8188
rect 14252 8132 14256 8188
rect 14192 8128 14256 8132
rect 19952 8188 20016 8192
rect 19952 8132 19956 8188
rect 19956 8132 20012 8188
rect 20012 8132 20016 8188
rect 19952 8128 20016 8132
rect 20032 8188 20096 8192
rect 20032 8132 20036 8188
rect 20036 8132 20092 8188
rect 20092 8132 20096 8188
rect 20032 8128 20096 8132
rect 20112 8188 20176 8192
rect 20112 8132 20116 8188
rect 20116 8132 20172 8188
rect 20172 8132 20176 8188
rect 20112 8128 20176 8132
rect 20192 8188 20256 8192
rect 20192 8132 20196 8188
rect 20196 8132 20252 8188
rect 20252 8132 20256 8188
rect 20192 8128 20256 8132
rect 25952 8188 26016 8192
rect 25952 8132 25956 8188
rect 25956 8132 26012 8188
rect 26012 8132 26016 8188
rect 25952 8128 26016 8132
rect 26032 8188 26096 8192
rect 26032 8132 26036 8188
rect 26036 8132 26092 8188
rect 26092 8132 26096 8188
rect 26032 8128 26096 8132
rect 26112 8188 26176 8192
rect 26112 8132 26116 8188
rect 26116 8132 26172 8188
rect 26172 8132 26176 8188
rect 26112 8128 26176 8132
rect 26192 8188 26256 8192
rect 26192 8132 26196 8188
rect 26196 8132 26252 8188
rect 26252 8132 26256 8188
rect 26192 8128 26256 8132
rect 31952 8188 32016 8192
rect 31952 8132 31956 8188
rect 31956 8132 32012 8188
rect 32012 8132 32016 8188
rect 31952 8128 32016 8132
rect 32032 8188 32096 8192
rect 32032 8132 32036 8188
rect 32036 8132 32092 8188
rect 32092 8132 32096 8188
rect 32032 8128 32096 8132
rect 32112 8188 32176 8192
rect 32112 8132 32116 8188
rect 32116 8132 32172 8188
rect 32172 8132 32176 8188
rect 32112 8128 32176 8132
rect 32192 8188 32256 8192
rect 32192 8132 32196 8188
rect 32196 8132 32252 8188
rect 32252 8132 32256 8188
rect 32192 8128 32256 8132
rect 37952 8188 38016 8192
rect 37952 8132 37956 8188
rect 37956 8132 38012 8188
rect 38012 8132 38016 8188
rect 37952 8128 38016 8132
rect 38032 8188 38096 8192
rect 38032 8132 38036 8188
rect 38036 8132 38092 8188
rect 38092 8132 38096 8188
rect 38032 8128 38096 8132
rect 38112 8188 38176 8192
rect 38112 8132 38116 8188
rect 38116 8132 38172 8188
rect 38172 8132 38176 8188
rect 38112 8128 38176 8132
rect 38192 8188 38256 8192
rect 38192 8132 38196 8188
rect 38196 8132 38252 8188
rect 38252 8132 38256 8188
rect 38192 8128 38256 8132
rect 43952 8188 44016 8192
rect 43952 8132 43956 8188
rect 43956 8132 44012 8188
rect 44012 8132 44016 8188
rect 43952 8128 44016 8132
rect 44032 8188 44096 8192
rect 44032 8132 44036 8188
rect 44036 8132 44092 8188
rect 44092 8132 44096 8188
rect 44032 8128 44096 8132
rect 44112 8188 44176 8192
rect 44112 8132 44116 8188
rect 44116 8132 44172 8188
rect 44172 8132 44176 8188
rect 44112 8128 44176 8132
rect 44192 8188 44256 8192
rect 44192 8132 44196 8188
rect 44196 8132 44252 8188
rect 44252 8132 44256 8188
rect 44192 8128 44256 8132
rect 3012 7644 3076 7648
rect 3012 7588 3016 7644
rect 3016 7588 3072 7644
rect 3072 7588 3076 7644
rect 3012 7584 3076 7588
rect 3092 7644 3156 7648
rect 3092 7588 3096 7644
rect 3096 7588 3152 7644
rect 3152 7588 3156 7644
rect 3092 7584 3156 7588
rect 3172 7644 3236 7648
rect 3172 7588 3176 7644
rect 3176 7588 3232 7644
rect 3232 7588 3236 7644
rect 3172 7584 3236 7588
rect 3252 7644 3316 7648
rect 3252 7588 3256 7644
rect 3256 7588 3312 7644
rect 3312 7588 3316 7644
rect 3252 7584 3316 7588
rect 9012 7644 9076 7648
rect 9012 7588 9016 7644
rect 9016 7588 9072 7644
rect 9072 7588 9076 7644
rect 9012 7584 9076 7588
rect 9092 7644 9156 7648
rect 9092 7588 9096 7644
rect 9096 7588 9152 7644
rect 9152 7588 9156 7644
rect 9092 7584 9156 7588
rect 9172 7644 9236 7648
rect 9172 7588 9176 7644
rect 9176 7588 9232 7644
rect 9232 7588 9236 7644
rect 9172 7584 9236 7588
rect 9252 7644 9316 7648
rect 9252 7588 9256 7644
rect 9256 7588 9312 7644
rect 9312 7588 9316 7644
rect 9252 7584 9316 7588
rect 15012 7644 15076 7648
rect 15012 7588 15016 7644
rect 15016 7588 15072 7644
rect 15072 7588 15076 7644
rect 15012 7584 15076 7588
rect 15092 7644 15156 7648
rect 15092 7588 15096 7644
rect 15096 7588 15152 7644
rect 15152 7588 15156 7644
rect 15092 7584 15156 7588
rect 15172 7644 15236 7648
rect 15172 7588 15176 7644
rect 15176 7588 15232 7644
rect 15232 7588 15236 7644
rect 15172 7584 15236 7588
rect 15252 7644 15316 7648
rect 15252 7588 15256 7644
rect 15256 7588 15312 7644
rect 15312 7588 15316 7644
rect 15252 7584 15316 7588
rect 21012 7644 21076 7648
rect 21012 7588 21016 7644
rect 21016 7588 21072 7644
rect 21072 7588 21076 7644
rect 21012 7584 21076 7588
rect 21092 7644 21156 7648
rect 21092 7588 21096 7644
rect 21096 7588 21152 7644
rect 21152 7588 21156 7644
rect 21092 7584 21156 7588
rect 21172 7644 21236 7648
rect 21172 7588 21176 7644
rect 21176 7588 21232 7644
rect 21232 7588 21236 7644
rect 21172 7584 21236 7588
rect 21252 7644 21316 7648
rect 21252 7588 21256 7644
rect 21256 7588 21312 7644
rect 21312 7588 21316 7644
rect 21252 7584 21316 7588
rect 27012 7644 27076 7648
rect 27012 7588 27016 7644
rect 27016 7588 27072 7644
rect 27072 7588 27076 7644
rect 27012 7584 27076 7588
rect 27092 7644 27156 7648
rect 27092 7588 27096 7644
rect 27096 7588 27152 7644
rect 27152 7588 27156 7644
rect 27092 7584 27156 7588
rect 27172 7644 27236 7648
rect 27172 7588 27176 7644
rect 27176 7588 27232 7644
rect 27232 7588 27236 7644
rect 27172 7584 27236 7588
rect 27252 7644 27316 7648
rect 27252 7588 27256 7644
rect 27256 7588 27312 7644
rect 27312 7588 27316 7644
rect 27252 7584 27316 7588
rect 33012 7644 33076 7648
rect 33012 7588 33016 7644
rect 33016 7588 33072 7644
rect 33072 7588 33076 7644
rect 33012 7584 33076 7588
rect 33092 7644 33156 7648
rect 33092 7588 33096 7644
rect 33096 7588 33152 7644
rect 33152 7588 33156 7644
rect 33092 7584 33156 7588
rect 33172 7644 33236 7648
rect 33172 7588 33176 7644
rect 33176 7588 33232 7644
rect 33232 7588 33236 7644
rect 33172 7584 33236 7588
rect 33252 7644 33316 7648
rect 33252 7588 33256 7644
rect 33256 7588 33312 7644
rect 33312 7588 33316 7644
rect 33252 7584 33316 7588
rect 39012 7644 39076 7648
rect 39012 7588 39016 7644
rect 39016 7588 39072 7644
rect 39072 7588 39076 7644
rect 39012 7584 39076 7588
rect 39092 7644 39156 7648
rect 39092 7588 39096 7644
rect 39096 7588 39152 7644
rect 39152 7588 39156 7644
rect 39092 7584 39156 7588
rect 39172 7644 39236 7648
rect 39172 7588 39176 7644
rect 39176 7588 39232 7644
rect 39232 7588 39236 7644
rect 39172 7584 39236 7588
rect 39252 7644 39316 7648
rect 39252 7588 39256 7644
rect 39256 7588 39312 7644
rect 39312 7588 39316 7644
rect 39252 7584 39316 7588
rect 45012 7644 45076 7648
rect 45012 7588 45016 7644
rect 45016 7588 45072 7644
rect 45072 7588 45076 7644
rect 45012 7584 45076 7588
rect 45092 7644 45156 7648
rect 45092 7588 45096 7644
rect 45096 7588 45152 7644
rect 45152 7588 45156 7644
rect 45092 7584 45156 7588
rect 45172 7644 45236 7648
rect 45172 7588 45176 7644
rect 45176 7588 45232 7644
rect 45232 7588 45236 7644
rect 45172 7584 45236 7588
rect 45252 7644 45316 7648
rect 45252 7588 45256 7644
rect 45256 7588 45312 7644
rect 45312 7588 45316 7644
rect 45252 7584 45316 7588
rect 14780 7380 14844 7444
rect 1952 7100 2016 7104
rect 1952 7044 1956 7100
rect 1956 7044 2012 7100
rect 2012 7044 2016 7100
rect 1952 7040 2016 7044
rect 2032 7100 2096 7104
rect 2032 7044 2036 7100
rect 2036 7044 2092 7100
rect 2092 7044 2096 7100
rect 2032 7040 2096 7044
rect 2112 7100 2176 7104
rect 2112 7044 2116 7100
rect 2116 7044 2172 7100
rect 2172 7044 2176 7100
rect 2112 7040 2176 7044
rect 2192 7100 2256 7104
rect 2192 7044 2196 7100
rect 2196 7044 2252 7100
rect 2252 7044 2256 7100
rect 2192 7040 2256 7044
rect 7952 7100 8016 7104
rect 7952 7044 7956 7100
rect 7956 7044 8012 7100
rect 8012 7044 8016 7100
rect 7952 7040 8016 7044
rect 8032 7100 8096 7104
rect 8032 7044 8036 7100
rect 8036 7044 8092 7100
rect 8092 7044 8096 7100
rect 8032 7040 8096 7044
rect 8112 7100 8176 7104
rect 8112 7044 8116 7100
rect 8116 7044 8172 7100
rect 8172 7044 8176 7100
rect 8112 7040 8176 7044
rect 8192 7100 8256 7104
rect 8192 7044 8196 7100
rect 8196 7044 8252 7100
rect 8252 7044 8256 7100
rect 8192 7040 8256 7044
rect 13952 7100 14016 7104
rect 13952 7044 13956 7100
rect 13956 7044 14012 7100
rect 14012 7044 14016 7100
rect 13952 7040 14016 7044
rect 14032 7100 14096 7104
rect 14032 7044 14036 7100
rect 14036 7044 14092 7100
rect 14092 7044 14096 7100
rect 14032 7040 14096 7044
rect 14112 7100 14176 7104
rect 14112 7044 14116 7100
rect 14116 7044 14172 7100
rect 14172 7044 14176 7100
rect 14112 7040 14176 7044
rect 14192 7100 14256 7104
rect 14192 7044 14196 7100
rect 14196 7044 14252 7100
rect 14252 7044 14256 7100
rect 14192 7040 14256 7044
rect 19952 7100 20016 7104
rect 19952 7044 19956 7100
rect 19956 7044 20012 7100
rect 20012 7044 20016 7100
rect 19952 7040 20016 7044
rect 20032 7100 20096 7104
rect 20032 7044 20036 7100
rect 20036 7044 20092 7100
rect 20092 7044 20096 7100
rect 20032 7040 20096 7044
rect 20112 7100 20176 7104
rect 20112 7044 20116 7100
rect 20116 7044 20172 7100
rect 20172 7044 20176 7100
rect 20112 7040 20176 7044
rect 20192 7100 20256 7104
rect 20192 7044 20196 7100
rect 20196 7044 20252 7100
rect 20252 7044 20256 7100
rect 20192 7040 20256 7044
rect 25952 7100 26016 7104
rect 25952 7044 25956 7100
rect 25956 7044 26012 7100
rect 26012 7044 26016 7100
rect 25952 7040 26016 7044
rect 26032 7100 26096 7104
rect 26032 7044 26036 7100
rect 26036 7044 26092 7100
rect 26092 7044 26096 7100
rect 26032 7040 26096 7044
rect 26112 7100 26176 7104
rect 26112 7044 26116 7100
rect 26116 7044 26172 7100
rect 26172 7044 26176 7100
rect 26112 7040 26176 7044
rect 26192 7100 26256 7104
rect 26192 7044 26196 7100
rect 26196 7044 26252 7100
rect 26252 7044 26256 7100
rect 26192 7040 26256 7044
rect 31952 7100 32016 7104
rect 31952 7044 31956 7100
rect 31956 7044 32012 7100
rect 32012 7044 32016 7100
rect 31952 7040 32016 7044
rect 32032 7100 32096 7104
rect 32032 7044 32036 7100
rect 32036 7044 32092 7100
rect 32092 7044 32096 7100
rect 32032 7040 32096 7044
rect 32112 7100 32176 7104
rect 32112 7044 32116 7100
rect 32116 7044 32172 7100
rect 32172 7044 32176 7100
rect 32112 7040 32176 7044
rect 32192 7100 32256 7104
rect 32192 7044 32196 7100
rect 32196 7044 32252 7100
rect 32252 7044 32256 7100
rect 32192 7040 32256 7044
rect 37952 7100 38016 7104
rect 37952 7044 37956 7100
rect 37956 7044 38012 7100
rect 38012 7044 38016 7100
rect 37952 7040 38016 7044
rect 38032 7100 38096 7104
rect 38032 7044 38036 7100
rect 38036 7044 38092 7100
rect 38092 7044 38096 7100
rect 38032 7040 38096 7044
rect 38112 7100 38176 7104
rect 38112 7044 38116 7100
rect 38116 7044 38172 7100
rect 38172 7044 38176 7100
rect 38112 7040 38176 7044
rect 38192 7100 38256 7104
rect 38192 7044 38196 7100
rect 38196 7044 38252 7100
rect 38252 7044 38256 7100
rect 38192 7040 38256 7044
rect 43952 7100 44016 7104
rect 43952 7044 43956 7100
rect 43956 7044 44012 7100
rect 44012 7044 44016 7100
rect 43952 7040 44016 7044
rect 44032 7100 44096 7104
rect 44032 7044 44036 7100
rect 44036 7044 44092 7100
rect 44092 7044 44096 7100
rect 44032 7040 44096 7044
rect 44112 7100 44176 7104
rect 44112 7044 44116 7100
rect 44116 7044 44172 7100
rect 44172 7044 44176 7100
rect 44112 7040 44176 7044
rect 44192 7100 44256 7104
rect 44192 7044 44196 7100
rect 44196 7044 44252 7100
rect 44252 7044 44256 7100
rect 44192 7040 44256 7044
rect 3012 6556 3076 6560
rect 3012 6500 3016 6556
rect 3016 6500 3072 6556
rect 3072 6500 3076 6556
rect 3012 6496 3076 6500
rect 3092 6556 3156 6560
rect 3092 6500 3096 6556
rect 3096 6500 3152 6556
rect 3152 6500 3156 6556
rect 3092 6496 3156 6500
rect 3172 6556 3236 6560
rect 3172 6500 3176 6556
rect 3176 6500 3232 6556
rect 3232 6500 3236 6556
rect 3172 6496 3236 6500
rect 3252 6556 3316 6560
rect 3252 6500 3256 6556
rect 3256 6500 3312 6556
rect 3312 6500 3316 6556
rect 3252 6496 3316 6500
rect 9012 6556 9076 6560
rect 9012 6500 9016 6556
rect 9016 6500 9072 6556
rect 9072 6500 9076 6556
rect 9012 6496 9076 6500
rect 9092 6556 9156 6560
rect 9092 6500 9096 6556
rect 9096 6500 9152 6556
rect 9152 6500 9156 6556
rect 9092 6496 9156 6500
rect 9172 6556 9236 6560
rect 9172 6500 9176 6556
rect 9176 6500 9232 6556
rect 9232 6500 9236 6556
rect 9172 6496 9236 6500
rect 9252 6556 9316 6560
rect 9252 6500 9256 6556
rect 9256 6500 9312 6556
rect 9312 6500 9316 6556
rect 9252 6496 9316 6500
rect 15012 6556 15076 6560
rect 15012 6500 15016 6556
rect 15016 6500 15072 6556
rect 15072 6500 15076 6556
rect 15012 6496 15076 6500
rect 15092 6556 15156 6560
rect 15092 6500 15096 6556
rect 15096 6500 15152 6556
rect 15152 6500 15156 6556
rect 15092 6496 15156 6500
rect 15172 6556 15236 6560
rect 15172 6500 15176 6556
rect 15176 6500 15232 6556
rect 15232 6500 15236 6556
rect 15172 6496 15236 6500
rect 15252 6556 15316 6560
rect 15252 6500 15256 6556
rect 15256 6500 15312 6556
rect 15312 6500 15316 6556
rect 15252 6496 15316 6500
rect 21012 6556 21076 6560
rect 21012 6500 21016 6556
rect 21016 6500 21072 6556
rect 21072 6500 21076 6556
rect 21012 6496 21076 6500
rect 21092 6556 21156 6560
rect 21092 6500 21096 6556
rect 21096 6500 21152 6556
rect 21152 6500 21156 6556
rect 21092 6496 21156 6500
rect 21172 6556 21236 6560
rect 21172 6500 21176 6556
rect 21176 6500 21232 6556
rect 21232 6500 21236 6556
rect 21172 6496 21236 6500
rect 21252 6556 21316 6560
rect 21252 6500 21256 6556
rect 21256 6500 21312 6556
rect 21312 6500 21316 6556
rect 21252 6496 21316 6500
rect 27012 6556 27076 6560
rect 27012 6500 27016 6556
rect 27016 6500 27072 6556
rect 27072 6500 27076 6556
rect 27012 6496 27076 6500
rect 27092 6556 27156 6560
rect 27092 6500 27096 6556
rect 27096 6500 27152 6556
rect 27152 6500 27156 6556
rect 27092 6496 27156 6500
rect 27172 6556 27236 6560
rect 27172 6500 27176 6556
rect 27176 6500 27232 6556
rect 27232 6500 27236 6556
rect 27172 6496 27236 6500
rect 27252 6556 27316 6560
rect 27252 6500 27256 6556
rect 27256 6500 27312 6556
rect 27312 6500 27316 6556
rect 27252 6496 27316 6500
rect 33012 6556 33076 6560
rect 33012 6500 33016 6556
rect 33016 6500 33072 6556
rect 33072 6500 33076 6556
rect 33012 6496 33076 6500
rect 33092 6556 33156 6560
rect 33092 6500 33096 6556
rect 33096 6500 33152 6556
rect 33152 6500 33156 6556
rect 33092 6496 33156 6500
rect 33172 6556 33236 6560
rect 33172 6500 33176 6556
rect 33176 6500 33232 6556
rect 33232 6500 33236 6556
rect 33172 6496 33236 6500
rect 33252 6556 33316 6560
rect 33252 6500 33256 6556
rect 33256 6500 33312 6556
rect 33312 6500 33316 6556
rect 33252 6496 33316 6500
rect 39012 6556 39076 6560
rect 39012 6500 39016 6556
rect 39016 6500 39072 6556
rect 39072 6500 39076 6556
rect 39012 6496 39076 6500
rect 39092 6556 39156 6560
rect 39092 6500 39096 6556
rect 39096 6500 39152 6556
rect 39152 6500 39156 6556
rect 39092 6496 39156 6500
rect 39172 6556 39236 6560
rect 39172 6500 39176 6556
rect 39176 6500 39232 6556
rect 39232 6500 39236 6556
rect 39172 6496 39236 6500
rect 39252 6556 39316 6560
rect 39252 6500 39256 6556
rect 39256 6500 39312 6556
rect 39312 6500 39316 6556
rect 39252 6496 39316 6500
rect 45012 6556 45076 6560
rect 45012 6500 45016 6556
rect 45016 6500 45072 6556
rect 45072 6500 45076 6556
rect 45012 6496 45076 6500
rect 45092 6556 45156 6560
rect 45092 6500 45096 6556
rect 45096 6500 45152 6556
rect 45152 6500 45156 6556
rect 45092 6496 45156 6500
rect 45172 6556 45236 6560
rect 45172 6500 45176 6556
rect 45176 6500 45232 6556
rect 45232 6500 45236 6556
rect 45172 6496 45236 6500
rect 45252 6556 45316 6560
rect 45252 6500 45256 6556
rect 45256 6500 45312 6556
rect 45312 6500 45316 6556
rect 45252 6496 45316 6500
rect 9812 6156 9876 6220
rect 1952 6012 2016 6016
rect 1952 5956 1956 6012
rect 1956 5956 2012 6012
rect 2012 5956 2016 6012
rect 1952 5952 2016 5956
rect 2032 6012 2096 6016
rect 2032 5956 2036 6012
rect 2036 5956 2092 6012
rect 2092 5956 2096 6012
rect 2032 5952 2096 5956
rect 2112 6012 2176 6016
rect 2112 5956 2116 6012
rect 2116 5956 2172 6012
rect 2172 5956 2176 6012
rect 2112 5952 2176 5956
rect 2192 6012 2256 6016
rect 2192 5956 2196 6012
rect 2196 5956 2252 6012
rect 2252 5956 2256 6012
rect 2192 5952 2256 5956
rect 7952 6012 8016 6016
rect 7952 5956 7956 6012
rect 7956 5956 8012 6012
rect 8012 5956 8016 6012
rect 7952 5952 8016 5956
rect 8032 6012 8096 6016
rect 8032 5956 8036 6012
rect 8036 5956 8092 6012
rect 8092 5956 8096 6012
rect 8032 5952 8096 5956
rect 8112 6012 8176 6016
rect 8112 5956 8116 6012
rect 8116 5956 8172 6012
rect 8172 5956 8176 6012
rect 8112 5952 8176 5956
rect 8192 6012 8256 6016
rect 8192 5956 8196 6012
rect 8196 5956 8252 6012
rect 8252 5956 8256 6012
rect 8192 5952 8256 5956
rect 13952 6012 14016 6016
rect 13952 5956 13956 6012
rect 13956 5956 14012 6012
rect 14012 5956 14016 6012
rect 13952 5952 14016 5956
rect 14032 6012 14096 6016
rect 14032 5956 14036 6012
rect 14036 5956 14092 6012
rect 14092 5956 14096 6012
rect 14032 5952 14096 5956
rect 14112 6012 14176 6016
rect 14112 5956 14116 6012
rect 14116 5956 14172 6012
rect 14172 5956 14176 6012
rect 14112 5952 14176 5956
rect 14192 6012 14256 6016
rect 14192 5956 14196 6012
rect 14196 5956 14252 6012
rect 14252 5956 14256 6012
rect 14192 5952 14256 5956
rect 19952 6012 20016 6016
rect 19952 5956 19956 6012
rect 19956 5956 20012 6012
rect 20012 5956 20016 6012
rect 19952 5952 20016 5956
rect 20032 6012 20096 6016
rect 20032 5956 20036 6012
rect 20036 5956 20092 6012
rect 20092 5956 20096 6012
rect 20032 5952 20096 5956
rect 20112 6012 20176 6016
rect 20112 5956 20116 6012
rect 20116 5956 20172 6012
rect 20172 5956 20176 6012
rect 20112 5952 20176 5956
rect 20192 6012 20256 6016
rect 20192 5956 20196 6012
rect 20196 5956 20252 6012
rect 20252 5956 20256 6012
rect 20192 5952 20256 5956
rect 25952 6012 26016 6016
rect 25952 5956 25956 6012
rect 25956 5956 26012 6012
rect 26012 5956 26016 6012
rect 25952 5952 26016 5956
rect 26032 6012 26096 6016
rect 26032 5956 26036 6012
rect 26036 5956 26092 6012
rect 26092 5956 26096 6012
rect 26032 5952 26096 5956
rect 26112 6012 26176 6016
rect 26112 5956 26116 6012
rect 26116 5956 26172 6012
rect 26172 5956 26176 6012
rect 26112 5952 26176 5956
rect 26192 6012 26256 6016
rect 26192 5956 26196 6012
rect 26196 5956 26252 6012
rect 26252 5956 26256 6012
rect 26192 5952 26256 5956
rect 31952 6012 32016 6016
rect 31952 5956 31956 6012
rect 31956 5956 32012 6012
rect 32012 5956 32016 6012
rect 31952 5952 32016 5956
rect 32032 6012 32096 6016
rect 32032 5956 32036 6012
rect 32036 5956 32092 6012
rect 32092 5956 32096 6012
rect 32032 5952 32096 5956
rect 32112 6012 32176 6016
rect 32112 5956 32116 6012
rect 32116 5956 32172 6012
rect 32172 5956 32176 6012
rect 32112 5952 32176 5956
rect 32192 6012 32256 6016
rect 32192 5956 32196 6012
rect 32196 5956 32252 6012
rect 32252 5956 32256 6012
rect 32192 5952 32256 5956
rect 37952 6012 38016 6016
rect 37952 5956 37956 6012
rect 37956 5956 38012 6012
rect 38012 5956 38016 6012
rect 37952 5952 38016 5956
rect 38032 6012 38096 6016
rect 38032 5956 38036 6012
rect 38036 5956 38092 6012
rect 38092 5956 38096 6012
rect 38032 5952 38096 5956
rect 38112 6012 38176 6016
rect 38112 5956 38116 6012
rect 38116 5956 38172 6012
rect 38172 5956 38176 6012
rect 38112 5952 38176 5956
rect 38192 6012 38256 6016
rect 38192 5956 38196 6012
rect 38196 5956 38252 6012
rect 38252 5956 38256 6012
rect 38192 5952 38256 5956
rect 43952 6012 44016 6016
rect 43952 5956 43956 6012
rect 43956 5956 44012 6012
rect 44012 5956 44016 6012
rect 43952 5952 44016 5956
rect 44032 6012 44096 6016
rect 44032 5956 44036 6012
rect 44036 5956 44092 6012
rect 44092 5956 44096 6012
rect 44032 5952 44096 5956
rect 44112 6012 44176 6016
rect 44112 5956 44116 6012
rect 44116 5956 44172 6012
rect 44172 5956 44176 6012
rect 44112 5952 44176 5956
rect 44192 6012 44256 6016
rect 44192 5956 44196 6012
rect 44196 5956 44252 6012
rect 44252 5956 44256 6012
rect 44192 5952 44256 5956
rect 3012 5468 3076 5472
rect 3012 5412 3016 5468
rect 3016 5412 3072 5468
rect 3072 5412 3076 5468
rect 3012 5408 3076 5412
rect 3092 5468 3156 5472
rect 3092 5412 3096 5468
rect 3096 5412 3152 5468
rect 3152 5412 3156 5468
rect 3092 5408 3156 5412
rect 3172 5468 3236 5472
rect 3172 5412 3176 5468
rect 3176 5412 3232 5468
rect 3232 5412 3236 5468
rect 3172 5408 3236 5412
rect 3252 5468 3316 5472
rect 3252 5412 3256 5468
rect 3256 5412 3312 5468
rect 3312 5412 3316 5468
rect 3252 5408 3316 5412
rect 9812 5612 9876 5676
rect 9012 5468 9076 5472
rect 9012 5412 9016 5468
rect 9016 5412 9072 5468
rect 9072 5412 9076 5468
rect 9012 5408 9076 5412
rect 9092 5468 9156 5472
rect 9092 5412 9096 5468
rect 9096 5412 9152 5468
rect 9152 5412 9156 5468
rect 9092 5408 9156 5412
rect 9172 5468 9236 5472
rect 9172 5412 9176 5468
rect 9176 5412 9232 5468
rect 9232 5412 9236 5468
rect 9172 5408 9236 5412
rect 9252 5468 9316 5472
rect 9252 5412 9256 5468
rect 9256 5412 9312 5468
rect 9312 5412 9316 5468
rect 9252 5408 9316 5412
rect 14780 5476 14844 5540
rect 15012 5468 15076 5472
rect 15012 5412 15016 5468
rect 15016 5412 15072 5468
rect 15072 5412 15076 5468
rect 15012 5408 15076 5412
rect 15092 5468 15156 5472
rect 15092 5412 15096 5468
rect 15096 5412 15152 5468
rect 15152 5412 15156 5468
rect 15092 5408 15156 5412
rect 15172 5468 15236 5472
rect 15172 5412 15176 5468
rect 15176 5412 15232 5468
rect 15232 5412 15236 5468
rect 15172 5408 15236 5412
rect 15252 5468 15316 5472
rect 15252 5412 15256 5468
rect 15256 5412 15312 5468
rect 15312 5412 15316 5468
rect 15252 5408 15316 5412
rect 21012 5468 21076 5472
rect 21012 5412 21016 5468
rect 21016 5412 21072 5468
rect 21072 5412 21076 5468
rect 21012 5408 21076 5412
rect 21092 5468 21156 5472
rect 21092 5412 21096 5468
rect 21096 5412 21152 5468
rect 21152 5412 21156 5468
rect 21092 5408 21156 5412
rect 21172 5468 21236 5472
rect 21172 5412 21176 5468
rect 21176 5412 21232 5468
rect 21232 5412 21236 5468
rect 21172 5408 21236 5412
rect 21252 5468 21316 5472
rect 21252 5412 21256 5468
rect 21256 5412 21312 5468
rect 21312 5412 21316 5468
rect 21252 5408 21316 5412
rect 27012 5468 27076 5472
rect 27012 5412 27016 5468
rect 27016 5412 27072 5468
rect 27072 5412 27076 5468
rect 27012 5408 27076 5412
rect 27092 5468 27156 5472
rect 27092 5412 27096 5468
rect 27096 5412 27152 5468
rect 27152 5412 27156 5468
rect 27092 5408 27156 5412
rect 27172 5468 27236 5472
rect 27172 5412 27176 5468
rect 27176 5412 27232 5468
rect 27232 5412 27236 5468
rect 27172 5408 27236 5412
rect 27252 5468 27316 5472
rect 27252 5412 27256 5468
rect 27256 5412 27312 5468
rect 27312 5412 27316 5468
rect 27252 5408 27316 5412
rect 33012 5468 33076 5472
rect 33012 5412 33016 5468
rect 33016 5412 33072 5468
rect 33072 5412 33076 5468
rect 33012 5408 33076 5412
rect 33092 5468 33156 5472
rect 33092 5412 33096 5468
rect 33096 5412 33152 5468
rect 33152 5412 33156 5468
rect 33092 5408 33156 5412
rect 33172 5468 33236 5472
rect 33172 5412 33176 5468
rect 33176 5412 33232 5468
rect 33232 5412 33236 5468
rect 33172 5408 33236 5412
rect 33252 5468 33316 5472
rect 33252 5412 33256 5468
rect 33256 5412 33312 5468
rect 33312 5412 33316 5468
rect 33252 5408 33316 5412
rect 39012 5468 39076 5472
rect 39012 5412 39016 5468
rect 39016 5412 39072 5468
rect 39072 5412 39076 5468
rect 39012 5408 39076 5412
rect 39092 5468 39156 5472
rect 39092 5412 39096 5468
rect 39096 5412 39152 5468
rect 39152 5412 39156 5468
rect 39092 5408 39156 5412
rect 39172 5468 39236 5472
rect 39172 5412 39176 5468
rect 39176 5412 39232 5468
rect 39232 5412 39236 5468
rect 39172 5408 39236 5412
rect 39252 5468 39316 5472
rect 39252 5412 39256 5468
rect 39256 5412 39312 5468
rect 39312 5412 39316 5468
rect 39252 5408 39316 5412
rect 45012 5468 45076 5472
rect 45012 5412 45016 5468
rect 45016 5412 45072 5468
rect 45072 5412 45076 5468
rect 45012 5408 45076 5412
rect 45092 5468 45156 5472
rect 45092 5412 45096 5468
rect 45096 5412 45152 5468
rect 45152 5412 45156 5468
rect 45092 5408 45156 5412
rect 45172 5468 45236 5472
rect 45172 5412 45176 5468
rect 45176 5412 45232 5468
rect 45232 5412 45236 5468
rect 45172 5408 45236 5412
rect 45252 5468 45316 5472
rect 45252 5412 45256 5468
rect 45256 5412 45312 5468
rect 45312 5412 45316 5468
rect 45252 5408 45316 5412
rect 1952 4924 2016 4928
rect 1952 4868 1956 4924
rect 1956 4868 2012 4924
rect 2012 4868 2016 4924
rect 1952 4864 2016 4868
rect 2032 4924 2096 4928
rect 2032 4868 2036 4924
rect 2036 4868 2092 4924
rect 2092 4868 2096 4924
rect 2032 4864 2096 4868
rect 2112 4924 2176 4928
rect 2112 4868 2116 4924
rect 2116 4868 2172 4924
rect 2172 4868 2176 4924
rect 2112 4864 2176 4868
rect 2192 4924 2256 4928
rect 2192 4868 2196 4924
rect 2196 4868 2252 4924
rect 2252 4868 2256 4924
rect 2192 4864 2256 4868
rect 7952 4924 8016 4928
rect 7952 4868 7956 4924
rect 7956 4868 8012 4924
rect 8012 4868 8016 4924
rect 7952 4864 8016 4868
rect 8032 4924 8096 4928
rect 8032 4868 8036 4924
rect 8036 4868 8092 4924
rect 8092 4868 8096 4924
rect 8032 4864 8096 4868
rect 8112 4924 8176 4928
rect 8112 4868 8116 4924
rect 8116 4868 8172 4924
rect 8172 4868 8176 4924
rect 8112 4864 8176 4868
rect 8192 4924 8256 4928
rect 8192 4868 8196 4924
rect 8196 4868 8252 4924
rect 8252 4868 8256 4924
rect 8192 4864 8256 4868
rect 13952 4924 14016 4928
rect 13952 4868 13956 4924
rect 13956 4868 14012 4924
rect 14012 4868 14016 4924
rect 13952 4864 14016 4868
rect 14032 4924 14096 4928
rect 14032 4868 14036 4924
rect 14036 4868 14092 4924
rect 14092 4868 14096 4924
rect 14032 4864 14096 4868
rect 14112 4924 14176 4928
rect 14112 4868 14116 4924
rect 14116 4868 14172 4924
rect 14172 4868 14176 4924
rect 14112 4864 14176 4868
rect 14192 4924 14256 4928
rect 14192 4868 14196 4924
rect 14196 4868 14252 4924
rect 14252 4868 14256 4924
rect 14192 4864 14256 4868
rect 19952 4924 20016 4928
rect 19952 4868 19956 4924
rect 19956 4868 20012 4924
rect 20012 4868 20016 4924
rect 19952 4864 20016 4868
rect 20032 4924 20096 4928
rect 20032 4868 20036 4924
rect 20036 4868 20092 4924
rect 20092 4868 20096 4924
rect 20032 4864 20096 4868
rect 20112 4924 20176 4928
rect 20112 4868 20116 4924
rect 20116 4868 20172 4924
rect 20172 4868 20176 4924
rect 20112 4864 20176 4868
rect 20192 4924 20256 4928
rect 20192 4868 20196 4924
rect 20196 4868 20252 4924
rect 20252 4868 20256 4924
rect 20192 4864 20256 4868
rect 25952 4924 26016 4928
rect 25952 4868 25956 4924
rect 25956 4868 26012 4924
rect 26012 4868 26016 4924
rect 25952 4864 26016 4868
rect 26032 4924 26096 4928
rect 26032 4868 26036 4924
rect 26036 4868 26092 4924
rect 26092 4868 26096 4924
rect 26032 4864 26096 4868
rect 26112 4924 26176 4928
rect 26112 4868 26116 4924
rect 26116 4868 26172 4924
rect 26172 4868 26176 4924
rect 26112 4864 26176 4868
rect 26192 4924 26256 4928
rect 26192 4868 26196 4924
rect 26196 4868 26252 4924
rect 26252 4868 26256 4924
rect 26192 4864 26256 4868
rect 31952 4924 32016 4928
rect 31952 4868 31956 4924
rect 31956 4868 32012 4924
rect 32012 4868 32016 4924
rect 31952 4864 32016 4868
rect 32032 4924 32096 4928
rect 32032 4868 32036 4924
rect 32036 4868 32092 4924
rect 32092 4868 32096 4924
rect 32032 4864 32096 4868
rect 32112 4924 32176 4928
rect 32112 4868 32116 4924
rect 32116 4868 32172 4924
rect 32172 4868 32176 4924
rect 32112 4864 32176 4868
rect 32192 4924 32256 4928
rect 32192 4868 32196 4924
rect 32196 4868 32252 4924
rect 32252 4868 32256 4924
rect 32192 4864 32256 4868
rect 37952 4924 38016 4928
rect 37952 4868 37956 4924
rect 37956 4868 38012 4924
rect 38012 4868 38016 4924
rect 37952 4864 38016 4868
rect 38032 4924 38096 4928
rect 38032 4868 38036 4924
rect 38036 4868 38092 4924
rect 38092 4868 38096 4924
rect 38032 4864 38096 4868
rect 38112 4924 38176 4928
rect 38112 4868 38116 4924
rect 38116 4868 38172 4924
rect 38172 4868 38176 4924
rect 38112 4864 38176 4868
rect 38192 4924 38256 4928
rect 38192 4868 38196 4924
rect 38196 4868 38252 4924
rect 38252 4868 38256 4924
rect 38192 4864 38256 4868
rect 43952 4924 44016 4928
rect 43952 4868 43956 4924
rect 43956 4868 44012 4924
rect 44012 4868 44016 4924
rect 43952 4864 44016 4868
rect 44032 4924 44096 4928
rect 44032 4868 44036 4924
rect 44036 4868 44092 4924
rect 44092 4868 44096 4924
rect 44032 4864 44096 4868
rect 44112 4924 44176 4928
rect 44112 4868 44116 4924
rect 44116 4868 44172 4924
rect 44172 4868 44176 4924
rect 44112 4864 44176 4868
rect 44192 4924 44256 4928
rect 44192 4868 44196 4924
rect 44196 4868 44252 4924
rect 44252 4868 44256 4924
rect 44192 4864 44256 4868
rect 3012 4380 3076 4384
rect 3012 4324 3016 4380
rect 3016 4324 3072 4380
rect 3072 4324 3076 4380
rect 3012 4320 3076 4324
rect 3092 4380 3156 4384
rect 3092 4324 3096 4380
rect 3096 4324 3152 4380
rect 3152 4324 3156 4380
rect 3092 4320 3156 4324
rect 3172 4380 3236 4384
rect 3172 4324 3176 4380
rect 3176 4324 3232 4380
rect 3232 4324 3236 4380
rect 3172 4320 3236 4324
rect 3252 4380 3316 4384
rect 3252 4324 3256 4380
rect 3256 4324 3312 4380
rect 3312 4324 3316 4380
rect 3252 4320 3316 4324
rect 9012 4380 9076 4384
rect 9012 4324 9016 4380
rect 9016 4324 9072 4380
rect 9072 4324 9076 4380
rect 9012 4320 9076 4324
rect 9092 4380 9156 4384
rect 9092 4324 9096 4380
rect 9096 4324 9152 4380
rect 9152 4324 9156 4380
rect 9092 4320 9156 4324
rect 9172 4380 9236 4384
rect 9172 4324 9176 4380
rect 9176 4324 9232 4380
rect 9232 4324 9236 4380
rect 9172 4320 9236 4324
rect 9252 4380 9316 4384
rect 9252 4324 9256 4380
rect 9256 4324 9312 4380
rect 9312 4324 9316 4380
rect 9252 4320 9316 4324
rect 15012 4380 15076 4384
rect 15012 4324 15016 4380
rect 15016 4324 15072 4380
rect 15072 4324 15076 4380
rect 15012 4320 15076 4324
rect 15092 4380 15156 4384
rect 15092 4324 15096 4380
rect 15096 4324 15152 4380
rect 15152 4324 15156 4380
rect 15092 4320 15156 4324
rect 15172 4380 15236 4384
rect 15172 4324 15176 4380
rect 15176 4324 15232 4380
rect 15232 4324 15236 4380
rect 15172 4320 15236 4324
rect 15252 4380 15316 4384
rect 15252 4324 15256 4380
rect 15256 4324 15312 4380
rect 15312 4324 15316 4380
rect 15252 4320 15316 4324
rect 21012 4380 21076 4384
rect 21012 4324 21016 4380
rect 21016 4324 21072 4380
rect 21072 4324 21076 4380
rect 21012 4320 21076 4324
rect 21092 4380 21156 4384
rect 21092 4324 21096 4380
rect 21096 4324 21152 4380
rect 21152 4324 21156 4380
rect 21092 4320 21156 4324
rect 21172 4380 21236 4384
rect 21172 4324 21176 4380
rect 21176 4324 21232 4380
rect 21232 4324 21236 4380
rect 21172 4320 21236 4324
rect 21252 4380 21316 4384
rect 21252 4324 21256 4380
rect 21256 4324 21312 4380
rect 21312 4324 21316 4380
rect 21252 4320 21316 4324
rect 27012 4380 27076 4384
rect 27012 4324 27016 4380
rect 27016 4324 27072 4380
rect 27072 4324 27076 4380
rect 27012 4320 27076 4324
rect 27092 4380 27156 4384
rect 27092 4324 27096 4380
rect 27096 4324 27152 4380
rect 27152 4324 27156 4380
rect 27092 4320 27156 4324
rect 27172 4380 27236 4384
rect 27172 4324 27176 4380
rect 27176 4324 27232 4380
rect 27232 4324 27236 4380
rect 27172 4320 27236 4324
rect 27252 4380 27316 4384
rect 27252 4324 27256 4380
rect 27256 4324 27312 4380
rect 27312 4324 27316 4380
rect 27252 4320 27316 4324
rect 33012 4380 33076 4384
rect 33012 4324 33016 4380
rect 33016 4324 33072 4380
rect 33072 4324 33076 4380
rect 33012 4320 33076 4324
rect 33092 4380 33156 4384
rect 33092 4324 33096 4380
rect 33096 4324 33152 4380
rect 33152 4324 33156 4380
rect 33092 4320 33156 4324
rect 33172 4380 33236 4384
rect 33172 4324 33176 4380
rect 33176 4324 33232 4380
rect 33232 4324 33236 4380
rect 33172 4320 33236 4324
rect 33252 4380 33316 4384
rect 33252 4324 33256 4380
rect 33256 4324 33312 4380
rect 33312 4324 33316 4380
rect 33252 4320 33316 4324
rect 39012 4380 39076 4384
rect 39012 4324 39016 4380
rect 39016 4324 39072 4380
rect 39072 4324 39076 4380
rect 39012 4320 39076 4324
rect 39092 4380 39156 4384
rect 39092 4324 39096 4380
rect 39096 4324 39152 4380
rect 39152 4324 39156 4380
rect 39092 4320 39156 4324
rect 39172 4380 39236 4384
rect 39172 4324 39176 4380
rect 39176 4324 39232 4380
rect 39232 4324 39236 4380
rect 39172 4320 39236 4324
rect 39252 4380 39316 4384
rect 39252 4324 39256 4380
rect 39256 4324 39312 4380
rect 39312 4324 39316 4380
rect 39252 4320 39316 4324
rect 45012 4380 45076 4384
rect 45012 4324 45016 4380
rect 45016 4324 45072 4380
rect 45072 4324 45076 4380
rect 45012 4320 45076 4324
rect 45092 4380 45156 4384
rect 45092 4324 45096 4380
rect 45096 4324 45152 4380
rect 45152 4324 45156 4380
rect 45092 4320 45156 4324
rect 45172 4380 45236 4384
rect 45172 4324 45176 4380
rect 45176 4324 45232 4380
rect 45232 4324 45236 4380
rect 45172 4320 45236 4324
rect 45252 4380 45316 4384
rect 45252 4324 45256 4380
rect 45256 4324 45312 4380
rect 45312 4324 45316 4380
rect 45252 4320 45316 4324
rect 1952 3836 2016 3840
rect 1952 3780 1956 3836
rect 1956 3780 2012 3836
rect 2012 3780 2016 3836
rect 1952 3776 2016 3780
rect 2032 3836 2096 3840
rect 2032 3780 2036 3836
rect 2036 3780 2092 3836
rect 2092 3780 2096 3836
rect 2032 3776 2096 3780
rect 2112 3836 2176 3840
rect 2112 3780 2116 3836
rect 2116 3780 2172 3836
rect 2172 3780 2176 3836
rect 2112 3776 2176 3780
rect 2192 3836 2256 3840
rect 2192 3780 2196 3836
rect 2196 3780 2252 3836
rect 2252 3780 2256 3836
rect 2192 3776 2256 3780
rect 7952 3836 8016 3840
rect 7952 3780 7956 3836
rect 7956 3780 8012 3836
rect 8012 3780 8016 3836
rect 7952 3776 8016 3780
rect 8032 3836 8096 3840
rect 8032 3780 8036 3836
rect 8036 3780 8092 3836
rect 8092 3780 8096 3836
rect 8032 3776 8096 3780
rect 8112 3836 8176 3840
rect 8112 3780 8116 3836
rect 8116 3780 8172 3836
rect 8172 3780 8176 3836
rect 8112 3776 8176 3780
rect 8192 3836 8256 3840
rect 8192 3780 8196 3836
rect 8196 3780 8252 3836
rect 8252 3780 8256 3836
rect 8192 3776 8256 3780
rect 13952 3836 14016 3840
rect 13952 3780 13956 3836
rect 13956 3780 14012 3836
rect 14012 3780 14016 3836
rect 13952 3776 14016 3780
rect 14032 3836 14096 3840
rect 14032 3780 14036 3836
rect 14036 3780 14092 3836
rect 14092 3780 14096 3836
rect 14032 3776 14096 3780
rect 14112 3836 14176 3840
rect 14112 3780 14116 3836
rect 14116 3780 14172 3836
rect 14172 3780 14176 3836
rect 14112 3776 14176 3780
rect 14192 3836 14256 3840
rect 14192 3780 14196 3836
rect 14196 3780 14252 3836
rect 14252 3780 14256 3836
rect 14192 3776 14256 3780
rect 19952 3836 20016 3840
rect 19952 3780 19956 3836
rect 19956 3780 20012 3836
rect 20012 3780 20016 3836
rect 19952 3776 20016 3780
rect 20032 3836 20096 3840
rect 20032 3780 20036 3836
rect 20036 3780 20092 3836
rect 20092 3780 20096 3836
rect 20032 3776 20096 3780
rect 20112 3836 20176 3840
rect 20112 3780 20116 3836
rect 20116 3780 20172 3836
rect 20172 3780 20176 3836
rect 20112 3776 20176 3780
rect 20192 3836 20256 3840
rect 20192 3780 20196 3836
rect 20196 3780 20252 3836
rect 20252 3780 20256 3836
rect 20192 3776 20256 3780
rect 25952 3836 26016 3840
rect 25952 3780 25956 3836
rect 25956 3780 26012 3836
rect 26012 3780 26016 3836
rect 25952 3776 26016 3780
rect 26032 3836 26096 3840
rect 26032 3780 26036 3836
rect 26036 3780 26092 3836
rect 26092 3780 26096 3836
rect 26032 3776 26096 3780
rect 26112 3836 26176 3840
rect 26112 3780 26116 3836
rect 26116 3780 26172 3836
rect 26172 3780 26176 3836
rect 26112 3776 26176 3780
rect 26192 3836 26256 3840
rect 26192 3780 26196 3836
rect 26196 3780 26252 3836
rect 26252 3780 26256 3836
rect 26192 3776 26256 3780
rect 31952 3836 32016 3840
rect 31952 3780 31956 3836
rect 31956 3780 32012 3836
rect 32012 3780 32016 3836
rect 31952 3776 32016 3780
rect 32032 3836 32096 3840
rect 32032 3780 32036 3836
rect 32036 3780 32092 3836
rect 32092 3780 32096 3836
rect 32032 3776 32096 3780
rect 32112 3836 32176 3840
rect 32112 3780 32116 3836
rect 32116 3780 32172 3836
rect 32172 3780 32176 3836
rect 32112 3776 32176 3780
rect 32192 3836 32256 3840
rect 32192 3780 32196 3836
rect 32196 3780 32252 3836
rect 32252 3780 32256 3836
rect 32192 3776 32256 3780
rect 37952 3836 38016 3840
rect 37952 3780 37956 3836
rect 37956 3780 38012 3836
rect 38012 3780 38016 3836
rect 37952 3776 38016 3780
rect 38032 3836 38096 3840
rect 38032 3780 38036 3836
rect 38036 3780 38092 3836
rect 38092 3780 38096 3836
rect 38032 3776 38096 3780
rect 38112 3836 38176 3840
rect 38112 3780 38116 3836
rect 38116 3780 38172 3836
rect 38172 3780 38176 3836
rect 38112 3776 38176 3780
rect 38192 3836 38256 3840
rect 38192 3780 38196 3836
rect 38196 3780 38252 3836
rect 38252 3780 38256 3836
rect 38192 3776 38256 3780
rect 43952 3836 44016 3840
rect 43952 3780 43956 3836
rect 43956 3780 44012 3836
rect 44012 3780 44016 3836
rect 43952 3776 44016 3780
rect 44032 3836 44096 3840
rect 44032 3780 44036 3836
rect 44036 3780 44092 3836
rect 44092 3780 44096 3836
rect 44032 3776 44096 3780
rect 44112 3836 44176 3840
rect 44112 3780 44116 3836
rect 44116 3780 44172 3836
rect 44172 3780 44176 3836
rect 44112 3776 44176 3780
rect 44192 3836 44256 3840
rect 44192 3780 44196 3836
rect 44196 3780 44252 3836
rect 44252 3780 44256 3836
rect 44192 3776 44256 3780
rect 3012 3292 3076 3296
rect 3012 3236 3016 3292
rect 3016 3236 3072 3292
rect 3072 3236 3076 3292
rect 3012 3232 3076 3236
rect 3092 3292 3156 3296
rect 3092 3236 3096 3292
rect 3096 3236 3152 3292
rect 3152 3236 3156 3292
rect 3092 3232 3156 3236
rect 3172 3292 3236 3296
rect 3172 3236 3176 3292
rect 3176 3236 3232 3292
rect 3232 3236 3236 3292
rect 3172 3232 3236 3236
rect 3252 3292 3316 3296
rect 3252 3236 3256 3292
rect 3256 3236 3312 3292
rect 3312 3236 3316 3292
rect 3252 3232 3316 3236
rect 9012 3292 9076 3296
rect 9012 3236 9016 3292
rect 9016 3236 9072 3292
rect 9072 3236 9076 3292
rect 9012 3232 9076 3236
rect 9092 3292 9156 3296
rect 9092 3236 9096 3292
rect 9096 3236 9152 3292
rect 9152 3236 9156 3292
rect 9092 3232 9156 3236
rect 9172 3292 9236 3296
rect 9172 3236 9176 3292
rect 9176 3236 9232 3292
rect 9232 3236 9236 3292
rect 9172 3232 9236 3236
rect 9252 3292 9316 3296
rect 9252 3236 9256 3292
rect 9256 3236 9312 3292
rect 9312 3236 9316 3292
rect 9252 3232 9316 3236
rect 15012 3292 15076 3296
rect 15012 3236 15016 3292
rect 15016 3236 15072 3292
rect 15072 3236 15076 3292
rect 15012 3232 15076 3236
rect 15092 3292 15156 3296
rect 15092 3236 15096 3292
rect 15096 3236 15152 3292
rect 15152 3236 15156 3292
rect 15092 3232 15156 3236
rect 15172 3292 15236 3296
rect 15172 3236 15176 3292
rect 15176 3236 15232 3292
rect 15232 3236 15236 3292
rect 15172 3232 15236 3236
rect 15252 3292 15316 3296
rect 15252 3236 15256 3292
rect 15256 3236 15312 3292
rect 15312 3236 15316 3292
rect 15252 3232 15316 3236
rect 21012 3292 21076 3296
rect 21012 3236 21016 3292
rect 21016 3236 21072 3292
rect 21072 3236 21076 3292
rect 21012 3232 21076 3236
rect 21092 3292 21156 3296
rect 21092 3236 21096 3292
rect 21096 3236 21152 3292
rect 21152 3236 21156 3292
rect 21092 3232 21156 3236
rect 21172 3292 21236 3296
rect 21172 3236 21176 3292
rect 21176 3236 21232 3292
rect 21232 3236 21236 3292
rect 21172 3232 21236 3236
rect 21252 3292 21316 3296
rect 21252 3236 21256 3292
rect 21256 3236 21312 3292
rect 21312 3236 21316 3292
rect 21252 3232 21316 3236
rect 27012 3292 27076 3296
rect 27012 3236 27016 3292
rect 27016 3236 27072 3292
rect 27072 3236 27076 3292
rect 27012 3232 27076 3236
rect 27092 3292 27156 3296
rect 27092 3236 27096 3292
rect 27096 3236 27152 3292
rect 27152 3236 27156 3292
rect 27092 3232 27156 3236
rect 27172 3292 27236 3296
rect 27172 3236 27176 3292
rect 27176 3236 27232 3292
rect 27232 3236 27236 3292
rect 27172 3232 27236 3236
rect 27252 3292 27316 3296
rect 27252 3236 27256 3292
rect 27256 3236 27312 3292
rect 27312 3236 27316 3292
rect 27252 3232 27316 3236
rect 33012 3292 33076 3296
rect 33012 3236 33016 3292
rect 33016 3236 33072 3292
rect 33072 3236 33076 3292
rect 33012 3232 33076 3236
rect 33092 3292 33156 3296
rect 33092 3236 33096 3292
rect 33096 3236 33152 3292
rect 33152 3236 33156 3292
rect 33092 3232 33156 3236
rect 33172 3292 33236 3296
rect 33172 3236 33176 3292
rect 33176 3236 33232 3292
rect 33232 3236 33236 3292
rect 33172 3232 33236 3236
rect 33252 3292 33316 3296
rect 33252 3236 33256 3292
rect 33256 3236 33312 3292
rect 33312 3236 33316 3292
rect 33252 3232 33316 3236
rect 39012 3292 39076 3296
rect 39012 3236 39016 3292
rect 39016 3236 39072 3292
rect 39072 3236 39076 3292
rect 39012 3232 39076 3236
rect 39092 3292 39156 3296
rect 39092 3236 39096 3292
rect 39096 3236 39152 3292
rect 39152 3236 39156 3292
rect 39092 3232 39156 3236
rect 39172 3292 39236 3296
rect 39172 3236 39176 3292
rect 39176 3236 39232 3292
rect 39232 3236 39236 3292
rect 39172 3232 39236 3236
rect 39252 3292 39316 3296
rect 39252 3236 39256 3292
rect 39256 3236 39312 3292
rect 39312 3236 39316 3292
rect 39252 3232 39316 3236
rect 45012 3292 45076 3296
rect 45012 3236 45016 3292
rect 45016 3236 45072 3292
rect 45072 3236 45076 3292
rect 45012 3232 45076 3236
rect 45092 3292 45156 3296
rect 45092 3236 45096 3292
rect 45096 3236 45152 3292
rect 45152 3236 45156 3292
rect 45092 3232 45156 3236
rect 45172 3292 45236 3296
rect 45172 3236 45176 3292
rect 45176 3236 45232 3292
rect 45232 3236 45236 3292
rect 45172 3232 45236 3236
rect 45252 3292 45316 3296
rect 45252 3236 45256 3292
rect 45256 3236 45312 3292
rect 45312 3236 45316 3292
rect 45252 3232 45316 3236
rect 1952 2748 2016 2752
rect 1952 2692 1956 2748
rect 1956 2692 2012 2748
rect 2012 2692 2016 2748
rect 1952 2688 2016 2692
rect 2032 2748 2096 2752
rect 2032 2692 2036 2748
rect 2036 2692 2092 2748
rect 2092 2692 2096 2748
rect 2032 2688 2096 2692
rect 2112 2748 2176 2752
rect 2112 2692 2116 2748
rect 2116 2692 2172 2748
rect 2172 2692 2176 2748
rect 2112 2688 2176 2692
rect 2192 2748 2256 2752
rect 2192 2692 2196 2748
rect 2196 2692 2252 2748
rect 2252 2692 2256 2748
rect 2192 2688 2256 2692
rect 7952 2748 8016 2752
rect 7952 2692 7956 2748
rect 7956 2692 8012 2748
rect 8012 2692 8016 2748
rect 7952 2688 8016 2692
rect 8032 2748 8096 2752
rect 8032 2692 8036 2748
rect 8036 2692 8092 2748
rect 8092 2692 8096 2748
rect 8032 2688 8096 2692
rect 8112 2748 8176 2752
rect 8112 2692 8116 2748
rect 8116 2692 8172 2748
rect 8172 2692 8176 2748
rect 8112 2688 8176 2692
rect 8192 2748 8256 2752
rect 8192 2692 8196 2748
rect 8196 2692 8252 2748
rect 8252 2692 8256 2748
rect 8192 2688 8256 2692
rect 13952 2748 14016 2752
rect 13952 2692 13956 2748
rect 13956 2692 14012 2748
rect 14012 2692 14016 2748
rect 13952 2688 14016 2692
rect 14032 2748 14096 2752
rect 14032 2692 14036 2748
rect 14036 2692 14092 2748
rect 14092 2692 14096 2748
rect 14032 2688 14096 2692
rect 14112 2748 14176 2752
rect 14112 2692 14116 2748
rect 14116 2692 14172 2748
rect 14172 2692 14176 2748
rect 14112 2688 14176 2692
rect 14192 2748 14256 2752
rect 14192 2692 14196 2748
rect 14196 2692 14252 2748
rect 14252 2692 14256 2748
rect 14192 2688 14256 2692
rect 19952 2748 20016 2752
rect 19952 2692 19956 2748
rect 19956 2692 20012 2748
rect 20012 2692 20016 2748
rect 19952 2688 20016 2692
rect 20032 2748 20096 2752
rect 20032 2692 20036 2748
rect 20036 2692 20092 2748
rect 20092 2692 20096 2748
rect 20032 2688 20096 2692
rect 20112 2748 20176 2752
rect 20112 2692 20116 2748
rect 20116 2692 20172 2748
rect 20172 2692 20176 2748
rect 20112 2688 20176 2692
rect 20192 2748 20256 2752
rect 20192 2692 20196 2748
rect 20196 2692 20252 2748
rect 20252 2692 20256 2748
rect 20192 2688 20256 2692
rect 25952 2748 26016 2752
rect 25952 2692 25956 2748
rect 25956 2692 26012 2748
rect 26012 2692 26016 2748
rect 25952 2688 26016 2692
rect 26032 2748 26096 2752
rect 26032 2692 26036 2748
rect 26036 2692 26092 2748
rect 26092 2692 26096 2748
rect 26032 2688 26096 2692
rect 26112 2748 26176 2752
rect 26112 2692 26116 2748
rect 26116 2692 26172 2748
rect 26172 2692 26176 2748
rect 26112 2688 26176 2692
rect 26192 2748 26256 2752
rect 26192 2692 26196 2748
rect 26196 2692 26252 2748
rect 26252 2692 26256 2748
rect 26192 2688 26256 2692
rect 31952 2748 32016 2752
rect 31952 2692 31956 2748
rect 31956 2692 32012 2748
rect 32012 2692 32016 2748
rect 31952 2688 32016 2692
rect 32032 2748 32096 2752
rect 32032 2692 32036 2748
rect 32036 2692 32092 2748
rect 32092 2692 32096 2748
rect 32032 2688 32096 2692
rect 32112 2748 32176 2752
rect 32112 2692 32116 2748
rect 32116 2692 32172 2748
rect 32172 2692 32176 2748
rect 32112 2688 32176 2692
rect 32192 2748 32256 2752
rect 32192 2692 32196 2748
rect 32196 2692 32252 2748
rect 32252 2692 32256 2748
rect 32192 2688 32256 2692
rect 37952 2748 38016 2752
rect 37952 2692 37956 2748
rect 37956 2692 38012 2748
rect 38012 2692 38016 2748
rect 37952 2688 38016 2692
rect 38032 2748 38096 2752
rect 38032 2692 38036 2748
rect 38036 2692 38092 2748
rect 38092 2692 38096 2748
rect 38032 2688 38096 2692
rect 38112 2748 38176 2752
rect 38112 2692 38116 2748
rect 38116 2692 38172 2748
rect 38172 2692 38176 2748
rect 38112 2688 38176 2692
rect 38192 2748 38256 2752
rect 38192 2692 38196 2748
rect 38196 2692 38252 2748
rect 38252 2692 38256 2748
rect 38192 2688 38256 2692
rect 43952 2748 44016 2752
rect 43952 2692 43956 2748
rect 43956 2692 44012 2748
rect 44012 2692 44016 2748
rect 43952 2688 44016 2692
rect 44032 2748 44096 2752
rect 44032 2692 44036 2748
rect 44036 2692 44092 2748
rect 44092 2692 44096 2748
rect 44032 2688 44096 2692
rect 44112 2748 44176 2752
rect 44112 2692 44116 2748
rect 44116 2692 44172 2748
rect 44172 2692 44176 2748
rect 44112 2688 44176 2692
rect 44192 2748 44256 2752
rect 44192 2692 44196 2748
rect 44196 2692 44252 2748
rect 44252 2692 44256 2748
rect 44192 2688 44256 2692
rect 3012 2204 3076 2208
rect 3012 2148 3016 2204
rect 3016 2148 3072 2204
rect 3072 2148 3076 2204
rect 3012 2144 3076 2148
rect 3092 2204 3156 2208
rect 3092 2148 3096 2204
rect 3096 2148 3152 2204
rect 3152 2148 3156 2204
rect 3092 2144 3156 2148
rect 3172 2204 3236 2208
rect 3172 2148 3176 2204
rect 3176 2148 3232 2204
rect 3232 2148 3236 2204
rect 3172 2144 3236 2148
rect 3252 2204 3316 2208
rect 3252 2148 3256 2204
rect 3256 2148 3312 2204
rect 3312 2148 3316 2204
rect 3252 2144 3316 2148
rect 9012 2204 9076 2208
rect 9012 2148 9016 2204
rect 9016 2148 9072 2204
rect 9072 2148 9076 2204
rect 9012 2144 9076 2148
rect 9092 2204 9156 2208
rect 9092 2148 9096 2204
rect 9096 2148 9152 2204
rect 9152 2148 9156 2204
rect 9092 2144 9156 2148
rect 9172 2204 9236 2208
rect 9172 2148 9176 2204
rect 9176 2148 9232 2204
rect 9232 2148 9236 2204
rect 9172 2144 9236 2148
rect 9252 2204 9316 2208
rect 9252 2148 9256 2204
rect 9256 2148 9312 2204
rect 9312 2148 9316 2204
rect 9252 2144 9316 2148
rect 15012 2204 15076 2208
rect 15012 2148 15016 2204
rect 15016 2148 15072 2204
rect 15072 2148 15076 2204
rect 15012 2144 15076 2148
rect 15092 2204 15156 2208
rect 15092 2148 15096 2204
rect 15096 2148 15152 2204
rect 15152 2148 15156 2204
rect 15092 2144 15156 2148
rect 15172 2204 15236 2208
rect 15172 2148 15176 2204
rect 15176 2148 15232 2204
rect 15232 2148 15236 2204
rect 15172 2144 15236 2148
rect 15252 2204 15316 2208
rect 15252 2148 15256 2204
rect 15256 2148 15312 2204
rect 15312 2148 15316 2204
rect 15252 2144 15316 2148
rect 21012 2204 21076 2208
rect 21012 2148 21016 2204
rect 21016 2148 21072 2204
rect 21072 2148 21076 2204
rect 21012 2144 21076 2148
rect 21092 2204 21156 2208
rect 21092 2148 21096 2204
rect 21096 2148 21152 2204
rect 21152 2148 21156 2204
rect 21092 2144 21156 2148
rect 21172 2204 21236 2208
rect 21172 2148 21176 2204
rect 21176 2148 21232 2204
rect 21232 2148 21236 2204
rect 21172 2144 21236 2148
rect 21252 2204 21316 2208
rect 21252 2148 21256 2204
rect 21256 2148 21312 2204
rect 21312 2148 21316 2204
rect 21252 2144 21316 2148
rect 27012 2204 27076 2208
rect 27012 2148 27016 2204
rect 27016 2148 27072 2204
rect 27072 2148 27076 2204
rect 27012 2144 27076 2148
rect 27092 2204 27156 2208
rect 27092 2148 27096 2204
rect 27096 2148 27152 2204
rect 27152 2148 27156 2204
rect 27092 2144 27156 2148
rect 27172 2204 27236 2208
rect 27172 2148 27176 2204
rect 27176 2148 27232 2204
rect 27232 2148 27236 2204
rect 27172 2144 27236 2148
rect 27252 2204 27316 2208
rect 27252 2148 27256 2204
rect 27256 2148 27312 2204
rect 27312 2148 27316 2204
rect 27252 2144 27316 2148
rect 33012 2204 33076 2208
rect 33012 2148 33016 2204
rect 33016 2148 33072 2204
rect 33072 2148 33076 2204
rect 33012 2144 33076 2148
rect 33092 2204 33156 2208
rect 33092 2148 33096 2204
rect 33096 2148 33152 2204
rect 33152 2148 33156 2204
rect 33092 2144 33156 2148
rect 33172 2204 33236 2208
rect 33172 2148 33176 2204
rect 33176 2148 33232 2204
rect 33232 2148 33236 2204
rect 33172 2144 33236 2148
rect 33252 2204 33316 2208
rect 33252 2148 33256 2204
rect 33256 2148 33312 2204
rect 33312 2148 33316 2204
rect 33252 2144 33316 2148
rect 39012 2204 39076 2208
rect 39012 2148 39016 2204
rect 39016 2148 39072 2204
rect 39072 2148 39076 2204
rect 39012 2144 39076 2148
rect 39092 2204 39156 2208
rect 39092 2148 39096 2204
rect 39096 2148 39152 2204
rect 39152 2148 39156 2204
rect 39092 2144 39156 2148
rect 39172 2204 39236 2208
rect 39172 2148 39176 2204
rect 39176 2148 39232 2204
rect 39232 2148 39236 2204
rect 39172 2144 39236 2148
rect 39252 2204 39316 2208
rect 39252 2148 39256 2204
rect 39256 2148 39312 2204
rect 39312 2148 39316 2204
rect 39252 2144 39316 2148
rect 45012 2204 45076 2208
rect 45012 2148 45016 2204
rect 45016 2148 45072 2204
rect 45072 2148 45076 2204
rect 45012 2144 45076 2148
rect 45092 2204 45156 2208
rect 45092 2148 45096 2204
rect 45096 2148 45152 2204
rect 45152 2148 45156 2204
rect 45092 2144 45156 2148
rect 45172 2204 45236 2208
rect 45172 2148 45176 2204
rect 45176 2148 45232 2204
rect 45232 2148 45236 2204
rect 45172 2144 45236 2148
rect 45252 2204 45316 2208
rect 45252 2148 45256 2204
rect 45256 2148 45312 2204
rect 45312 2148 45316 2204
rect 45252 2144 45316 2148
<< metal4 >>
rect 1944 8192 2264 11250
rect 1944 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2264 8192
rect 1944 7104 2264 8128
rect 1944 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2264 7104
rect 1944 6016 2264 7040
rect 1944 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2264 6016
rect 1944 4928 2264 5952
rect 1944 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2264 4928
rect 1944 3840 2264 4864
rect 1944 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2264 3840
rect 1944 2752 2264 3776
rect 1944 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2264 2752
rect 1944 0 2264 2688
rect 3004 8736 3324 11250
rect 3004 8672 3012 8736
rect 3076 8672 3092 8736
rect 3156 8672 3172 8736
rect 3236 8672 3252 8736
rect 3316 8672 3324 8736
rect 3004 7648 3324 8672
rect 3004 7584 3012 7648
rect 3076 7584 3092 7648
rect 3156 7584 3172 7648
rect 3236 7584 3252 7648
rect 3316 7584 3324 7648
rect 3004 6560 3324 7584
rect 3004 6496 3012 6560
rect 3076 6496 3092 6560
rect 3156 6496 3172 6560
rect 3236 6496 3252 6560
rect 3316 6496 3324 6560
rect 3004 5472 3324 6496
rect 3004 5408 3012 5472
rect 3076 5408 3092 5472
rect 3156 5408 3172 5472
rect 3236 5408 3252 5472
rect 3316 5408 3324 5472
rect 3004 4384 3324 5408
rect 3004 4320 3012 4384
rect 3076 4320 3092 4384
rect 3156 4320 3172 4384
rect 3236 4320 3252 4384
rect 3316 4320 3324 4384
rect 3004 3296 3324 4320
rect 3004 3232 3012 3296
rect 3076 3232 3092 3296
rect 3156 3232 3172 3296
rect 3236 3232 3252 3296
rect 3316 3232 3324 3296
rect 3004 2208 3324 3232
rect 3004 2144 3012 2208
rect 3076 2144 3092 2208
rect 3156 2144 3172 2208
rect 3236 2144 3252 2208
rect 3316 2144 3324 2208
rect 3004 0 3324 2144
rect 7944 8192 8264 11250
rect 7944 8128 7952 8192
rect 8016 8128 8032 8192
rect 8096 8128 8112 8192
rect 8176 8128 8192 8192
rect 8256 8128 8264 8192
rect 7944 7104 8264 8128
rect 7944 7040 7952 7104
rect 8016 7040 8032 7104
rect 8096 7040 8112 7104
rect 8176 7040 8192 7104
rect 8256 7040 8264 7104
rect 7944 6016 8264 7040
rect 7944 5952 7952 6016
rect 8016 5952 8032 6016
rect 8096 5952 8112 6016
rect 8176 5952 8192 6016
rect 8256 5952 8264 6016
rect 7944 4928 8264 5952
rect 7944 4864 7952 4928
rect 8016 4864 8032 4928
rect 8096 4864 8112 4928
rect 8176 4864 8192 4928
rect 8256 4864 8264 4928
rect 7944 3840 8264 4864
rect 7944 3776 7952 3840
rect 8016 3776 8032 3840
rect 8096 3776 8112 3840
rect 8176 3776 8192 3840
rect 8256 3776 8264 3840
rect 7944 2752 8264 3776
rect 7944 2688 7952 2752
rect 8016 2688 8032 2752
rect 8096 2688 8112 2752
rect 8176 2688 8192 2752
rect 8256 2688 8264 2752
rect 7944 0 8264 2688
rect 9004 8736 9324 11250
rect 9004 8672 9012 8736
rect 9076 8672 9092 8736
rect 9156 8672 9172 8736
rect 9236 8672 9252 8736
rect 9316 8672 9324 8736
rect 9004 7648 9324 8672
rect 9004 7584 9012 7648
rect 9076 7584 9092 7648
rect 9156 7584 9172 7648
rect 9236 7584 9252 7648
rect 9316 7584 9324 7648
rect 9004 6560 9324 7584
rect 9004 6496 9012 6560
rect 9076 6496 9092 6560
rect 9156 6496 9172 6560
rect 9236 6496 9252 6560
rect 9316 6496 9324 6560
rect 9004 5472 9324 6496
rect 13944 8192 14264 11250
rect 13944 8128 13952 8192
rect 14016 8128 14032 8192
rect 14096 8128 14112 8192
rect 14176 8128 14192 8192
rect 14256 8128 14264 8192
rect 13944 7104 14264 8128
rect 15004 8736 15324 11250
rect 15004 8672 15012 8736
rect 15076 8672 15092 8736
rect 15156 8672 15172 8736
rect 15236 8672 15252 8736
rect 15316 8672 15324 8736
rect 15004 7648 15324 8672
rect 15004 7584 15012 7648
rect 15076 7584 15092 7648
rect 15156 7584 15172 7648
rect 15236 7584 15252 7648
rect 15316 7584 15324 7648
rect 14779 7444 14845 7445
rect 14779 7380 14780 7444
rect 14844 7380 14845 7444
rect 14779 7379 14845 7380
rect 13944 7040 13952 7104
rect 14016 7040 14032 7104
rect 14096 7040 14112 7104
rect 14176 7040 14192 7104
rect 14256 7040 14264 7104
rect 9811 6220 9877 6221
rect 9811 6156 9812 6220
rect 9876 6156 9877 6220
rect 9811 6155 9877 6156
rect 9814 5677 9874 6155
rect 13944 6016 14264 7040
rect 13944 5952 13952 6016
rect 14016 5952 14032 6016
rect 14096 5952 14112 6016
rect 14176 5952 14192 6016
rect 14256 5952 14264 6016
rect 9811 5676 9877 5677
rect 9811 5612 9812 5676
rect 9876 5612 9877 5676
rect 9811 5611 9877 5612
rect 9004 5408 9012 5472
rect 9076 5408 9092 5472
rect 9156 5408 9172 5472
rect 9236 5408 9252 5472
rect 9316 5408 9324 5472
rect 9004 4384 9324 5408
rect 9004 4320 9012 4384
rect 9076 4320 9092 4384
rect 9156 4320 9172 4384
rect 9236 4320 9252 4384
rect 9316 4320 9324 4384
rect 9004 3296 9324 4320
rect 9004 3232 9012 3296
rect 9076 3232 9092 3296
rect 9156 3232 9172 3296
rect 9236 3232 9252 3296
rect 9316 3232 9324 3296
rect 9004 2208 9324 3232
rect 9004 2144 9012 2208
rect 9076 2144 9092 2208
rect 9156 2144 9172 2208
rect 9236 2144 9252 2208
rect 9316 2144 9324 2208
rect 9004 0 9324 2144
rect 13944 4928 14264 5952
rect 14782 5541 14842 7379
rect 15004 6560 15324 7584
rect 15004 6496 15012 6560
rect 15076 6496 15092 6560
rect 15156 6496 15172 6560
rect 15236 6496 15252 6560
rect 15316 6496 15324 6560
rect 14779 5540 14845 5541
rect 14779 5476 14780 5540
rect 14844 5476 14845 5540
rect 14779 5475 14845 5476
rect 13944 4864 13952 4928
rect 14016 4864 14032 4928
rect 14096 4864 14112 4928
rect 14176 4864 14192 4928
rect 14256 4864 14264 4928
rect 13944 3840 14264 4864
rect 13944 3776 13952 3840
rect 14016 3776 14032 3840
rect 14096 3776 14112 3840
rect 14176 3776 14192 3840
rect 14256 3776 14264 3840
rect 13944 2752 14264 3776
rect 13944 2688 13952 2752
rect 14016 2688 14032 2752
rect 14096 2688 14112 2752
rect 14176 2688 14192 2752
rect 14256 2688 14264 2752
rect 13944 0 14264 2688
rect 15004 5472 15324 6496
rect 15004 5408 15012 5472
rect 15076 5408 15092 5472
rect 15156 5408 15172 5472
rect 15236 5408 15252 5472
rect 15316 5408 15324 5472
rect 15004 4384 15324 5408
rect 15004 4320 15012 4384
rect 15076 4320 15092 4384
rect 15156 4320 15172 4384
rect 15236 4320 15252 4384
rect 15316 4320 15324 4384
rect 15004 3296 15324 4320
rect 15004 3232 15012 3296
rect 15076 3232 15092 3296
rect 15156 3232 15172 3296
rect 15236 3232 15252 3296
rect 15316 3232 15324 3296
rect 15004 2208 15324 3232
rect 15004 2144 15012 2208
rect 15076 2144 15092 2208
rect 15156 2144 15172 2208
rect 15236 2144 15252 2208
rect 15316 2144 15324 2208
rect 15004 0 15324 2144
rect 19944 8192 20264 11250
rect 19944 8128 19952 8192
rect 20016 8128 20032 8192
rect 20096 8128 20112 8192
rect 20176 8128 20192 8192
rect 20256 8128 20264 8192
rect 19944 7104 20264 8128
rect 19944 7040 19952 7104
rect 20016 7040 20032 7104
rect 20096 7040 20112 7104
rect 20176 7040 20192 7104
rect 20256 7040 20264 7104
rect 19944 6016 20264 7040
rect 19944 5952 19952 6016
rect 20016 5952 20032 6016
rect 20096 5952 20112 6016
rect 20176 5952 20192 6016
rect 20256 5952 20264 6016
rect 19944 4928 20264 5952
rect 19944 4864 19952 4928
rect 20016 4864 20032 4928
rect 20096 4864 20112 4928
rect 20176 4864 20192 4928
rect 20256 4864 20264 4928
rect 19944 3840 20264 4864
rect 19944 3776 19952 3840
rect 20016 3776 20032 3840
rect 20096 3776 20112 3840
rect 20176 3776 20192 3840
rect 20256 3776 20264 3840
rect 19944 2752 20264 3776
rect 19944 2688 19952 2752
rect 20016 2688 20032 2752
rect 20096 2688 20112 2752
rect 20176 2688 20192 2752
rect 20256 2688 20264 2752
rect 19944 0 20264 2688
rect 21004 8736 21324 11250
rect 21004 8672 21012 8736
rect 21076 8672 21092 8736
rect 21156 8672 21172 8736
rect 21236 8672 21252 8736
rect 21316 8672 21324 8736
rect 21004 7648 21324 8672
rect 21004 7584 21012 7648
rect 21076 7584 21092 7648
rect 21156 7584 21172 7648
rect 21236 7584 21252 7648
rect 21316 7584 21324 7648
rect 21004 6560 21324 7584
rect 21004 6496 21012 6560
rect 21076 6496 21092 6560
rect 21156 6496 21172 6560
rect 21236 6496 21252 6560
rect 21316 6496 21324 6560
rect 21004 5472 21324 6496
rect 21004 5408 21012 5472
rect 21076 5408 21092 5472
rect 21156 5408 21172 5472
rect 21236 5408 21252 5472
rect 21316 5408 21324 5472
rect 21004 4384 21324 5408
rect 21004 4320 21012 4384
rect 21076 4320 21092 4384
rect 21156 4320 21172 4384
rect 21236 4320 21252 4384
rect 21316 4320 21324 4384
rect 21004 3296 21324 4320
rect 21004 3232 21012 3296
rect 21076 3232 21092 3296
rect 21156 3232 21172 3296
rect 21236 3232 21252 3296
rect 21316 3232 21324 3296
rect 21004 2208 21324 3232
rect 21004 2144 21012 2208
rect 21076 2144 21092 2208
rect 21156 2144 21172 2208
rect 21236 2144 21252 2208
rect 21316 2144 21324 2208
rect 21004 0 21324 2144
rect 25944 8192 26264 11250
rect 25944 8128 25952 8192
rect 26016 8128 26032 8192
rect 26096 8128 26112 8192
rect 26176 8128 26192 8192
rect 26256 8128 26264 8192
rect 25944 7104 26264 8128
rect 25944 7040 25952 7104
rect 26016 7040 26032 7104
rect 26096 7040 26112 7104
rect 26176 7040 26192 7104
rect 26256 7040 26264 7104
rect 25944 6016 26264 7040
rect 25944 5952 25952 6016
rect 26016 5952 26032 6016
rect 26096 5952 26112 6016
rect 26176 5952 26192 6016
rect 26256 5952 26264 6016
rect 25944 4928 26264 5952
rect 25944 4864 25952 4928
rect 26016 4864 26032 4928
rect 26096 4864 26112 4928
rect 26176 4864 26192 4928
rect 26256 4864 26264 4928
rect 25944 3840 26264 4864
rect 25944 3776 25952 3840
rect 26016 3776 26032 3840
rect 26096 3776 26112 3840
rect 26176 3776 26192 3840
rect 26256 3776 26264 3840
rect 25944 2752 26264 3776
rect 25944 2688 25952 2752
rect 26016 2688 26032 2752
rect 26096 2688 26112 2752
rect 26176 2688 26192 2752
rect 26256 2688 26264 2752
rect 25944 0 26264 2688
rect 27004 8736 27324 11250
rect 27004 8672 27012 8736
rect 27076 8672 27092 8736
rect 27156 8672 27172 8736
rect 27236 8672 27252 8736
rect 27316 8672 27324 8736
rect 27004 7648 27324 8672
rect 27004 7584 27012 7648
rect 27076 7584 27092 7648
rect 27156 7584 27172 7648
rect 27236 7584 27252 7648
rect 27316 7584 27324 7648
rect 27004 6560 27324 7584
rect 27004 6496 27012 6560
rect 27076 6496 27092 6560
rect 27156 6496 27172 6560
rect 27236 6496 27252 6560
rect 27316 6496 27324 6560
rect 27004 5472 27324 6496
rect 27004 5408 27012 5472
rect 27076 5408 27092 5472
rect 27156 5408 27172 5472
rect 27236 5408 27252 5472
rect 27316 5408 27324 5472
rect 27004 4384 27324 5408
rect 27004 4320 27012 4384
rect 27076 4320 27092 4384
rect 27156 4320 27172 4384
rect 27236 4320 27252 4384
rect 27316 4320 27324 4384
rect 27004 3296 27324 4320
rect 27004 3232 27012 3296
rect 27076 3232 27092 3296
rect 27156 3232 27172 3296
rect 27236 3232 27252 3296
rect 27316 3232 27324 3296
rect 27004 2208 27324 3232
rect 27004 2144 27012 2208
rect 27076 2144 27092 2208
rect 27156 2144 27172 2208
rect 27236 2144 27252 2208
rect 27316 2144 27324 2208
rect 27004 0 27324 2144
rect 31944 8192 32264 11250
rect 31944 8128 31952 8192
rect 32016 8128 32032 8192
rect 32096 8128 32112 8192
rect 32176 8128 32192 8192
rect 32256 8128 32264 8192
rect 31944 7104 32264 8128
rect 31944 7040 31952 7104
rect 32016 7040 32032 7104
rect 32096 7040 32112 7104
rect 32176 7040 32192 7104
rect 32256 7040 32264 7104
rect 31944 6016 32264 7040
rect 31944 5952 31952 6016
rect 32016 5952 32032 6016
rect 32096 5952 32112 6016
rect 32176 5952 32192 6016
rect 32256 5952 32264 6016
rect 31944 4928 32264 5952
rect 31944 4864 31952 4928
rect 32016 4864 32032 4928
rect 32096 4864 32112 4928
rect 32176 4864 32192 4928
rect 32256 4864 32264 4928
rect 31944 3840 32264 4864
rect 31944 3776 31952 3840
rect 32016 3776 32032 3840
rect 32096 3776 32112 3840
rect 32176 3776 32192 3840
rect 32256 3776 32264 3840
rect 31944 2752 32264 3776
rect 31944 2688 31952 2752
rect 32016 2688 32032 2752
rect 32096 2688 32112 2752
rect 32176 2688 32192 2752
rect 32256 2688 32264 2752
rect 31944 0 32264 2688
rect 33004 8736 33324 11250
rect 33004 8672 33012 8736
rect 33076 8672 33092 8736
rect 33156 8672 33172 8736
rect 33236 8672 33252 8736
rect 33316 8672 33324 8736
rect 33004 7648 33324 8672
rect 33004 7584 33012 7648
rect 33076 7584 33092 7648
rect 33156 7584 33172 7648
rect 33236 7584 33252 7648
rect 33316 7584 33324 7648
rect 33004 6560 33324 7584
rect 33004 6496 33012 6560
rect 33076 6496 33092 6560
rect 33156 6496 33172 6560
rect 33236 6496 33252 6560
rect 33316 6496 33324 6560
rect 33004 5472 33324 6496
rect 33004 5408 33012 5472
rect 33076 5408 33092 5472
rect 33156 5408 33172 5472
rect 33236 5408 33252 5472
rect 33316 5408 33324 5472
rect 33004 4384 33324 5408
rect 33004 4320 33012 4384
rect 33076 4320 33092 4384
rect 33156 4320 33172 4384
rect 33236 4320 33252 4384
rect 33316 4320 33324 4384
rect 33004 3296 33324 4320
rect 33004 3232 33012 3296
rect 33076 3232 33092 3296
rect 33156 3232 33172 3296
rect 33236 3232 33252 3296
rect 33316 3232 33324 3296
rect 33004 2208 33324 3232
rect 33004 2144 33012 2208
rect 33076 2144 33092 2208
rect 33156 2144 33172 2208
rect 33236 2144 33252 2208
rect 33316 2144 33324 2208
rect 33004 0 33324 2144
rect 37944 8192 38264 11250
rect 37944 8128 37952 8192
rect 38016 8128 38032 8192
rect 38096 8128 38112 8192
rect 38176 8128 38192 8192
rect 38256 8128 38264 8192
rect 37944 7104 38264 8128
rect 37944 7040 37952 7104
rect 38016 7040 38032 7104
rect 38096 7040 38112 7104
rect 38176 7040 38192 7104
rect 38256 7040 38264 7104
rect 37944 6016 38264 7040
rect 37944 5952 37952 6016
rect 38016 5952 38032 6016
rect 38096 5952 38112 6016
rect 38176 5952 38192 6016
rect 38256 5952 38264 6016
rect 37944 4928 38264 5952
rect 37944 4864 37952 4928
rect 38016 4864 38032 4928
rect 38096 4864 38112 4928
rect 38176 4864 38192 4928
rect 38256 4864 38264 4928
rect 37944 3840 38264 4864
rect 37944 3776 37952 3840
rect 38016 3776 38032 3840
rect 38096 3776 38112 3840
rect 38176 3776 38192 3840
rect 38256 3776 38264 3840
rect 37944 2752 38264 3776
rect 37944 2688 37952 2752
rect 38016 2688 38032 2752
rect 38096 2688 38112 2752
rect 38176 2688 38192 2752
rect 38256 2688 38264 2752
rect 37944 0 38264 2688
rect 39004 8736 39324 11250
rect 39004 8672 39012 8736
rect 39076 8672 39092 8736
rect 39156 8672 39172 8736
rect 39236 8672 39252 8736
rect 39316 8672 39324 8736
rect 39004 7648 39324 8672
rect 39004 7584 39012 7648
rect 39076 7584 39092 7648
rect 39156 7584 39172 7648
rect 39236 7584 39252 7648
rect 39316 7584 39324 7648
rect 39004 6560 39324 7584
rect 39004 6496 39012 6560
rect 39076 6496 39092 6560
rect 39156 6496 39172 6560
rect 39236 6496 39252 6560
rect 39316 6496 39324 6560
rect 39004 5472 39324 6496
rect 39004 5408 39012 5472
rect 39076 5408 39092 5472
rect 39156 5408 39172 5472
rect 39236 5408 39252 5472
rect 39316 5408 39324 5472
rect 39004 4384 39324 5408
rect 39004 4320 39012 4384
rect 39076 4320 39092 4384
rect 39156 4320 39172 4384
rect 39236 4320 39252 4384
rect 39316 4320 39324 4384
rect 39004 3296 39324 4320
rect 39004 3232 39012 3296
rect 39076 3232 39092 3296
rect 39156 3232 39172 3296
rect 39236 3232 39252 3296
rect 39316 3232 39324 3296
rect 39004 2208 39324 3232
rect 39004 2144 39012 2208
rect 39076 2144 39092 2208
rect 39156 2144 39172 2208
rect 39236 2144 39252 2208
rect 39316 2144 39324 2208
rect 39004 0 39324 2144
rect 43944 8192 44264 11250
rect 43944 8128 43952 8192
rect 44016 8128 44032 8192
rect 44096 8128 44112 8192
rect 44176 8128 44192 8192
rect 44256 8128 44264 8192
rect 43944 7104 44264 8128
rect 43944 7040 43952 7104
rect 44016 7040 44032 7104
rect 44096 7040 44112 7104
rect 44176 7040 44192 7104
rect 44256 7040 44264 7104
rect 43944 6016 44264 7040
rect 43944 5952 43952 6016
rect 44016 5952 44032 6016
rect 44096 5952 44112 6016
rect 44176 5952 44192 6016
rect 44256 5952 44264 6016
rect 43944 4928 44264 5952
rect 43944 4864 43952 4928
rect 44016 4864 44032 4928
rect 44096 4864 44112 4928
rect 44176 4864 44192 4928
rect 44256 4864 44264 4928
rect 43944 3840 44264 4864
rect 43944 3776 43952 3840
rect 44016 3776 44032 3840
rect 44096 3776 44112 3840
rect 44176 3776 44192 3840
rect 44256 3776 44264 3840
rect 43944 2752 44264 3776
rect 43944 2688 43952 2752
rect 44016 2688 44032 2752
rect 44096 2688 44112 2752
rect 44176 2688 44192 2752
rect 44256 2688 44264 2752
rect 43944 0 44264 2688
rect 45004 8736 45324 11250
rect 45004 8672 45012 8736
rect 45076 8672 45092 8736
rect 45156 8672 45172 8736
rect 45236 8672 45252 8736
rect 45316 8672 45324 8736
rect 45004 7648 45324 8672
rect 45004 7584 45012 7648
rect 45076 7584 45092 7648
rect 45156 7584 45172 7648
rect 45236 7584 45252 7648
rect 45316 7584 45324 7648
rect 45004 6560 45324 7584
rect 45004 6496 45012 6560
rect 45076 6496 45092 6560
rect 45156 6496 45172 6560
rect 45236 6496 45252 6560
rect 45316 6496 45324 6560
rect 45004 5472 45324 6496
rect 45004 5408 45012 5472
rect 45076 5408 45092 5472
rect 45156 5408 45172 5472
rect 45236 5408 45252 5472
rect 45316 5408 45324 5472
rect 45004 4384 45324 5408
rect 45004 4320 45012 4384
rect 45076 4320 45092 4384
rect 45156 4320 45172 4384
rect 45236 4320 45252 4384
rect 45316 4320 45324 4384
rect 45004 3296 45324 4320
rect 45004 3232 45012 3296
rect 45076 3232 45092 3296
rect 45156 3232 45172 3296
rect 45236 3232 45252 3296
rect 45316 3232 45324 3296
rect 45004 2208 45324 3232
rect 45004 2144 45012 2208
rect 45076 2144 45092 2208
rect 45156 2144 45172 2208
rect 45236 2144 45252 2208
rect 45316 2144 45324 2208
rect 45004 0 45324 2144
use sky130_fd_sc_hd__clkbuf_2  _000_
timestamp -3599
transform 1 0 8280 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _001_
timestamp -3599
transform 1 0 12972 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _002_
timestamp -3599
transform 1 0 20240 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _003_
timestamp -3599
transform 1 0 20884 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _004_
timestamp -3599
transform 1 0 16652 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _005_
timestamp -3599
transform 1 0 25116 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _006_
timestamp -3599
transform 1 0 23368 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _007_
timestamp -3599
transform 1 0 22724 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _008_
timestamp -3599
transform 1 0 25024 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _009_
timestamp -3599
transform 1 0 18124 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _010_
timestamp -3599
transform -1 0 25760 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _011_
timestamp -3599
transform 1 0 23460 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _012_
timestamp -3599
transform 1 0 21804 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _013_
timestamp -3599
transform 1 0 21528 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _014_
timestamp -3599
transform 1 0 18584 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _015_
timestamp -3599
transform 1 0 17572 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _016_
timestamp -3599
transform 1 0 20240 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _017_
timestamp -3599
transform 1 0 27508 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _018_
timestamp -3599
transform 1 0 14628 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _019_
timestamp -3599
transform 1 0 25300 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _020_
timestamp -3599
transform 1 0 17848 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _021_
timestamp -3599
transform 1 0 9108 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _022_
timestamp -3599
transform 1 0 37444 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _023_
timestamp -3599
transform 1 0 22908 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _024_
timestamp -3599
transform 1 0 36708 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _025_
timestamp -3599
transform 1 0 32936 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _026_
timestamp -3599
transform -1 0 42044 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _027_
timestamp -3599
transform 1 0 7636 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _028_
timestamp -3599
transform 1 0 30360 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _029_
timestamp -3599
transform 1 0 2116 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _030_
timestamp -3599
transform 1 0 5060 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _031_
timestamp -3599
transform -1 0 46092 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _032_
timestamp -3599
transform -1 0 39744 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _033_
timestamp -3599
transform -1 0 40572 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _034_
timestamp -3599
transform 1 0 8648 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _035_
timestamp -3599
transform 1 0 10764 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _036_
timestamp -3599
transform 1 0 12604 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _037_
timestamp -3599
transform 1 0 15640 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _038_
timestamp -3599
transform 1 0 18676 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _039_
timestamp -3599
transform 1 0 21896 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _040_
timestamp -3599
transform 1 0 24564 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _041_
timestamp -3599
transform 1 0 27232 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _042_
timestamp -3599
transform 1 0 29256 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _043_
timestamp -3599
transform -1 0 42044 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _044_
timestamp -3599
transform -1 0 43332 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _045_
timestamp -3599
transform -1 0 44068 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _046_
timestamp -3599
transform -1 0 43608 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _047_
timestamp -3599
transform -1 0 37076 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _048_
timestamp -3599
transform -1 0 42780 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _049_
timestamp -3599
transform -1 0 44620 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _050_
timestamp -3599
transform -1 0 45632 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _051_
timestamp -3599
transform -1 0 45356 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _052_
timestamp -3599
transform -1 0 16928 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _053_
timestamp -3599
transform -1 0 15916 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _054_
timestamp -3599
transform -1 0 14352 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _055_
timestamp -3599
transform -1 0 12788 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _056_
timestamp -3599
transform 1 0 23644 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _057_
timestamp -3599
transform -1 0 22724 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _058_
timestamp -3599
transform -1 0 22080 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _059_
timestamp -3599
transform -1 0 21620 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _060_
timestamp -3599
transform -1 0 21528 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _061_
timestamp -3599
transform -1 0 21068 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _062_
timestamp -3599
transform -1 0 20240 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _063_
timestamp -3599
transform -1 0 18308 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _064_
timestamp -3599
transform -1 0 29808 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _065_
timestamp -3599
transform -1 0 28520 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _066_
timestamp -3599
transform -1 0 27324 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _067_
timestamp -3599
transform -1 0 26312 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _068_
timestamp -3599
transform -1 0 26680 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _069_
timestamp -3599
transform -1 0 26496 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _070_
timestamp -3599
transform -1 0 26036 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _071_
timestamp -3599
transform -1 0 24748 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _072_
timestamp -3599
transform -1 0 37904 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _073_
timestamp -3599
transform -1 0 36524 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _074_
timestamp -3599
transform -1 0 35604 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _075_
timestamp -3599
transform -1 0 34500 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _076_
timestamp -3599
transform -1 0 33580 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _077_
timestamp -3599
transform 1 0 32292 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _078_
timestamp -3599
transform -1 0 31740 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _079_
timestamp -3599
transform -1 0 30452 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _080_
timestamp -3599
transform -1 0 29072 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _081_
timestamp -3599
transform -1 0 29440 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _082_
timestamp -3599
transform -1 0 30084 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _083_
timestamp -3599
transform -1 0 30912 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _084_
timestamp -3599
transform -1 0 11408 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _085_
timestamp -3599
transform -1 0 11132 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _086_
timestamp -3599
transform -1 0 12236 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _087_
timestamp -3599
transform -1 0 13156 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _088_
timestamp -3599
transform -1 0 13984 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _089_
timestamp -3599
transform -1 0 14812 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _090_
timestamp -3599
transform -1 0 14720 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _091_
timestamp -3599
transform -1 0 15732 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _092_
timestamp -3599
transform -1 0 16008 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _093_
timestamp -3599
transform -1 0 15824 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _094_
timestamp -3599
transform -1 0 16560 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _095_
timestamp -3599
transform 1 0 17112 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _096_
timestamp -3599
transform 1 0 17756 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _097_
timestamp -3599
transform 1 0 18124 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _098_
timestamp -3599
transform 1 0 19412 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _099_
timestamp -3599
transform 1 0 20148 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _100_
timestamp -3599
transform -1 0 40756 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _101_
timestamp -3599
transform -1 0 39744 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _102_
timestamp -3599
transform -1 0 39928 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _103_
timestamp -3599
transform -1 0 39192 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp -3599
transform 1 0 38548 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp -3599
transform 1 0 8096 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp -3599
transform 1 0 25300 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp -3599
transform -1 0 18584 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp -3599
transform -1 0 17572 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp -3599
transform 1 0 20056 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp -3599
transform 1 0 14444 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp -3599
transform -1 0 17848 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp -3599
transform -1 0 37444 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp -3599
transform -1 0 22908 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp -3599
transform -1 0 36708 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp -3599
transform 1 0 41584 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp -3599
transform 1 0 30176 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp -3599
transform 1 0 20056 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp -3599
transform 1 0 45632 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp -3599
transform 1 0 20700 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp -3599
transform -1 0 25116 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp -3599
transform -1 0 23368 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp -3599
transform 1 0 22540 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp -3599
transform -1 0 25024 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp -3599
transform 1 0 17940 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp -3599
transform 1 0 41584 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_22
timestamp -3599
transform -1 0 2944 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_23
timestamp -3599
transform -1 0 20056 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_24
timestamp -3599
transform 1 0 20792 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_25
timestamp -3599
transform -1 0 12880 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_26
timestamp -3599
transform -1 0 11960 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_27
timestamp -3599
transform -1 0 10856 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_28
timestamp -3599
transform -1 0 15548 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_29
timestamp -3599
transform -1 0 15180 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_30
timestamp -3599
transform -1 0 20148 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_31
timestamp -3599
transform -1 0 19412 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_32
timestamp -3599
transform -1 0 16284 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_33
timestamp -3599
transform -1 0 6624 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_34
timestamp -3599
transform -1 0 15456 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_35
timestamp -3599
transform -1 0 13708 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3
timestamp 1636964856
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1636964856
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27
timestamp -3599
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1636964856
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1636964856
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53
timestamp -3599
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1636964856
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1636964856
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp -3599
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1636964856
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1636964856
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp -3599
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1636964856
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1636964856
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp -3599
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1636964856
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1636964856
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp -3599
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1636964856
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1636964856
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp -3599
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 1636964856
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_209
timestamp 1636964856
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp -3599
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_225
timestamp 1636964856
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_237
timestamp 1636964856
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp -3599
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_253
timestamp 1636964856
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_265
timestamp 1636964856
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp -3599
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_281
timestamp 1636964856
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_293
timestamp 1636964856
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp -3599
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_309
timestamp 1636964856
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_321
timestamp 1636964856
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_333
timestamp -3599
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_337
timestamp 1636964856
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_349
timestamp 1636964856
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361
timestamp -3599
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_365
timestamp 1636964856
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_377
timestamp 1636964856
transform 1 0 35788 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_389
timestamp -3599
transform 1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_393
timestamp 1636964856
transform 1 0 37260 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_405
timestamp 1636964856
transform 1 0 38364 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_417
timestamp -3599
transform 1 0 39468 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_421
timestamp 1636964856
transform 1 0 39836 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_433
timestamp 1636964856
transform 1 0 40940 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_445
timestamp -3599
transform 1 0 42044 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_449
timestamp 1636964856
transform 1 0 42412 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_461
timestamp 1636964856
transform 1 0 43516 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_473
timestamp -3599
transform 1 0 44620 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_477
timestamp -3599
transform 1 0 44988 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_483
timestamp -3599
transform 1 0 45540 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1636964856
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1636964856
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1636964856
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1636964856
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp -3599
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp -3599
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1636964856
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_69
timestamp -3599
transform 1 0 7452 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_75
timestamp -3599
transform 1 0 8004 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_86
timestamp 1636964856
transform 1 0 9016 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_98
timestamp -3599
transform 1 0 10120 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_104
timestamp -3599
transform 1 0 10672 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_109
timestamp -3599
transform 1 0 11132 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1636964856
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_133
timestamp 1636964856
transform 1 0 13340 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_145
timestamp 1636964856
transform 1 0 14444 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_157
timestamp -3599
transform 1 0 15548 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_162
timestamp -3599
transform 1 0 16008 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_1_173
timestamp -3599
transform 1 0 17020 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_179
timestamp -3599
transform 1 0 17572 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_186
timestamp -3599
transform 1 0 18216 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_190
timestamp -3599
transform 1 0 18584 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_194
timestamp 1636964856
transform 1 0 18952 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_211
timestamp -3599
transform 1 0 20516 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_218
timestamp -3599
transform 1 0 21160 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_225
timestamp -3599
transform 1 0 21804 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_229
timestamp -3599
transform 1 0 22172 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_240
timestamp 1636964856
transform 1 0 23184 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_252
timestamp -3599
transform 1 0 24288 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_260
timestamp -3599
transform 1 0 25024 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_266
timestamp 1636964856
transform 1 0 25576 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_278
timestamp -3599
transform 1 0 26680 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_281
timestamp -3599
transform 1 0 26956 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_290
timestamp 1636964856
transform 1 0 27784 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_302
timestamp -3599
transform 1 0 28888 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_309
timestamp 1636964856
transform 1 0 29532 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_321
timestamp 1636964856
transform 1 0 30636 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_333
timestamp -3599
transform 1 0 31740 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1636964856
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1636964856
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_361
timestamp 1636964856
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_373
timestamp 1636964856
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_390
timestamp -3599
transform 1 0 36984 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_398
timestamp -3599
transform 1 0 37720 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_406
timestamp -3599
transform 1 0 38456 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_411
timestamp -3599
transform 1 0 38916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_1_420
timestamp -3599
transform 1 0 39744 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_429
timestamp 1636964856
transform 1 0 40572 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_441
timestamp -3599
transform 1 0 41676 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp -3599
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_449
timestamp -3599
transform 1 0 42412 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_455
timestamp -3599
transform 1 0 42964 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_459
timestamp -3599
transform 1 0 43332 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_463
timestamp -3599
transform 1 0 43700 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_467
timestamp 1636964856
transform 1 0 44068 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_479
timestamp 1636964856
transform 1 0 45172 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_491
timestamp -3599
transform 1 0 46276 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_495
timestamp -3599
transform 1 0 46644 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1636964856
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1636964856
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp -3599
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1636964856
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1636964856
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1636964856
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1636964856
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp -3599
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp -3599
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1636964856
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1636964856
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1636964856
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1636964856
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp -3599
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp -3599
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_144
timestamp 1636964856
transform 1 0 14352 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_156
timestamp 1636964856
transform 1 0 15456 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_168
timestamp 1636964856
transform 1 0 16560 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_180
timestamp 1636964856
transform 1 0 17664 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_192
timestamp -3599
transform 1 0 18768 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_197
timestamp -3599
transform 1 0 19228 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_208
timestamp 1636964856
transform 1 0 20240 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_220
timestamp 1636964856
transform 1 0 21344 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_232
timestamp 1636964856
transform 1 0 22448 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_244
timestamp -3599
transform 1 0 23552 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_253
timestamp -3599
transform 1 0 24380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_258
timestamp -3599
transform 1 0 24840 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_264
timestamp 1636964856
transform 1 0 25392 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_276
timestamp 1636964856
transform 1 0 26496 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_288
timestamp 1636964856
transform 1 0 27600 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_300
timestamp -3599
transform 1 0 28704 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1636964856
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1636964856
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1636964856
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1636964856
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp -3599
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp -3599
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1636964856
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1636964856
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_389
timestamp 1636964856
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_401
timestamp 1636964856
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_413
timestamp -3599
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp -3599
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_421
timestamp 1636964856
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_433
timestamp 1636964856
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_445
timestamp 1636964856
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_457
timestamp 1636964856
transform 1 0 43148 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_469
timestamp -3599
transform 1 0 44252 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_475
timestamp -3599
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_477
timestamp 1636964856
transform 1 0 44988 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_489
timestamp -3599
transform 1 0 46092 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1636964856
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1636964856
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1636964856
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1636964856
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp -3599
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp -3599
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1636964856
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1636964856
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1636964856
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1636964856
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp -3599
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp -3599
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_113
timestamp -3599
transform 1 0 11500 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_121
timestamp -3599
transform 1 0 12236 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_127
timestamp 1636964856
transform 1 0 12788 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_139
timestamp 1636964856
transform 1 0 13892 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_151
timestamp -3599
transform 1 0 14996 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_157
timestamp -3599
transform 1 0 15548 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp -3599
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp -3599
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_172
timestamp -3599
transform 1 0 16928 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_180
timestamp -3599
transform 1 0 17664 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_189
timestamp 1636964856
transform 1 0 18492 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_201
timestamp 1636964856
transform 1 0 19596 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_213
timestamp -3599
transform 1 0 20700 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_221
timestamp -3599
transform 1 0 21436 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_225
timestamp -3599
transform 1 0 21804 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_3_238
timestamp 1636964856
transform 1 0 23000 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_250
timestamp 1636964856
transform 1 0 24104 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_262
timestamp 1636964856
transform 1 0 25208 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_274
timestamp -3599
transform 1 0 26312 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1636964856
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1636964856
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1636964856
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1636964856
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp -3599
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp -3599
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1636964856
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1636964856
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1636964856
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1636964856
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp -3599
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp -3599
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1636964856
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_405
timestamp 1636964856
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_417
timestamp 1636964856
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_429
timestamp 1636964856
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp -3599
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp -3599
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_449
timestamp 1636964856
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_461
timestamp 1636964856
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_473
timestamp 1636964856
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_485
timestamp -3599
transform 1 0 45724 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_493
timestamp -3599
transform 1 0 46460 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1636964856
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1636964856
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp -3599
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1636964856
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1636964856
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1636964856
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1636964856
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp -3599
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp -3599
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1636964856
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1636964856
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1636964856
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1636964856
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp -3599
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp -3599
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1636964856
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1636964856
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1636964856
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_177
timestamp -3599
transform 1 0 17388 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_183
timestamp -3599
transform 1 0 17940 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_187
timestamp -3599
transform 1 0 18308 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp -3599
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_197
timestamp -3599
transform 1 0 19228 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_205
timestamp -3599
transform 1 0 19964 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_211
timestamp -3599
transform 1 0 20516 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_217
timestamp -3599
transform 1 0 21068 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_222
timestamp 1636964856
transform 1 0 21528 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_234
timestamp -3599
transform 1 0 22632 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp -3599
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp -3599
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_253
timestamp -3599
transform 1 0 24380 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_257
timestamp -3599
transform 1 0 24748 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_263
timestamp 1636964856
transform 1 0 25300 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_275
timestamp 1636964856
transform 1 0 26404 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_287
timestamp 1636964856
transform 1 0 27508 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_299
timestamp -3599
transform 1 0 28612 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp -3599
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1636964856
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1636964856
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1636964856
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1636964856
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp -3599
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp -3599
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1636964856
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1636964856
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1636964856
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_401
timestamp 1636964856
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp -3599
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp -3599
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1636964856
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 1636964856
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_445
timestamp 1636964856
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_457
timestamp 1636964856
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp -3599
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp -3599
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_477
timestamp 1636964856
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_489
timestamp -3599
transform 1 0 46092 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1636964856
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1636964856
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1636964856
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1636964856
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp -3599
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp -3599
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1636964856
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1636964856
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_81
timestamp -3599
transform 1 0 8556 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_5_91
timestamp 1636964856
transform 1 0 9476 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_103
timestamp -3599
transform 1 0 10580 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp -3599
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1636964856
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1636964856
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1636964856
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1636964856
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp -3599
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp -3599
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1636964856
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1636964856
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1636964856
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1636964856
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_217
timestamp -3599
transform 1 0 21068 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp -3599
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_228
timestamp 1636964856
transform 1 0 22080 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_240
timestamp -3599
transform 1 0 23184 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_244
timestamp -3599
transform 1 0 23552 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_248
timestamp 1636964856
transform 1 0 23920 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_260
timestamp 1636964856
transform 1 0 25024 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_272
timestamp -3599
transform 1 0 26128 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1636964856
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1636964856
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1636964856
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_317
timestamp 1636964856
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp -3599
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp -3599
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1636964856
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1636964856
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1636964856
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1636964856
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp -3599
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp -3599
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_393
timestamp -3599
transform 1 0 37260 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_400
timestamp 1636964856
transform 1 0 37904 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_412
timestamp 1636964856
transform 1 0 39008 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_424
timestamp 1636964856
transform 1 0 40112 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_436
timestamp 1636964856
transform 1 0 41216 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_449
timestamp 1636964856
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_461
timestamp 1636964856
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_473
timestamp 1636964856
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_485
timestamp -3599
transform 1 0 45724 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_493
timestamp -3599
transform 1 0 46460 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1636964856
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1636964856
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp -3599
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1636964856
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1636964856
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1636964856
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1636964856
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp -3599
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp -3599
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1636964856
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1636964856
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1636964856
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1636964856
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp -3599
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp -3599
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_141
timestamp -3599
transform 1 0 14076 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_151
timestamp 1636964856
transform 1 0 14996 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_163
timestamp 1636964856
transform 1 0 16100 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_175
timestamp -3599
transform 1 0 17204 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_183
timestamp 1636964856
transform 1 0 17940 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp -3599
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1636964856
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1636964856
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_221
timestamp -3599
transform 1 0 21436 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_229
timestamp -3599
transform 1 0 22172 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_235
timestamp 1636964856
transform 1 0 22724 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_247
timestamp -3599
transform 1 0 23828 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp -3599
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1636964856
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1636964856
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1636964856
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1636964856
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_304
timestamp -3599
transform 1 0 29072 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_309
timestamp -3599
transform 1 0 29532 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_315
timestamp -3599
transform 1 0 30084 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_319
timestamp -3599
transform 1 0 30452 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_327
timestamp -3599
transform 1 0 31188 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1636964856
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1636964856
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp -3599
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp -3599
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1636964856
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1636964856
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1636964856
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_401
timestamp -3599
transform 1 0 37996 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_409
timestamp -3599
transform 1 0 38732 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_414
timestamp -3599
transform 1 0 39192 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1636964856
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 1636964856
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_445
timestamp 1636964856
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_457
timestamp 1636964856
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp -3599
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp -3599
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_477
timestamp 1636964856
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_489
timestamp -3599
transform 1 0 46092 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1636964856
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1636964856
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1636964856
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1636964856
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp -3599
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp -3599
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1636964856
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1636964856
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1636964856
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1636964856
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp -3599
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp -3599
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1636964856
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1636964856
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1636964856
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1636964856
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp -3599
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp -3599
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1636964856
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1636964856
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1636964856
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1636964856
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp -3599
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp -3599
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1636964856
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1636964856
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_249
timestamp -3599
transform 1 0 24012 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_253
timestamp -3599
transform 1 0 24380 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_257
timestamp -3599
transform 1 0 24748 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_271
timestamp -3599
transform 1 0 26036 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_276
timestamp -3599
transform 1 0 26496 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1636964856
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1636964856
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1636964856
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1636964856
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp -3599
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp -3599
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_337
timestamp -3599
transform 1 0 32108 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_345
timestamp -3599
transform 1 0 32844 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1636964856
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1636964856
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_373
timestamp -3599
transform 1 0 35420 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp -3599
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp -3599
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1636964856
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_405
timestamp 1636964856
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_417
timestamp -3599
transform 1 0 39468 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_422
timestamp 1636964856
transform 1 0 39928 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_434
timestamp 1636964856
transform 1 0 41032 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_446
timestamp -3599
transform 1 0 42136 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_449
timestamp 1636964856
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_461
timestamp 1636964856
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_473
timestamp 1636964856
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_485
timestamp -3599
transform 1 0 45724 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_491
timestamp -3599
transform 1 0 46276 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1636964856
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1636964856
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp -3599
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1636964856
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1636964856
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1636964856
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1636964856
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp -3599
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp -3599
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1636964856
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1636964856
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1636964856
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1636964856
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp -3599
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp -3599
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1636964856
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_153
timestamp -3599
transform 1 0 15180 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_160
timestamp -3599
transform 1 0 15824 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_168
timestamp 1636964856
transform 1 0 16560 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_180
timestamp 1636964856
transform 1 0 17664 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_192
timestamp -3599
transform 1 0 18768 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1636964856
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1636964856
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1636964856
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_233
timestamp -3599
transform 1 0 22540 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_241
timestamp -3599
transform 1 0 23276 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_246
timestamp -3599
transform 1 0 23736 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1636964856
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1636964856
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1636964856
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1636964856
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_301
timestamp -3599
transform 1 0 28796 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1636964856
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1636964856
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_333
timestamp -3599
transform 1 0 31740 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_342
timestamp 1636964856
transform 1 0 32568 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_354
timestamp -3599
transform 1 0 33672 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_362
timestamp -3599
transform 1 0 34408 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_365
timestamp -3599
transform 1 0 34684 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_371
timestamp -3599
transform 1 0 35236 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_375
timestamp 1636964856
transform 1 0 35604 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_387
timestamp 1636964856
transform 1 0 36708 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_399
timestamp 1636964856
transform 1 0 37812 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_411
timestamp -3599
transform 1 0 38916 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp -3599
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_421
timestamp 1636964856
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_433
timestamp 1636964856
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_445
timestamp 1636964856
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_457
timestamp 1636964856
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp -3599
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp -3599
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_477
timestamp -3599
transform 1 0 44988 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_483
timestamp -3599
transform 1 0 45540 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1636964856
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1636964856
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1636964856
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1636964856
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp -3599
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp -3599
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1636964856
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_69
timestamp -3599
transform 1 0 7452 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_75
timestamp 1636964856
transform 1 0 8004 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_87
timestamp 1636964856
transform 1 0 9108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_99
timestamp 1636964856
transform 1 0 10212 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp -3599
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1636964856
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1636964856
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_137
timestamp -3599
transform 1 0 13708 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_148
timestamp -3599
transform 1 0 14720 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_153
timestamp -3599
transform 1 0 15180 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_162
timestamp -3599
transform 1 0 16008 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_169
timestamp -3599
transform 1 0 16652 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_173
timestamp -3599
transform 1 0 17020 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_177
timestamp 1636964856
transform 1 0 17388 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_189
timestamp 1636964856
transform 1 0 18492 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_201
timestamp 1636964856
transform 1 0 19596 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_213
timestamp -3599
transform 1 0 20700 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_221
timestamp -3599
transform 1 0 21436 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_228
timestamp 1636964856
transform 1 0 22080 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_240
timestamp 1636964856
transform 1 0 23184 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_252
timestamp 1636964856
transform 1 0 24288 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_264
timestamp -3599
transform 1 0 25392 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_272
timestamp -3599
transform 1 0 26128 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_278
timestamp -3599
transform 1 0 26680 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1636964856
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1636964856
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1636964856
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_317
timestamp 1636964856
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp -3599
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp -3599
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1636964856
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_349
timestamp -3599
transform 1 0 33212 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_353
timestamp 1636964856
transform 1 0 33580 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_365
timestamp 1636964856
transform 1 0 34684 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_377
timestamp 1636964856
transform 1 0 35788 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_389
timestamp -3599
transform 1 0 36892 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_393
timestamp 1636964856
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_405
timestamp 1636964856
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_417
timestamp 1636964856
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_429
timestamp -3599
transform 1 0 40572 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_437
timestamp -3599
transform 1 0 41308 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_445
timestamp -3599
transform 1 0 42044 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_449
timestamp -3599
transform 1 0 42412 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_453
timestamp -3599
transform 1 0 42780 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_9_462
timestamp -3599
transform 1 0 43608 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_473
timestamp -3599
transform 1 0 44620 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_477
timestamp -3599
transform 1 0 44988 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_3
timestamp -3599
transform 1 0 1380 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_8
timestamp -3599
transform 1 0 1840 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1636964856
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp -3599
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_29
timestamp -3599
transform 1 0 3772 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_34
timestamp -3599
transform 1 0 4232 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_42
timestamp -3599
transform 1 0 4968 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_47
timestamp -3599
transform 1 0 5428 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_55
timestamp -3599
transform 1 0 6164 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_62
timestamp 1636964856
transform 1 0 6808 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_74
timestamp -3599
transform 1 0 7912 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_82
timestamp -3599
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_85
timestamp -3599
transform 1 0 8924 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_90
timestamp 1636964856
transform 1 0 9384 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_102
timestamp -3599
transform 1 0 10488 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_112
timestamp -3599
transform 1 0 11408 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_125
timestamp -3599
transform 1 0 12604 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_131
timestamp -3599
transform 1 0 13156 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_141
timestamp -3599
transform 1 0 14076 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_149
timestamp 1636964856
transform 1 0 14812 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_161
timestamp -3599
transform 1 0 15916 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_169
timestamp -3599
transform 1 0 16652 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_178
timestamp -3599
transform 1 0 17480 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_184
timestamp -3599
transform 1 0 18032 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_194
timestamp -3599
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_202
timestamp -3599
transform 1 0 19688 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_210
timestamp 1636964856
transform 1 0 20424 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_225
timestamp 1636964856
transform 1 0 21804 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_237
timestamp 1636964856
transform 1 0 22908 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_249
timestamp -3599
transform 1 0 24012 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1636964856
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_265
timestamp -3599
transform 1 0 25484 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_10_274
timestamp -3599
transform 1 0 26312 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_285
timestamp -3599
transform 1 0 27324 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_293
timestamp -3599
transform 1 0 28060 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_298
timestamp -3599
transform 1 0 28520 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_306
timestamp -3599
transform 1 0 29256 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_315
timestamp -3599
transform 1 0 30084 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_324
timestamp 1636964856
transform 1 0 30912 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_336
timestamp 1636964856
transform 1 0 32016 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_348
timestamp 1636964856
transform 1 0 33120 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp -3599
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1636964856
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_377
timestamp -3599
transform 1 0 35788 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_385
timestamp -3599
transform 1 0 36524 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_391
timestamp 1636964856
transform 1 0 37076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_403
timestamp 1636964856
transform 1 0 38180 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_415
timestamp -3599
transform 1 0 39284 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_421
timestamp -3599
transform 1 0 39836 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_427
timestamp -3599
transform 1 0 40388 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_431
timestamp -3599
transform 1 0 40756 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_439
timestamp -3599
transform 1 0 41492 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_445
timestamp 1636964856
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_457
timestamp 1636964856
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp -3599
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp -3599
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_477
timestamp -3599
transform 1 0 44988 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_502
timestamp -3599
transform 1 0 47288 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_3
timestamp -3599
transform 1 0 1380 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_29
timestamp -3599
transform 1 0 3772 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_57
timestamp -3599
transform 1 0 6348 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_85
timestamp -3599
transform 1 0 8924 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_113
timestamp -3599
transform 1 0 11500 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_141
timestamp -3599
transform 1 0 14076 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_169
timestamp -3599
transform 1 0 16652 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_197
timestamp -3599
transform 1 0 19228 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_216
timestamp -3599
transform 1 0 20976 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1636964856
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1636964856
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_249
timestamp -3599
transform 1 0 24012 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_253
timestamp 1636964856
transform 1 0 24380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_265
timestamp 1636964856
transform 1 0 25484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_277
timestamp -3599
transform 1 0 26588 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1636964856
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_293
timestamp 1636964856
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_305
timestamp -3599
transform 1 0 29164 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_309
timestamp 1636964856
transform 1 0 29532 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_321
timestamp 1636964856
transform 1 0 30636 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_333
timestamp -3599
transform 1 0 31740 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1636964856
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_349
timestamp 1636964856
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_361
timestamp -3599
transform 1 0 34316 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_365
timestamp 1636964856
transform 1 0 34684 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_377
timestamp 1636964856
transform 1 0 35788 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_389
timestamp -3599
transform 1 0 36892 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_393
timestamp 1636964856
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_405
timestamp 1636964856
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_417
timestamp -3599
transform 1 0 39468 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_421
timestamp -3599
transform 1 0 39836 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_425
timestamp -3599
transform 1 0 40204 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_446
timestamp -3599
transform 1 0 42136 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_473
timestamp -3599
transform 1 0 44620 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_501
timestamp -3599
transform 1 0 47196 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output1
timestamp -3599
transform 1 0 46368 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output2
timestamp -3599
transform 1 0 47104 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output3
timestamp -3599
transform 1 0 46828 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output4
timestamp -3599
transform 1 0 47196 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output5
timestamp -3599
transform 1 0 46736 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output6
timestamp -3599
transform 1 0 47104 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output7
timestamp -3599
transform 1 0 46828 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output8
timestamp -3599
transform 1 0 46368 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output9
timestamp -3599
transform 1 0 47196 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp -3599
transform 1 0 46092 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp -3599
transform 1 0 46736 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp -3599
transform 1 0 46000 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp -3599
transform 1 0 46460 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp -3599
transform 1 0 47196 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output15
timestamp -3599
transform 1 0 46736 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output16
timestamp -3599
transform 1 0 47104 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output17
timestamp -3599
transform 1 0 45816 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output18
timestamp -3599
transform 1 0 46368 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output19
timestamp -3599
transform 1 0 46828 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output20
timestamp -3599
transform 1 0 46000 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output21
timestamp -3599
transform 1 0 45448 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output22
timestamp -3599
transform 1 0 45632 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output23
timestamp -3599
transform 1 0 45632 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output24
timestamp -3599
transform 1 0 45080 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output25
timestamp -3599
transform 1 0 47104 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output26
timestamp -3599
transform 1 0 46736 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output27
timestamp -3599
transform 1 0 47104 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output28
timestamp -3599
transform 1 0 46736 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output29
timestamp -3599
transform 1 0 47104 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output30
timestamp -3599
transform 1 0 46828 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output31
timestamp -3599
transform 1 0 47196 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output32
timestamp -3599
transform 1 0 46736 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output33
timestamp -3599
transform 1 0 40296 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output34
timestamp -3599
transform 1 0 44252 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output35
timestamp -3599
transform 1 0 44988 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output36
timestamp -3599
transform 1 0 45356 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output37
timestamp -3599
transform 1 0 45724 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output38
timestamp -3599
transform 1 0 46092 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output39
timestamp -3599
transform 1 0 46460 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output40
timestamp -3599
transform 1 0 46828 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output41
timestamp -3599
transform 1 0 46552 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output42
timestamp -3599
transform 1 0 46920 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output43
timestamp -3599
transform 1 0 46184 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output44
timestamp -3599
transform 1 0 40664 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output45
timestamp -3599
transform 1 0 41032 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output46
timestamp -3599
transform 1 0 41400 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output47
timestamp -3599
transform 1 0 41768 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output48
timestamp -3599
transform 1 0 42412 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output49
timestamp -3599
transform 1 0 42780 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output50
timestamp -3599
transform 1 0 43148 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output51
timestamp -3599
transform 1 0 43516 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output52
timestamp -3599
transform 1 0 43884 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output53
timestamp -3599
transform -1 0 1840 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output54
timestamp -3599
transform -1 0 2024 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output55
timestamp -3599
transform -1 0 2392 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output56
timestamp -3599
transform -1 0 2760 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output57
timestamp -3599
transform -1 0 3312 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output58
timestamp -3599
transform -1 0 3680 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output59
timestamp -3599
transform -1 0 4232 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output60
timestamp -3599
transform -1 0 4416 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output61
timestamp -3599
transform -1 0 4784 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp -3599
transform -1 0 5152 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output63
timestamp -3599
transform -1 0 5520 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp -3599
transform -1 0 5888 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp -3599
transform -1 0 6256 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp -3599
transform -1 0 6808 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp -3599
transform -1 0 6992 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp -3599
transform -1 0 7360 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp -3599
transform -1 0 7728 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp -3599
transform -1 0 8096 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp -3599
transform -1 0 8464 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp -3599
transform -1 0 8832 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp -3599
transform -1 0 9384 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp -3599
transform -1 0 12880 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp -3599
transform -1 0 13248 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp -3599
transform 1 0 13248 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp -3599
transform 1 0 13616 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp -3599
transform 1 0 14168 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp -3599
transform 1 0 14352 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp -3599
transform -1 0 9568 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp -3599
transform -1 0 9936 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp -3599
transform -1 0 10304 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp -3599
transform -1 0 10672 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp -3599
transform -1 0 11040 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp -3599
transform -1 0 11408 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp -3599
transform -1 0 12604 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp -3599
transform -1 0 12144 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp -3599
transform -1 0 12512 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp -3599
transform 1 0 14720 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp -3599
transform -1 0 18400 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp -3599
transform -1 0 18768 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp -3599
transform -1 0 19136 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp -3599
transform -1 0 19872 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp -3599
transform -1 0 20424 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp -3599
transform -1 0 20792 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp -3599
transform 1 0 15088 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp -3599
transform 1 0 15456 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp -3599
transform 1 0 15824 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp -3599
transform 1 0 16192 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output100
timestamp -3599
transform 1 0 16744 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output101
timestamp -3599
transform 1 0 17112 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp -3599
transform 1 0 16928 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output103
timestamp -3599
transform -1 0 17664 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output104
timestamp -3599
transform -1 0 18032 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  output105
timestamp -3599
transform -1 0 40204 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_12
timestamp -3599
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp -3599
transform -1 0 47840 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_13
timestamp -3599
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp -3599
transform -1 0 47840 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_14
timestamp -3599
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp -3599
transform -1 0 47840 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_15
timestamp -3599
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp -3599
transform -1 0 47840 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_16
timestamp -3599
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp -3599
transform -1 0 47840 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_17
timestamp -3599
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp -3599
transform -1 0 47840 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_18
timestamp -3599
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp -3599
transform -1 0 47840 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_19
timestamp -3599
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp -3599
transform -1 0 47840 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_20
timestamp -3599
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp -3599
transform -1 0 47840 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_21
timestamp -3599
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp -3599
transform -1 0 47840 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_22
timestamp -3599
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp -3599
transform -1 0 47840 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_23
timestamp -3599
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp -3599
transform -1 0 47840 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_24
timestamp -3599
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_25
timestamp -3599
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_26
timestamp -3599
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_27
timestamp -3599
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_28
timestamp -3599
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_29
timestamp -3599
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_30
timestamp -3599
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_31
timestamp -3599
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_32
timestamp -3599
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_33
timestamp -3599
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_34
timestamp -3599
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_35
timestamp -3599
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_36
timestamp -3599
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_37
timestamp -3599
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_38
timestamp -3599
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_39
timestamp -3599
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_40
timestamp -3599
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_41
timestamp -3599
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_42
timestamp -3599
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_43
timestamp -3599
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_44
timestamp -3599
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_45
timestamp -3599
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_46
timestamp -3599
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_47
timestamp -3599
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_48
timestamp -3599
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_49
timestamp -3599
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_50
timestamp -3599
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_51
timestamp -3599
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_52
timestamp -3599
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_53
timestamp -3599
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_54
timestamp -3599
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_55
timestamp -3599
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_56
timestamp -3599
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_57
timestamp -3599
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_58
timestamp -3599
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_59
timestamp -3599
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_60
timestamp -3599
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_61
timestamp -3599
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_62
timestamp -3599
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_63
timestamp -3599
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_64
timestamp -3599
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_65
timestamp -3599
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_66
timestamp -3599
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_67
timestamp -3599
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_68
timestamp -3599
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_69
timestamp -3599
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_70
timestamp -3599
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_71
timestamp -3599
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_72
timestamp -3599
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_73
timestamp -3599
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_74
timestamp -3599
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_75
timestamp -3599
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_76
timestamp -3599
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_77
timestamp -3599
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_78
timestamp -3599
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_79
timestamp -3599
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_80
timestamp -3599
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_81
timestamp -3599
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_82
timestamp -3599
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_83
timestamp -3599
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_84
timestamp -3599
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_85
timestamp -3599
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_86
timestamp -3599
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_87
timestamp -3599
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_88
timestamp -3599
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_89
timestamp -3599
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_90
timestamp -3599
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_91
timestamp -3599
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_92
timestamp -3599
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_93
timestamp -3599
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_94
timestamp -3599
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_95
timestamp -3599
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_96
timestamp -3599
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_97
timestamp -3599
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_98
timestamp -3599
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_99
timestamp -3599
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_100
timestamp -3599
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_101
timestamp -3599
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_102
timestamp -3599
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_103
timestamp -3599
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_104
timestamp -3599
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_105
timestamp -3599
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_106
timestamp -3599
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_107
timestamp -3599
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_108
timestamp -3599
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_109
timestamp -3599
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_110
timestamp -3599
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_111
timestamp -3599
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_112
timestamp -3599
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_113
timestamp -3599
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_114
timestamp -3599
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_115
timestamp -3599
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_116
timestamp -3599
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_117
timestamp -3599
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_118
timestamp -3599
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_119
timestamp -3599
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_120
timestamp -3599
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_121
timestamp -3599
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_122
timestamp -3599
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_123
timestamp -3599
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_124
timestamp -3599
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_125
timestamp -3599
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_126
timestamp -3599
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_127
timestamp -3599
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_128
timestamp -3599
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_129
timestamp -3599
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_130
timestamp -3599
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_131
timestamp -3599
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_132
timestamp -3599
transform 1 0 3680 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_133
timestamp -3599
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_134
timestamp -3599
transform 1 0 8832 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_135
timestamp -3599
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_136
timestamp -3599
transform 1 0 13984 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_137
timestamp -3599
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_138
timestamp -3599
transform 1 0 19136 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_139
timestamp -3599
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_140
timestamp -3599
transform 1 0 24288 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_141
timestamp -3599
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_142
timestamp -3599
transform 1 0 29440 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_143
timestamp -3599
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_144
timestamp -3599
transform 1 0 34592 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_145
timestamp -3599
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_146
timestamp -3599
transform 1 0 39744 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_147
timestamp -3599
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_148
timestamp -3599
transform 1 0 44896 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_149
timestamp -3599
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
<< labels >>
flabel metal3 s 0 1368 120 1488 0 FreeSans 480 0 0 0 FrameData[0]
port 0 nsew signal input
flabel metal3 s 0 4088 120 4208 0 FreeSans 480 0 0 0 FrameData[10]
port 1 nsew signal input
flabel metal3 s 0 4360 120 4480 0 FreeSans 480 0 0 0 FrameData[11]
port 2 nsew signal input
flabel metal3 s 0 4632 120 4752 0 FreeSans 480 0 0 0 FrameData[12]
port 3 nsew signal input
flabel metal3 s 0 4904 120 5024 0 FreeSans 480 0 0 0 FrameData[13]
port 4 nsew signal input
flabel metal3 s 0 5176 120 5296 0 FreeSans 480 0 0 0 FrameData[14]
port 5 nsew signal input
flabel metal3 s 0 5448 120 5568 0 FreeSans 480 0 0 0 FrameData[15]
port 6 nsew signal input
flabel metal3 s 0 5720 120 5840 0 FreeSans 480 0 0 0 FrameData[16]
port 7 nsew signal input
flabel metal3 s 0 5992 120 6112 0 FreeSans 480 0 0 0 FrameData[17]
port 8 nsew signal input
flabel metal3 s 0 6264 120 6384 0 FreeSans 480 0 0 0 FrameData[18]
port 9 nsew signal input
flabel metal3 s 0 6536 120 6656 0 FreeSans 480 0 0 0 FrameData[19]
port 10 nsew signal input
flabel metal3 s 0 1640 120 1760 0 FreeSans 480 0 0 0 FrameData[1]
port 11 nsew signal input
flabel metal3 s 0 6808 120 6928 0 FreeSans 480 0 0 0 FrameData[20]
port 12 nsew signal input
flabel metal3 s 0 7080 120 7200 0 FreeSans 480 0 0 0 FrameData[21]
port 13 nsew signal input
flabel metal3 s 0 7352 120 7472 0 FreeSans 480 0 0 0 FrameData[22]
port 14 nsew signal input
flabel metal3 s 0 7624 120 7744 0 FreeSans 480 0 0 0 FrameData[23]
port 15 nsew signal input
flabel metal3 s 0 7896 120 8016 0 FreeSans 480 0 0 0 FrameData[24]
port 16 nsew signal input
flabel metal3 s 0 8168 120 8288 0 FreeSans 480 0 0 0 FrameData[25]
port 17 nsew signal input
flabel metal3 s 0 8440 120 8560 0 FreeSans 480 0 0 0 FrameData[26]
port 18 nsew signal input
flabel metal3 s 0 8712 120 8832 0 FreeSans 480 0 0 0 FrameData[27]
port 19 nsew signal input
flabel metal3 s 0 8984 120 9104 0 FreeSans 480 0 0 0 FrameData[28]
port 20 nsew signal input
flabel metal3 s 0 9256 120 9376 0 FreeSans 480 0 0 0 FrameData[29]
port 21 nsew signal input
flabel metal3 s 0 1912 120 2032 0 FreeSans 480 0 0 0 FrameData[2]
port 22 nsew signal input
flabel metal3 s 0 9528 120 9648 0 FreeSans 480 0 0 0 FrameData[30]
port 23 nsew signal input
flabel metal3 s 0 9800 120 9920 0 FreeSans 480 0 0 0 FrameData[31]
port 24 nsew signal input
flabel metal3 s 0 2184 120 2304 0 FreeSans 480 0 0 0 FrameData[3]
port 25 nsew signal input
flabel metal3 s 0 2456 120 2576 0 FreeSans 480 0 0 0 FrameData[4]
port 26 nsew signal input
flabel metal3 s 0 2728 120 2848 0 FreeSans 480 0 0 0 FrameData[5]
port 27 nsew signal input
flabel metal3 s 0 3000 120 3120 0 FreeSans 480 0 0 0 FrameData[6]
port 28 nsew signal input
flabel metal3 s 0 3272 120 3392 0 FreeSans 480 0 0 0 FrameData[7]
port 29 nsew signal input
flabel metal3 s 0 3544 120 3664 0 FreeSans 480 0 0 0 FrameData[8]
port 30 nsew signal input
flabel metal3 s 0 3816 120 3936 0 FreeSans 480 0 0 0 FrameData[9]
port 31 nsew signal input
flabel metal3 s 48880 1368 49000 1488 0 FreeSans 480 0 0 0 FrameData_O[0]
port 32 nsew signal output
flabel metal3 s 48880 4088 49000 4208 0 FreeSans 480 0 0 0 FrameData_O[10]
port 33 nsew signal output
flabel metal3 s 48880 4360 49000 4480 0 FreeSans 480 0 0 0 FrameData_O[11]
port 34 nsew signal output
flabel metal3 s 48880 4632 49000 4752 0 FreeSans 480 0 0 0 FrameData_O[12]
port 35 nsew signal output
flabel metal3 s 48880 4904 49000 5024 0 FreeSans 480 0 0 0 FrameData_O[13]
port 36 nsew signal output
flabel metal3 s 48880 5176 49000 5296 0 FreeSans 480 0 0 0 FrameData_O[14]
port 37 nsew signal output
flabel metal3 s 48880 5448 49000 5568 0 FreeSans 480 0 0 0 FrameData_O[15]
port 38 nsew signal output
flabel metal3 s 48880 5720 49000 5840 0 FreeSans 480 0 0 0 FrameData_O[16]
port 39 nsew signal output
flabel metal3 s 48880 5992 49000 6112 0 FreeSans 480 0 0 0 FrameData_O[17]
port 40 nsew signal output
flabel metal3 s 48880 6264 49000 6384 0 FreeSans 480 0 0 0 FrameData_O[18]
port 41 nsew signal output
flabel metal3 s 48880 6536 49000 6656 0 FreeSans 480 0 0 0 FrameData_O[19]
port 42 nsew signal output
flabel metal3 s 48880 1640 49000 1760 0 FreeSans 480 0 0 0 FrameData_O[1]
port 43 nsew signal output
flabel metal3 s 48880 6808 49000 6928 0 FreeSans 480 0 0 0 FrameData_O[20]
port 44 nsew signal output
flabel metal3 s 48880 7080 49000 7200 0 FreeSans 480 0 0 0 FrameData_O[21]
port 45 nsew signal output
flabel metal3 s 48880 7352 49000 7472 0 FreeSans 480 0 0 0 FrameData_O[22]
port 46 nsew signal output
flabel metal3 s 48880 7624 49000 7744 0 FreeSans 480 0 0 0 FrameData_O[23]
port 47 nsew signal output
flabel metal3 s 48880 7896 49000 8016 0 FreeSans 480 0 0 0 FrameData_O[24]
port 48 nsew signal output
flabel metal3 s 48880 8168 49000 8288 0 FreeSans 480 0 0 0 FrameData_O[25]
port 49 nsew signal output
flabel metal3 s 48880 8440 49000 8560 0 FreeSans 480 0 0 0 FrameData_O[26]
port 50 nsew signal output
flabel metal3 s 48880 8712 49000 8832 0 FreeSans 480 0 0 0 FrameData_O[27]
port 51 nsew signal output
flabel metal3 s 48880 8984 49000 9104 0 FreeSans 480 0 0 0 FrameData_O[28]
port 52 nsew signal output
flabel metal3 s 48880 9256 49000 9376 0 FreeSans 480 0 0 0 FrameData_O[29]
port 53 nsew signal output
flabel metal3 s 48880 1912 49000 2032 0 FreeSans 480 0 0 0 FrameData_O[2]
port 54 nsew signal output
flabel metal3 s 48880 9528 49000 9648 0 FreeSans 480 0 0 0 FrameData_O[30]
port 55 nsew signal output
flabel metal3 s 48880 9800 49000 9920 0 FreeSans 480 0 0 0 FrameData_O[31]
port 56 nsew signal output
flabel metal3 s 48880 2184 49000 2304 0 FreeSans 480 0 0 0 FrameData_O[3]
port 57 nsew signal output
flabel metal3 s 48880 2456 49000 2576 0 FreeSans 480 0 0 0 FrameData_O[4]
port 58 nsew signal output
flabel metal3 s 48880 2728 49000 2848 0 FreeSans 480 0 0 0 FrameData_O[5]
port 59 nsew signal output
flabel metal3 s 48880 3000 49000 3120 0 FreeSans 480 0 0 0 FrameData_O[6]
port 60 nsew signal output
flabel metal3 s 48880 3272 49000 3392 0 FreeSans 480 0 0 0 FrameData_O[7]
port 61 nsew signal output
flabel metal3 s 48880 3544 49000 3664 0 FreeSans 480 0 0 0 FrameData_O[8]
port 62 nsew signal output
flabel metal3 s 48880 3816 49000 3936 0 FreeSans 480 0 0 0 FrameData_O[9]
port 63 nsew signal output
flabel metal2 s 3698 0 3754 56 0 FreeSans 224 0 0 0 FrameStrobe[0]
port 64 nsew signal input
flabel metal2 s 26698 0 26754 56 0 FreeSans 224 0 0 0 FrameStrobe[10]
port 65 nsew signal input
flabel metal2 s 28998 0 29054 56 0 FreeSans 224 0 0 0 FrameStrobe[11]
port 66 nsew signal input
flabel metal2 s 31298 0 31354 56 0 FreeSans 224 0 0 0 FrameStrobe[12]
port 67 nsew signal input
flabel metal2 s 33598 0 33654 56 0 FreeSans 224 0 0 0 FrameStrobe[13]
port 68 nsew signal input
flabel metal2 s 35898 0 35954 56 0 FreeSans 224 0 0 0 FrameStrobe[14]
port 69 nsew signal input
flabel metal2 s 38198 0 38254 56 0 FreeSans 224 0 0 0 FrameStrobe[15]
port 70 nsew signal input
flabel metal2 s 40498 0 40554 56 0 FreeSans 224 0 0 0 FrameStrobe[16]
port 71 nsew signal input
flabel metal2 s 42798 0 42854 56 0 FreeSans 224 0 0 0 FrameStrobe[17]
port 72 nsew signal input
flabel metal2 s 45098 0 45154 56 0 FreeSans 224 0 0 0 FrameStrobe[18]
port 73 nsew signal input
flabel metal2 s 47398 0 47454 56 0 FreeSans 224 0 0 0 FrameStrobe[19]
port 74 nsew signal input
flabel metal2 s 5998 0 6054 56 0 FreeSans 224 0 0 0 FrameStrobe[1]
port 75 nsew signal input
flabel metal2 s 8298 0 8354 56 0 FreeSans 224 0 0 0 FrameStrobe[2]
port 76 nsew signal input
flabel metal2 s 10598 0 10654 56 0 FreeSans 224 0 0 0 FrameStrobe[3]
port 77 nsew signal input
flabel metal2 s 12898 0 12954 56 0 FreeSans 224 0 0 0 FrameStrobe[4]
port 78 nsew signal input
flabel metal2 s 15198 0 15254 56 0 FreeSans 224 0 0 0 FrameStrobe[5]
port 79 nsew signal input
flabel metal2 s 17498 0 17554 56 0 FreeSans 224 0 0 0 FrameStrobe[6]
port 80 nsew signal input
flabel metal2 s 19798 0 19854 56 0 FreeSans 224 0 0 0 FrameStrobe[7]
port 81 nsew signal input
flabel metal2 s 22098 0 22154 56 0 FreeSans 224 0 0 0 FrameStrobe[8]
port 82 nsew signal input
flabel metal2 s 24398 0 24454 56 0 FreeSans 224 0 0 0 FrameStrobe[9]
port 83 nsew signal input
flabel metal2 s 40222 11194 40278 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[0]
port 84 nsew signal output
flabel metal2 s 43902 11194 43958 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[10]
port 85 nsew signal output
flabel metal2 s 44270 11194 44326 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[11]
port 86 nsew signal output
flabel metal2 s 44638 11194 44694 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[12]
port 87 nsew signal output
flabel metal2 s 45006 11194 45062 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[13]
port 88 nsew signal output
flabel metal2 s 45374 11194 45430 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[14]
port 89 nsew signal output
flabel metal2 s 45742 11194 45798 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[15]
port 90 nsew signal output
flabel metal2 s 46110 11194 46166 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[16]
port 91 nsew signal output
flabel metal2 s 46478 11194 46534 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[17]
port 92 nsew signal output
flabel metal2 s 46846 11194 46902 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[18]
port 93 nsew signal output
flabel metal2 s 47214 11194 47270 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[19]
port 94 nsew signal output
flabel metal2 s 40590 11194 40646 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[1]
port 95 nsew signal output
flabel metal2 s 40958 11194 41014 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[2]
port 96 nsew signal output
flabel metal2 s 41326 11194 41382 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[3]
port 97 nsew signal output
flabel metal2 s 41694 11194 41750 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[4]
port 98 nsew signal output
flabel metal2 s 42062 11194 42118 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[5]
port 99 nsew signal output
flabel metal2 s 42430 11194 42486 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[6]
port 100 nsew signal output
flabel metal2 s 42798 11194 42854 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[7]
port 101 nsew signal output
flabel metal2 s 43166 11194 43222 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[8]
port 102 nsew signal output
flabel metal2 s 43534 11194 43590 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[9]
port 103 nsew signal output
flabel metal2 s 1582 11194 1638 11250 0 FreeSans 224 0 0 0 N1BEG[0]
port 104 nsew signal output
flabel metal2 s 1950 11194 2006 11250 0 FreeSans 224 0 0 0 N1BEG[1]
port 105 nsew signal output
flabel metal2 s 2318 11194 2374 11250 0 FreeSans 224 0 0 0 N1BEG[2]
port 106 nsew signal output
flabel metal2 s 2686 11194 2742 11250 0 FreeSans 224 0 0 0 N1BEG[3]
port 107 nsew signal output
flabel metal2 s 3054 11194 3110 11250 0 FreeSans 224 0 0 0 N2BEG[0]
port 108 nsew signal output
flabel metal2 s 3422 11194 3478 11250 0 FreeSans 224 0 0 0 N2BEG[1]
port 109 nsew signal output
flabel metal2 s 3790 11194 3846 11250 0 FreeSans 224 0 0 0 N2BEG[2]
port 110 nsew signal output
flabel metal2 s 4158 11194 4214 11250 0 FreeSans 224 0 0 0 N2BEG[3]
port 111 nsew signal output
flabel metal2 s 4526 11194 4582 11250 0 FreeSans 224 0 0 0 N2BEG[4]
port 112 nsew signal output
flabel metal2 s 4894 11194 4950 11250 0 FreeSans 224 0 0 0 N2BEG[5]
port 113 nsew signal output
flabel metal2 s 5262 11194 5318 11250 0 FreeSans 224 0 0 0 N2BEG[6]
port 114 nsew signal output
flabel metal2 s 5630 11194 5686 11250 0 FreeSans 224 0 0 0 N2BEG[7]
port 115 nsew signal output
flabel metal2 s 5998 11194 6054 11250 0 FreeSans 224 0 0 0 N2BEGb[0]
port 116 nsew signal output
flabel metal2 s 6366 11194 6422 11250 0 FreeSans 224 0 0 0 N2BEGb[1]
port 117 nsew signal output
flabel metal2 s 6734 11194 6790 11250 0 FreeSans 224 0 0 0 N2BEGb[2]
port 118 nsew signal output
flabel metal2 s 7102 11194 7158 11250 0 FreeSans 224 0 0 0 N2BEGb[3]
port 119 nsew signal output
flabel metal2 s 7470 11194 7526 11250 0 FreeSans 224 0 0 0 N2BEGb[4]
port 120 nsew signal output
flabel metal2 s 7838 11194 7894 11250 0 FreeSans 224 0 0 0 N2BEGb[5]
port 121 nsew signal output
flabel metal2 s 8206 11194 8262 11250 0 FreeSans 224 0 0 0 N2BEGb[6]
port 122 nsew signal output
flabel metal2 s 8574 11194 8630 11250 0 FreeSans 224 0 0 0 N2BEGb[7]
port 123 nsew signal output
flabel metal2 s 8942 11194 8998 11250 0 FreeSans 224 0 0 0 N4BEG[0]
port 124 nsew signal output
flabel metal2 s 12622 11194 12678 11250 0 FreeSans 224 0 0 0 N4BEG[10]
port 125 nsew signal output
flabel metal2 s 12990 11194 13046 11250 0 FreeSans 224 0 0 0 N4BEG[11]
port 126 nsew signal output
flabel metal2 s 13358 11194 13414 11250 0 FreeSans 224 0 0 0 N4BEG[12]
port 127 nsew signal output
flabel metal2 s 13726 11194 13782 11250 0 FreeSans 224 0 0 0 N4BEG[13]
port 128 nsew signal output
flabel metal2 s 14094 11194 14150 11250 0 FreeSans 224 0 0 0 N4BEG[14]
port 129 nsew signal output
flabel metal2 s 14462 11194 14518 11250 0 FreeSans 224 0 0 0 N4BEG[15]
port 130 nsew signal output
flabel metal2 s 9310 11194 9366 11250 0 FreeSans 224 0 0 0 N4BEG[1]
port 131 nsew signal output
flabel metal2 s 9678 11194 9734 11250 0 FreeSans 224 0 0 0 N4BEG[2]
port 132 nsew signal output
flabel metal2 s 10046 11194 10102 11250 0 FreeSans 224 0 0 0 N4BEG[3]
port 133 nsew signal output
flabel metal2 s 10414 11194 10470 11250 0 FreeSans 224 0 0 0 N4BEG[4]
port 134 nsew signal output
flabel metal2 s 10782 11194 10838 11250 0 FreeSans 224 0 0 0 N4BEG[5]
port 135 nsew signal output
flabel metal2 s 11150 11194 11206 11250 0 FreeSans 224 0 0 0 N4BEG[6]
port 136 nsew signal output
flabel metal2 s 11518 11194 11574 11250 0 FreeSans 224 0 0 0 N4BEG[7]
port 137 nsew signal output
flabel metal2 s 11886 11194 11942 11250 0 FreeSans 224 0 0 0 N4BEG[8]
port 138 nsew signal output
flabel metal2 s 12254 11194 12310 11250 0 FreeSans 224 0 0 0 N4BEG[9]
port 139 nsew signal output
flabel metal2 s 14830 11194 14886 11250 0 FreeSans 224 0 0 0 NN4BEG[0]
port 140 nsew signal output
flabel metal2 s 18510 11194 18566 11250 0 FreeSans 224 0 0 0 NN4BEG[10]
port 141 nsew signal output
flabel metal2 s 18878 11194 18934 11250 0 FreeSans 224 0 0 0 NN4BEG[11]
port 142 nsew signal output
flabel metal2 s 19246 11194 19302 11250 0 FreeSans 224 0 0 0 NN4BEG[12]
port 143 nsew signal output
flabel metal2 s 19614 11194 19670 11250 0 FreeSans 224 0 0 0 NN4BEG[13]
port 144 nsew signal output
flabel metal2 s 19982 11194 20038 11250 0 FreeSans 224 0 0 0 NN4BEG[14]
port 145 nsew signal output
flabel metal2 s 20350 11194 20406 11250 0 FreeSans 224 0 0 0 NN4BEG[15]
port 146 nsew signal output
flabel metal2 s 15198 11194 15254 11250 0 FreeSans 224 0 0 0 NN4BEG[1]
port 147 nsew signal output
flabel metal2 s 15566 11194 15622 11250 0 FreeSans 224 0 0 0 NN4BEG[2]
port 148 nsew signal output
flabel metal2 s 15934 11194 15990 11250 0 FreeSans 224 0 0 0 NN4BEG[3]
port 149 nsew signal output
flabel metal2 s 16302 11194 16358 11250 0 FreeSans 224 0 0 0 NN4BEG[4]
port 150 nsew signal output
flabel metal2 s 16670 11194 16726 11250 0 FreeSans 224 0 0 0 NN4BEG[5]
port 151 nsew signal output
flabel metal2 s 17038 11194 17094 11250 0 FreeSans 224 0 0 0 NN4BEG[6]
port 152 nsew signal output
flabel metal2 s 17406 11194 17462 11250 0 FreeSans 224 0 0 0 NN4BEG[7]
port 153 nsew signal output
flabel metal2 s 17774 11194 17830 11250 0 FreeSans 224 0 0 0 NN4BEG[8]
port 154 nsew signal output
flabel metal2 s 18142 11194 18198 11250 0 FreeSans 224 0 0 0 NN4BEG[9]
port 155 nsew signal output
flabel metal2 s 20718 11194 20774 11250 0 FreeSans 224 0 0 0 S1END[0]
port 156 nsew signal input
flabel metal2 s 21086 11194 21142 11250 0 FreeSans 224 0 0 0 S1END[1]
port 157 nsew signal input
flabel metal2 s 21454 11194 21510 11250 0 FreeSans 224 0 0 0 S1END[2]
port 158 nsew signal input
flabel metal2 s 21822 11194 21878 11250 0 FreeSans 224 0 0 0 S1END[3]
port 159 nsew signal input
flabel metal2 s 25134 11194 25190 11250 0 FreeSans 224 0 0 0 S2END[0]
port 160 nsew signal input
flabel metal2 s 25502 11194 25558 11250 0 FreeSans 224 0 0 0 S2END[1]
port 161 nsew signal input
flabel metal2 s 25870 11194 25926 11250 0 FreeSans 224 0 0 0 S2END[2]
port 162 nsew signal input
flabel metal2 s 26238 11194 26294 11250 0 FreeSans 224 0 0 0 S2END[3]
port 163 nsew signal input
flabel metal2 s 26606 11194 26662 11250 0 FreeSans 224 0 0 0 S2END[4]
port 164 nsew signal input
flabel metal2 s 26974 11194 27030 11250 0 FreeSans 224 0 0 0 S2END[5]
port 165 nsew signal input
flabel metal2 s 27342 11194 27398 11250 0 FreeSans 224 0 0 0 S2END[6]
port 166 nsew signal input
flabel metal2 s 27710 11194 27766 11250 0 FreeSans 224 0 0 0 S2END[7]
port 167 nsew signal input
flabel metal2 s 22190 11194 22246 11250 0 FreeSans 224 0 0 0 S2MID[0]
port 168 nsew signal input
flabel metal2 s 22558 11194 22614 11250 0 FreeSans 224 0 0 0 S2MID[1]
port 169 nsew signal input
flabel metal2 s 22926 11194 22982 11250 0 FreeSans 224 0 0 0 S2MID[2]
port 170 nsew signal input
flabel metal2 s 23294 11194 23350 11250 0 FreeSans 224 0 0 0 S2MID[3]
port 171 nsew signal input
flabel metal2 s 23662 11194 23718 11250 0 FreeSans 224 0 0 0 S2MID[4]
port 172 nsew signal input
flabel metal2 s 24030 11194 24086 11250 0 FreeSans 224 0 0 0 S2MID[5]
port 173 nsew signal input
flabel metal2 s 24398 11194 24454 11250 0 FreeSans 224 0 0 0 S2MID[6]
port 174 nsew signal input
flabel metal2 s 24766 11194 24822 11250 0 FreeSans 224 0 0 0 S2MID[7]
port 175 nsew signal input
flabel metal2 s 28078 11194 28134 11250 0 FreeSans 224 0 0 0 S4END[0]
port 176 nsew signal input
flabel metal2 s 31758 11194 31814 11250 0 FreeSans 224 0 0 0 S4END[10]
port 177 nsew signal input
flabel metal2 s 32126 11194 32182 11250 0 FreeSans 224 0 0 0 S4END[11]
port 178 nsew signal input
flabel metal2 s 32494 11194 32550 11250 0 FreeSans 224 0 0 0 S4END[12]
port 179 nsew signal input
flabel metal2 s 32862 11194 32918 11250 0 FreeSans 224 0 0 0 S4END[13]
port 180 nsew signal input
flabel metal2 s 33230 11194 33286 11250 0 FreeSans 224 0 0 0 S4END[14]
port 181 nsew signal input
flabel metal2 s 33598 11194 33654 11250 0 FreeSans 224 0 0 0 S4END[15]
port 182 nsew signal input
flabel metal2 s 28446 11194 28502 11250 0 FreeSans 224 0 0 0 S4END[1]
port 183 nsew signal input
flabel metal2 s 28814 11194 28870 11250 0 FreeSans 224 0 0 0 S4END[2]
port 184 nsew signal input
flabel metal2 s 29182 11194 29238 11250 0 FreeSans 224 0 0 0 S4END[3]
port 185 nsew signal input
flabel metal2 s 29550 11194 29606 11250 0 FreeSans 224 0 0 0 S4END[4]
port 186 nsew signal input
flabel metal2 s 29918 11194 29974 11250 0 FreeSans 224 0 0 0 S4END[5]
port 187 nsew signal input
flabel metal2 s 30286 11194 30342 11250 0 FreeSans 224 0 0 0 S4END[6]
port 188 nsew signal input
flabel metal2 s 30654 11194 30710 11250 0 FreeSans 224 0 0 0 S4END[7]
port 189 nsew signal input
flabel metal2 s 31022 11194 31078 11250 0 FreeSans 224 0 0 0 S4END[8]
port 190 nsew signal input
flabel metal2 s 31390 11194 31446 11250 0 FreeSans 224 0 0 0 S4END[9]
port 191 nsew signal input
flabel metal2 s 33966 11194 34022 11250 0 FreeSans 224 0 0 0 SS4END[0]
port 192 nsew signal input
flabel metal2 s 37646 11194 37702 11250 0 FreeSans 224 0 0 0 SS4END[10]
port 193 nsew signal input
flabel metal2 s 38014 11194 38070 11250 0 FreeSans 224 0 0 0 SS4END[11]
port 194 nsew signal input
flabel metal2 s 38382 11194 38438 11250 0 FreeSans 224 0 0 0 SS4END[12]
port 195 nsew signal input
flabel metal2 s 38750 11194 38806 11250 0 FreeSans 224 0 0 0 SS4END[13]
port 196 nsew signal input
flabel metal2 s 39118 11194 39174 11250 0 FreeSans 224 0 0 0 SS4END[14]
port 197 nsew signal input
flabel metal2 s 39486 11194 39542 11250 0 FreeSans 224 0 0 0 SS4END[15]
port 198 nsew signal input
flabel metal2 s 34334 11194 34390 11250 0 FreeSans 224 0 0 0 SS4END[1]
port 199 nsew signal input
flabel metal2 s 34702 11194 34758 11250 0 FreeSans 224 0 0 0 SS4END[2]
port 200 nsew signal input
flabel metal2 s 35070 11194 35126 11250 0 FreeSans 224 0 0 0 SS4END[3]
port 201 nsew signal input
flabel metal2 s 35438 11194 35494 11250 0 FreeSans 224 0 0 0 SS4END[4]
port 202 nsew signal input
flabel metal2 s 35806 11194 35862 11250 0 FreeSans 224 0 0 0 SS4END[5]
port 203 nsew signal input
flabel metal2 s 36174 11194 36230 11250 0 FreeSans 224 0 0 0 SS4END[6]
port 204 nsew signal input
flabel metal2 s 36542 11194 36598 11250 0 FreeSans 224 0 0 0 SS4END[7]
port 205 nsew signal input
flabel metal2 s 36910 11194 36966 11250 0 FreeSans 224 0 0 0 SS4END[8]
port 206 nsew signal input
flabel metal2 s 37278 11194 37334 11250 0 FreeSans 224 0 0 0 SS4END[9]
port 207 nsew signal input
flabel metal2 s 1398 0 1454 56 0 FreeSans 224 0 0 0 UserCLK
port 208 nsew signal input
flabel metal2 s 39854 11194 39910 11250 0 FreeSans 224 0 0 0 UserCLKo
port 209 nsew signal output
flabel metal4 s 3004 0 3324 11250 0 FreeSans 1920 90 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 3004 0 3324 60 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 3004 11190 3324 11250 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 9004 0 9324 11250 0 FreeSans 1920 90 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 9004 0 9324 60 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 9004 11190 9324 11250 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 15004 0 15324 11250 0 FreeSans 1920 90 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 15004 0 15324 60 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 15004 11190 15324 11250 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 21004 0 21324 11250 0 FreeSans 1920 90 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 21004 0 21324 60 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 21004 11190 21324 11250 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 27004 0 27324 11250 0 FreeSans 1920 90 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 27004 0 27324 60 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 27004 11190 27324 11250 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 33004 0 33324 11250 0 FreeSans 1920 90 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 33004 0 33324 60 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 33004 11190 33324 11250 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 39004 0 39324 11250 0 FreeSans 1920 90 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 39004 0 39324 60 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 39004 11190 39324 11250 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 45004 0 45324 11250 0 FreeSans 1920 90 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 45004 0 45324 60 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 45004 11190 45324 11250 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 1944 0 2264 11250 0 FreeSans 1920 90 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 1944 0 2264 60 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 1944 11190 2264 11250 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 7944 0 8264 11250 0 FreeSans 1920 90 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 7944 0 8264 60 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 7944 11190 8264 11250 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 13944 0 14264 11250 0 FreeSans 1920 90 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 13944 0 14264 60 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 13944 11190 14264 11250 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 19944 0 20264 11250 0 FreeSans 1920 90 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 19944 0 20264 60 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 19944 11190 20264 11250 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 25944 0 26264 11250 0 FreeSans 1920 90 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 25944 0 26264 60 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 25944 11190 26264 11250 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 31944 0 32264 11250 0 FreeSans 1920 90 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 31944 0 32264 60 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 31944 11190 32264 11250 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 37944 0 38264 11250 0 FreeSans 1920 90 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 37944 0 38264 60 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 37944 11190 38264 11250 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 43944 0 44264 11250 0 FreeSans 1920 90 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 43944 0 44264 60 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 43944 11190 44264 11250 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
rlabel metal1 24472 8704 24472 8704 0 VGND
rlabel metal1 24472 8160 24472 8160 0 VPWR
rlabel metal3 712 1428 712 1428 0 FrameData[0]
rlabel metal1 25024 6086 25024 6086 0 FrameData[10]
rlabel metal2 13662 5695 13662 5695 0 FrameData[11]
rlabel metal4 14812 6460 14812 6460 0 FrameData[12]
rlabel metal3 919 4964 919 4964 0 FrameData[13]
rlabel metal3 1402 5236 1402 5236 0 FrameData[14]
rlabel metal2 17434 5253 17434 5253 0 FrameData[15]
rlabel metal1 19964 4794 19964 4794 0 FrameData[16]
rlabel metal3 919 6052 919 6052 0 FrameData[17]
rlabel metal1 14674 5678 14674 5678 0 FrameData[18]
rlabel metal1 14122 2074 14122 2074 0 FrameData[19]
rlabel metal3 4852 1700 4852 1700 0 FrameData[1]
rlabel metal1 15640 3162 15640 3162 0 FrameData[20]
rlabel metal3 919 7140 919 7140 0 FrameData[21]
rlabel metal3 620 7412 620 7412 0 FrameData[22]
rlabel metal3 20516 7140 20516 7140 0 FrameData[23]
rlabel metal1 36524 3026 36524 3026 0 FrameData[24]
rlabel metal3 712 8228 712 8228 0 FrameData[25]
rlabel metal2 41630 8279 41630 8279 0 FrameData[26]
rlabel metal3 1425 8772 1425 8772 0 FrameData[27]
rlabel metal2 30222 8551 30222 8551 0 FrameData[28]
rlabel metal3 160 9316 160 9316 0 FrameData[29]
rlabel metal3 9912 1972 9912 1972 0 FrameData[2]
rlabel metal2 5198 8721 5198 8721 0 FrameData[30]
rlabel metal2 34454 9503 34454 9503 0 FrameData[31]
rlabel metal3 1471 2244 1471 2244 0 FrameData[3]
rlabel metal3 4806 2516 4806 2516 0 FrameData[4]
rlabel metal3 919 2788 919 2788 0 FrameData[5]
rlabel metal2 17250 3859 17250 3859 0 FrameData[6]
rlabel metal2 20746 3689 20746 3689 0 FrameData[7]
rlabel metal2 24886 4029 24886 4029 0 FrameData[8]
rlabel metal3 919 3876 919 3876 0 FrameData[9]
rlabel metal3 47754 1428 47754 1428 0 FrameData_O[0]
rlabel metal3 48122 4148 48122 4148 0 FrameData_O[10]
rlabel metal3 47984 4420 47984 4420 0 FrameData_O[11]
rlabel metal3 48168 4692 48168 4692 0 FrameData_O[12]
rlabel metal3 47938 4964 47938 4964 0 FrameData_O[13]
rlabel metal3 48122 5236 48122 5236 0 FrameData_O[14]
rlabel metal3 47984 5508 47984 5508 0 FrameData_O[15]
rlabel metal3 47754 5780 47754 5780 0 FrameData_O[16]
rlabel metal2 47426 5967 47426 5967 0 FrameData_O[17]
rlabel metal3 47616 6324 47616 6324 0 FrameData_O[18]
rlabel metal2 46966 6511 46966 6511 0 FrameData_O[19]
rlabel metal3 47570 1700 47570 1700 0 FrameData_O[1]
rlabel metal3 47800 6868 47800 6868 0 FrameData_O[20]
rlabel metal2 47426 6885 47426 6885 0 FrameData_O[21]
rlabel metal3 47938 7412 47938 7412 0 FrameData_O[22]
rlabel metal2 47334 7599 47334 7599 0 FrameData_O[23]
rlabel metal3 47478 7956 47478 7956 0 FrameData_O[24]
rlabel metal2 46598 7871 46598 7871 0 FrameData_O[25]
rlabel metal2 47058 7565 47058 7565 0 FrameData_O[26]
rlabel metal1 46276 7174 46276 7174 0 FrameData_O[27]
rlabel metal2 45678 8551 45678 8551 0 FrameData_O[28]
rlabel metal1 45908 7174 45908 7174 0 FrameData_O[29]
rlabel metal3 47386 1972 47386 1972 0 FrameData_O[2]
rlabel metal1 45080 8058 45080 8058 0 FrameData_O[30]
rlabel metal1 47426 6426 47426 6426 0 FrameData_O[31]
rlabel metal3 47938 2244 47938 2244 0 FrameData_O[3]
rlabel metal3 48122 2516 48122 2516 0 FrameData_O[4]
rlabel metal3 47938 2788 47938 2788 0 FrameData_O[5]
rlabel metal3 48122 3060 48122 3060 0 FrameData_O[6]
rlabel metal3 47984 3332 47984 3332 0 FrameData_O[7]
rlabel metal3 48168 3604 48168 3604 0 FrameData_O[8]
rlabel metal3 47938 3876 47938 3876 0 FrameData_O[9]
rlabel metal2 3726 106 3726 106 0 FrameStrobe[0]
rlabel metal1 28014 3162 28014 3162 0 FrameStrobe[10]
rlabel metal2 29026 1823 29026 1823 0 FrameStrobe[11]
rlabel metal2 31326 1058 31326 1058 0 FrameStrobe[12]
rlabel metal2 33626 1704 33626 1704 0 FrameStrobe[13]
rlabel metal2 35926 3744 35926 3744 0 FrameStrobe[14]
rlabel metal2 38226 735 38226 735 0 FrameStrobe[15]
rlabel metal2 40526 3676 40526 3676 0 FrameStrobe[16]
rlabel metal1 43608 7310 43608 7310 0 FrameStrobe[17]
rlabel metal2 45126 55 45126 55 0 FrameStrobe[18]
rlabel metal2 47426 55 47426 55 0 FrameStrobe[19]
rlabel metal2 6026 106 6026 106 0 FrameStrobe[1]
rlabel metal1 8556 3094 8556 3094 0 FrameStrobe[2]
rlabel metal1 10764 3026 10764 3026 0 FrameStrobe[3]
rlabel metal1 12834 3026 12834 3026 0 FrameStrobe[4]
rlabel metal2 15226 55 15226 55 0 FrameStrobe[5]
rlabel metal1 18124 2958 18124 2958 0 FrameStrobe[6]
rlabel metal1 20884 3094 20884 3094 0 FrameStrobe[7]
rlabel metal1 23368 3502 23368 3502 0 FrameStrobe[8]
rlabel metal1 25852 3094 25852 3094 0 FrameStrobe[9]
rlabel metal1 40388 8602 40388 8602 0 FrameStrobe_O[0]
rlabel metal1 44206 8602 44206 8602 0 FrameStrobe_O[10]
rlabel metal1 44758 8330 44758 8330 0 FrameStrobe_O[11]
rlabel metal1 45126 8602 45126 8602 0 FrameStrobe_O[12]
rlabel metal1 45954 8568 45954 8568 0 FrameStrobe_O[13]
rlabel metal1 46368 8330 46368 8330 0 FrameStrobe_O[14]
rlabel metal1 46368 8602 46368 8602 0 FrameStrobe_O[15]
rlabel metal1 47058 8364 47058 8364 0 FrameStrobe_O[16]
rlabel metal1 46644 8058 46644 8058 0 FrameStrobe_O[17]
rlabel metal1 47012 8058 47012 8058 0 FrameStrobe_O[18]
rlabel metal1 46828 7990 46828 7990 0 FrameStrobe_O[19]
rlabel metal1 40756 8602 40756 8602 0 FrameStrobe_O[1]
rlabel metal1 41124 8602 41124 8602 0 FrameStrobe_O[2]
rlabel metal2 41354 9904 41354 9904 0 FrameStrobe_O[3]
rlabel metal1 41860 8602 41860 8602 0 FrameStrobe_O[4]
rlabel metal1 42366 8602 42366 8602 0 FrameStrobe_O[5]
rlabel metal1 42734 8330 42734 8330 0 FrameStrobe_O[6]
rlabel metal1 43102 8602 43102 8602 0 FrameStrobe_O[7]
rlabel metal1 43470 8330 43470 8330 0 FrameStrobe_O[8]
rlabel metal1 44114 8364 44114 8364 0 FrameStrobe_O[9]
rlabel metal2 1610 9632 1610 9632 0 N1BEG[0]
rlabel metal1 1886 8602 1886 8602 0 N1BEG[1]
rlabel metal1 2254 8602 2254 8602 0 N1BEG[2]
rlabel metal1 2622 8602 2622 8602 0 N1BEG[3]
rlabel metal1 2990 8602 2990 8602 0 N2BEG[0]
rlabel metal2 3450 9904 3450 9904 0 N2BEG[1]
rlabel metal1 3910 8058 3910 8058 0 N2BEG[2]
rlabel metal2 4186 9904 4186 9904 0 N2BEG[3]
rlabel metal2 4554 9904 4554 9904 0 N2BEG[4]
rlabel metal2 4922 9904 4922 9904 0 N2BEG[5]
rlabel metal2 5290 9904 5290 9904 0 N2BEG[6]
rlabel metal2 5658 9904 5658 9904 0 N2BEG[7]
rlabel metal2 6026 9904 6026 9904 0 N2BEGb[0]
rlabel metal1 6486 8058 6486 8058 0 N2BEGb[1]
rlabel metal2 6762 9904 6762 9904 0 N2BEGb[2]
rlabel metal2 7130 9904 7130 9904 0 N2BEGb[3]
rlabel metal2 7498 9904 7498 9904 0 N2BEGb[4]
rlabel metal2 7866 9904 7866 9904 0 N2BEGb[5]
rlabel metal2 8234 9904 8234 9904 0 N2BEGb[6]
rlabel metal2 8602 9904 8602 9904 0 N2BEGb[7]
rlabel metal1 9016 8058 9016 8058 0 N4BEG[0]
rlabel metal2 12650 9904 12650 9904 0 N4BEG[10]
rlabel metal2 13018 9904 13018 9904 0 N4BEG[11]
rlabel metal1 13432 8602 13432 8602 0 N4BEG[12]
rlabel metal1 13800 8602 13800 8602 0 N4BEG[13]
rlabel metal1 14352 8058 14352 8058 0 N4BEG[14]
rlabel metal1 14536 8602 14536 8602 0 N4BEG[15]
rlabel metal1 9384 8602 9384 8602 0 N4BEG[1]
rlabel metal2 9706 9904 9706 9904 0 N4BEG[2]
rlabel metal2 10074 9904 10074 9904 0 N4BEG[3]
rlabel metal2 10442 9904 10442 9904 0 N4BEG[4]
rlabel metal2 10810 9904 10810 9904 0 N4BEG[5]
rlabel metal2 11178 9904 11178 9904 0 N4BEG[6]
rlabel metal1 11960 8058 11960 8058 0 N4BEG[7]
rlabel metal2 11914 9904 11914 9904 0 N4BEG[8]
rlabel metal2 12282 9904 12282 9904 0 N4BEG[9]
rlabel metal1 14904 8602 14904 8602 0 NN4BEG[0]
rlabel metal1 18354 8602 18354 8602 0 NN4BEG[10]
rlabel metal1 18722 8330 18722 8330 0 NN4BEG[11]
rlabel metal1 19090 8602 19090 8602 0 NN4BEG[12]
rlabel metal2 19642 9904 19642 9904 0 NN4BEG[13]
rlabel metal1 20102 8602 20102 8602 0 NN4BEG[14]
rlabel metal1 20470 8602 20470 8602 0 NN4BEG[15]
rlabel metal1 15364 8602 15364 8602 0 NN4BEG[1]
rlabel metal1 15640 8602 15640 8602 0 NN4BEG[2]
rlabel metal1 16008 8602 16008 8602 0 NN4BEG[3]
rlabel metal1 16376 8602 16376 8602 0 NN4BEG[4]
rlabel metal1 16836 8058 16836 8058 0 NN4BEG[5]
rlabel metal1 17204 8058 17204 8058 0 NN4BEG[6]
rlabel metal1 17296 8602 17296 8602 0 NN4BEG[7]
rlabel metal1 17434 8364 17434 8364 0 NN4BEG[8]
rlabel metal1 17940 8602 17940 8602 0 NN4BEG[9]
rlabel metal2 20746 10465 20746 10465 0 S1END[0]
rlabel metal2 21114 10057 21114 10057 0 S1END[1]
rlabel metal2 21482 7660 21482 7660 0 S1END[2]
rlabel metal2 21850 7626 21850 7626 0 S1END[3]
rlabel metal2 25162 8748 25162 8748 0 S2END[0]
rlabel metal2 25530 9989 25530 9989 0 S2END[1]
rlabel metal2 25898 8714 25898 8714 0 S2END[2]
rlabel metal2 26266 10261 26266 10261 0 S2END[3]
rlabel metal2 26634 9530 26634 9530 0 S2END[4]
rlabel metal2 27002 10397 27002 10397 0 S2END[5]
rlabel metal2 27370 9530 27370 9530 0 S2END[6]
rlabel metal2 27738 9564 27738 9564 0 S2END[7]
rlabel metal2 18262 5457 18262 5457 0 S2MID[0]
rlabel metal1 20194 3468 20194 3468 0 S2MID[1]
rlabel metal1 21022 4624 21022 4624 0 S2MID[2]
rlabel metal2 23322 9581 23322 9581 0 S2MID[3]
rlabel metal1 21574 5236 21574 5236 0 S2MID[4]
rlabel metal2 21942 7956 21942 7956 0 S2MID[5]
rlabel metal2 24426 8442 24426 8442 0 S2MID[6]
rlabel metal2 24794 8204 24794 8204 0 S2MID[7]
rlabel metal1 14214 7718 14214 7718 0 S4END[0]
rlabel metal2 31786 8986 31786 8986 0 S4END[10]
rlabel metal2 32154 10261 32154 10261 0 S4END[11]
rlabel metal2 32522 9530 32522 9530 0 S4END[12]
rlabel metal2 32890 8986 32890 8986 0 S4END[13]
rlabel metal2 33258 10057 33258 10057 0 S4END[14]
rlabel metal2 33626 8204 33626 8204 0 S4END[15]
rlabel metal2 12006 9333 12006 9333 0 S4END[1]
rlabel metal1 10856 8058 10856 8058 0 S4END[2]
rlabel metal2 11822 9418 11822 9418 0 S4END[3]
rlabel metal2 29578 9564 29578 9564 0 S4END[4]
rlabel metal2 29946 9530 29946 9530 0 S4END[5]
rlabel metal2 30314 8986 30314 8986 0 S4END[6]
rlabel metal2 30682 8476 30682 8476 0 S4END[7]
rlabel metal2 31050 8442 31050 8442 0 S4END[8]
rlabel metal2 31418 8442 31418 8442 0 S4END[9]
rlabel metal2 33994 8442 33994 8442 0 SS4END[0]
rlabel metal1 15778 6766 15778 6766 0 SS4END[10]
rlabel metal1 16192 7378 16192 7378 0 SS4END[11]
rlabel metal2 38410 10142 38410 10142 0 SS4END[12]
rlabel metal2 14950 9248 14950 9248 0 SS4END[13]
rlabel metal2 14582 8432 14582 8432 0 SS4END[14]
rlabel metal2 13570 9520 13570 9520 0 SS4END[15]
rlabel metal2 34362 8748 34362 8748 0 SS4END[1]
rlabel metal2 34730 9564 34730 9564 0 SS4END[2]
rlabel metal2 35098 9632 35098 9632 0 SS4END[3]
rlabel metal1 20424 7854 20424 7854 0 SS4END[4]
rlabel metal1 19734 7854 19734 7854 0 SS4END[5]
rlabel metal2 18354 9384 18354 9384 0 SS4END[6]
rlabel metal2 18262 9452 18262 9452 0 SS4END[7]
rlabel metal2 19182 8296 19182 8296 0 SS4END[8]
rlabel viali 16330 6766 16330 6766 0 SS4END[9]
rlabel metal2 1426 55 1426 55 0 UserCLK
rlabel metal1 39928 8602 39928 8602 0 UserCLKo
rlabel metal2 8602 2652 8602 2652 0 net1
rlabel via2 14950 5661 14950 5661 0 net10
rlabel metal1 15778 6664 15778 6664 0 net100
rlabel metal1 16836 6630 16836 6630 0 net101
rlabel metal1 17066 7514 17066 7514 0 net102
rlabel metal1 17710 8058 17710 8058 0 net103
rlabel metal1 18078 8058 18078 8058 0 net104
rlabel metal2 38778 5814 38778 5814 0 net105
rlabel metal1 26036 2822 26036 2822 0 net11
rlabel metal2 13294 2686 13294 2686 0 net12
rlabel metal2 18170 4080 18170 4080 0 net13
rlabel metal2 32798 5967 32798 5967 0 net14
rlabel metal2 37674 3366 37674 3366 0 net15
rlabel metal2 23138 3910 23138 3910 0 net16
rlabel metal2 36938 4896 36938 4896 0 net17
rlabel metal2 33166 5916 33166 5916 0 net18
rlabel metal1 46874 6800 46874 6800 0 net19
rlabel metal2 34454 5610 34454 5610 0 net2
rlabel metal1 8142 7446 8142 7446 0 net20
rlabel metal2 39606 7650 39606 7650 0 net21
rlabel via2 2438 7837 2438 7837 0 net22
rlabel metal2 20470 2720 20470 2720 0 net23
rlabel via2 5382 7973 5382 7973 0 net24
rlabel metal1 47150 6256 47150 6256 0 net25
rlabel metal1 31740 2312 31740 2312 0 net26
rlabel metal2 16882 2686 16882 2686 0 net27
rlabel metal2 28566 3213 28566 3213 0 net28
rlabel metal1 23598 4488 23598 4488 0 net29
rlabel metal1 36478 6392 36478 6392 0 net3
rlabel metal2 25898 3689 25898 3689 0 net30
rlabel metal2 25254 4352 25254 4352 0 net31
rlabel metal1 31740 4046 31740 4046 0 net32
rlabel metal2 39698 5780 39698 5780 0 net33
rlabel metal2 35834 5610 35834 5610 0 net34
rlabel metal1 43056 7514 43056 7514 0 net35
rlabel metal2 43286 6018 43286 6018 0 net36
rlabel metal1 43976 3162 43976 3162 0 net37
rlabel metal1 44528 7242 44528 7242 0 net38
rlabel metal2 39974 8126 39974 8126 0 net39
rlabel metal1 47242 4624 47242 4624 0 net4
rlabel metal1 42826 7242 42826 7242 0 net40
rlabel metal2 44574 7718 44574 7718 0 net41
rlabel metal1 46138 7242 46138 7242 0 net42
rlabel metal1 45770 7514 45770 7514 0 net43
rlabel metal1 40618 3162 40618 3162 0 net44
rlabel metal1 41078 8500 41078 8500 0 net45
rlabel metal2 41354 3944 41354 3944 0 net46
rlabel metal2 12834 3400 12834 3400 0 net47
rlabel metal1 18998 2856 18998 2856 0 net48
rlabel metal1 18906 2924 18906 2924 0 net49
rlabel metal2 21758 6392 21758 6392 0 net5
rlabel metal1 31878 2992 31878 2992 0 net50
rlabel metal2 43378 6086 43378 6086 0 net51
rlabel metal2 40802 6120 40802 6120 0 net52
rlabel metal1 1794 7888 1794 7888 0 net53
rlabel metal1 15732 3910 15732 3910 0 net54
rlabel metal2 2346 5950 2346 5950 0 net55
rlabel metal1 2668 8466 2668 8466 0 net56
rlabel metal1 23552 5338 23552 5338 0 net57
rlabel metal2 6854 7208 6854 7208 0 net58
rlabel metal1 17802 5338 17802 5338 0 net59
rlabel metal2 18814 6426 18814 6426 0 net6
rlabel metal1 20884 4998 20884 4998 0 net60
rlabel metal1 21298 4488 21298 4488 0 net61
rlabel metal2 8694 6766 8694 6766 0 net62
rlabel metal1 20010 3400 20010 3400 0 net63
rlabel metal2 18078 5695 18078 5695 0 net64
rlabel metal1 17250 9248 17250 9248 0 net65
rlabel metal2 6762 7582 6762 7582 0 net66
rlabel metal1 12558 8296 12558 8296 0 net67
rlabel metal1 7498 8398 7498 8398 0 net68
rlabel metal2 7682 7854 7682 7854 0 net69
rlabel metal2 17802 6358 17802 6358 0 net7
rlabel metal2 7866 7344 7866 7344 0 net70
rlabel metal2 8418 7310 8418 7310 0 net71
rlabel metal2 16882 7820 16882 7820 0 net72
rlabel metal2 14858 5236 14858 5236 0 net73
rlabel metal2 18906 7684 18906 7684 0 net74
rlabel metal2 16330 7548 16330 7548 0 net75
rlabel metal1 13294 8500 13294 8500 0 net76
rlabel metal2 13662 8228 13662 8228 0 net77
rlabel metal1 14214 7820 14214 7820 0 net78
rlabel metal1 13432 8058 13432 8058 0 net79
rlabel metal2 24978 5202 24978 5202 0 net8
rlabel metal3 13708 6120 13708 6120 0 net80
rlabel metal2 35374 6681 35374 6681 0 net81
rlabel metal2 18998 8262 18998 8262 0 net82
rlabel metal2 14858 7038 14858 7038 0 net83
rlabel metal2 10994 7412 10994 7412 0 net84
rlabel metal2 12466 8279 12466 8279 0 net85
rlabel metal2 19366 6358 19366 6358 0 net86
rlabel metal2 12650 7106 12650 7106 0 net87
rlabel metal2 17250 6562 17250 6562 0 net88
rlabel metal1 14214 7990 14214 7990 0 net89
rlabel metal1 31970 3094 31970 3094 0 net9
rlabel metal2 19458 8296 19458 8296 0 net90
rlabel metal1 19964 8058 19964 8058 0 net91
rlabel metal2 19734 8704 19734 8704 0 net92
rlabel metal1 19826 8432 19826 8432 0 net93
rlabel metal1 20194 8466 20194 8466 0 net94
rlabel metal1 20838 8466 20838 8466 0 net95
rlabel metal1 14950 8058 14950 8058 0 net96
rlabel metal1 15088 7514 15088 7514 0 net97
rlabel metal1 15778 7514 15778 7514 0 net98
rlabel metal1 16100 7514 16100 7514 0 net99
<< properties >>
string FIXED_BBOX 0 0 49000 11250
<< end >>
