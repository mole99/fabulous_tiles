* NGSPICE file created from N_IO.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlxtp_1 abstract view
.subckt sky130_fd_sc_hd__dlxtp_1 D GATE VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_1 abstract view
.subckt sky130_fd_sc_hd__inv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

.subckt N_IO A_I_top A_O_top A_T_top A_config_C_bit0 A_config_C_bit1 A_config_C_bit2
+ A_config_C_bit3 B_I_top B_O_top B_T_top B_config_C_bit0 B_config_C_bit1 B_config_C_bit2
+ B_config_C_bit3 Ci FrameData[0] FrameData[10] FrameData[11] FrameData[12] FrameData[13]
+ FrameData[14] FrameData[15] FrameData[16] FrameData[17] FrameData[18] FrameData[19]
+ FrameData[1] FrameData[20] FrameData[21] FrameData[22] FrameData[23] FrameData[24]
+ FrameData[25] FrameData[26] FrameData[27] FrameData[28] FrameData[29] FrameData[2]
+ FrameData[30] FrameData[31] FrameData[3] FrameData[4] FrameData[5] FrameData[6]
+ FrameData[7] FrameData[8] FrameData[9] FrameData_O[0] FrameData_O[10] FrameData_O[11]
+ FrameData_O[12] FrameData_O[13] FrameData_O[14] FrameData_O[15] FrameData_O[16]
+ FrameData_O[17] FrameData_O[18] FrameData_O[19] FrameData_O[1] FrameData_O[20] FrameData_O[21]
+ FrameData_O[22] FrameData_O[23] FrameData_O[24] FrameData_O[25] FrameData_O[26]
+ FrameData_O[27] FrameData_O[28] FrameData_O[29] FrameData_O[2] FrameData_O[30] FrameData_O[31]
+ FrameData_O[3] FrameData_O[4] FrameData_O[5] FrameData_O[6] FrameData_O[7] FrameData_O[8]
+ FrameData_O[9] FrameStrobe[0] FrameStrobe[10] FrameStrobe[11] FrameStrobe[12] FrameStrobe[13]
+ FrameStrobe[14] FrameStrobe[15] FrameStrobe[16] FrameStrobe[17] FrameStrobe[18]
+ FrameStrobe[19] FrameStrobe[1] FrameStrobe[2] FrameStrobe[3] FrameStrobe[4] FrameStrobe[5]
+ FrameStrobe[6] FrameStrobe[7] FrameStrobe[8] FrameStrobe[9] FrameStrobe_O[0] FrameStrobe_O[10]
+ FrameStrobe_O[11] FrameStrobe_O[12] FrameStrobe_O[13] FrameStrobe_O[14] FrameStrobe_O[15]
+ FrameStrobe_O[16] FrameStrobe_O[17] FrameStrobe_O[18] FrameStrobe_O[19] FrameStrobe_O[1]
+ FrameStrobe_O[2] FrameStrobe_O[3] FrameStrobe_O[4] FrameStrobe_O[5] FrameStrobe_O[6]
+ FrameStrobe_O[7] FrameStrobe_O[8] FrameStrobe_O[9] N1END[0] N1END[1] N1END[2] N1END[3]
+ N2END[0] N2END[1] N2END[2] N2END[3] N2END[4] N2END[5] N2END[6] N2END[7] N2MID[0]
+ N2MID[1] N2MID[2] N2MID[3] N2MID[4] N2MID[5] N2MID[6] N2MID[7] N4END[0] N4END[10]
+ N4END[11] N4END[12] N4END[13] N4END[14] N4END[15] N4END[1] N4END[2] N4END[3] N4END[4]
+ N4END[5] N4END[6] N4END[7] N4END[8] N4END[9] NN4END[0] NN4END[10] NN4END[11] NN4END[12]
+ NN4END[13] NN4END[14] NN4END[15] NN4END[1] NN4END[2] NN4END[3] NN4END[4] NN4END[5]
+ NN4END[6] NN4END[7] NN4END[8] NN4END[9] S1BEG[0] S1BEG[1] S1BEG[2] S1BEG[3] S2BEG[0]
+ S2BEG[1] S2BEG[2] S2BEG[3] S2BEG[4] S2BEG[5] S2BEG[6] S2BEG[7] S2BEGb[0] S2BEGb[1]
+ S2BEGb[2] S2BEGb[3] S2BEGb[4] S2BEGb[5] S2BEGb[6] S2BEGb[7] S4BEG[0] S4BEG[10] S4BEG[11]
+ S4BEG[12] S4BEG[13] S4BEG[14] S4BEG[15] S4BEG[1] S4BEG[2] S4BEG[3] S4BEG[4] S4BEG[5]
+ S4BEG[6] S4BEG[7] S4BEG[8] S4BEG[9] SS4BEG[0] SS4BEG[10] SS4BEG[11] SS4BEG[12] SS4BEG[13]
+ SS4BEG[14] SS4BEG[15] SS4BEG[1] SS4BEG[2] SS4BEG[3] SS4BEG[4] SS4BEG[5] SS4BEG[6]
+ SS4BEG[7] SS4BEG[8] SS4BEG[9] UserCLK UserCLKo VGND VPWR
X_294_ FrameStrobe[18] VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__clkbuf_1
XFILLER_5_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_8_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_0_Left_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_346_ Inst_N_IO_switch_matrix.SS4BEG14 VGND VGND VPWR VPWR net209 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_11_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_277_ net63 VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__clkbuf_1
X_131_ net11 net54 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame3_bit17.Q sky130_fd_sc_hd__dlxtp_1
X_200_ net17 net62 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame1_bit22.Q sky130_fd_sc_hd__dlxtp_1
X_062_ Inst_N_IO_ConfigMem.Inst_frame0_bit27.Q _006_ VGND VGND VPWR VPWR _007_ sky130_fd_sc_hd__or2_1
X_329_ Inst_N_IO_switch_matrix.S4BEG13 VGND VGND VPWR VPWR net192 sky130_fd_sc_hd__clkbuf_1
XFILLER_11_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_045_ net43 Inst_N_IO_ConfigMem.Inst_frame0_bit23.Q Inst_N_IO_ConfigMem.Inst_frame0_bit24.Q
+ VGND VGND VPWR VPWR _024_ sky130_fd_sc_hd__o21ai_1
X_114_ net44 net83 net99 net92 Inst_N_IO_ConfigMem.Inst_frame2_bit6.Q Inst_N_IO_ConfigMem.Inst_frame2_bit7.Q
+ VGND VGND VPWR VPWR Inst_N_IO_switch_matrix.S2BEGb2 sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_5_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_5 net143 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput97 net114 VGND VGND VPWR VPWR B_config_C_bit2 sky130_fd_sc_hd__buf_2
XFILLER_8_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_2_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_293_ FrameStrobe[17] VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__clkbuf_1
XFILLER_2_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_276_ net68 VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__clkbuf_1
X_345_ Inst_N_IO_switch_matrix.SS4BEG13 VGND VGND VPWR VPWR net208 sky130_fd_sc_hd__clkbuf_1
X_130_ net10 net54 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame3_bit16.Q sky130_fd_sc_hd__dlxtp_1
X_259_ net9 VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__clkbuf_2
X_061_ net39 net40 net41 net42 Inst_N_IO_ConfigMem.Inst_frame0_bit25.Q Inst_N_IO_ConfigMem.Inst_frame0_bit26.Q
+ VGND VGND VPWR VPWR _006_ sky130_fd_sc_hd__mux4_1
X_328_ Inst_N_IO_switch_matrix.S4BEG12 VGND VGND VPWR VPWR net191 sky130_fd_sc_hd__clkbuf_1
XFILLER_4_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_113_ net43 net82 net98 net91 Inst_N_IO_ConfigMem.Inst_frame2_bit8.Q Inst_N_IO_ConfigMem.Inst_frame2_bit9.Q
+ VGND VGND VPWR VPWR Inst_N_IO_switch_matrix.S2BEGb3 sky130_fd_sc_hd__mux4_1
XFILLER_7_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_044_ Inst_N_IO_ConfigMem.Inst_frame0_bit23.Q Inst_N_IO_ConfigMem.Inst_frame0_bit24.Q
+ net39 VGND VGND VPWR VPWR _023_ sky130_fd_sc_hd__or3b_1
XANTENNA_6 FrameStrobe[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput98 net115 VGND VGND VPWR VPWR B_config_C_bit3 sky130_fd_sc_hd__buf_2
Xoutput87 net104 VGND VGND VPWR VPWR A_I_top sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_2_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_292_ FrameStrobe[16] VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__clkbuf_1
XFILLER_5_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_275_ net27 VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__clkbuf_2
X_344_ Inst_N_IO_switch_matrix.SS4BEG12 VGND VGND VPWR VPWR net207 sky130_fd_sc_hd__clkbuf_1
Xoutput200 net217 VGND VGND VPWR VPWR SS4BEG[7] sky130_fd_sc_hd__buf_2
X_060_ Inst_N_IO_ConfigMem.Inst_frame0_bit31.Q VGND VGND VPWR VPWR _005_ sky130_fd_sc_hd__inv_1
X_327_ Inst_N_IO_switch_matrix.S4BEG11 VGND VGND VPWR VPWR net190 sky130_fd_sc_hd__clkbuf_1
XFILLER_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_189_ net5 net60 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame1_bit11.Q sky130_fd_sc_hd__dlxtp_1
X_258_ net8 VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_5_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_043_ _004_ _020_ _021_ Inst_N_IO_ConfigMem.Inst_frame0_bit22.Q VGND VGND VPWR VPWR
+ _022_ sky130_fd_sc_hd__a211oi_1
X_112_ net42 net81 net97 net90 Inst_N_IO_ConfigMem.Inst_frame2_bit10.Q Inst_N_IO_ConfigMem.Inst_frame2_bit11.Q
+ VGND VGND VPWR VPWR Inst_N_IO_switch_matrix.S2BEGb4 sky130_fd_sc_hd__mux4_1
XFILLER_4_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_7 FrameStrobe[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput88 net105 VGND VGND VPWR VPWR A_T_top sky130_fd_sc_hd__buf_2
Xoutput99 net116 VGND VGND VPWR VPWR FrameData_O[0] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_2_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_291_ FrameStrobe[15] VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__clkbuf_1
XFILLER_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_343_ Inst_N_IO_switch_matrix.SS4BEG11 VGND VGND VPWR VPWR net206 sky130_fd_sc_hd__clkbuf_1
X_274_ net26 VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__clkbuf_2
XFILLER_5_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput201 net218 VGND VGND VPWR VPWR SS4BEG[8] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_4_Left_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_257_ net7 VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__buf_1
X_326_ Inst_N_IO_switch_matrix.S4BEG10 VGND VGND VPWR VPWR net189 sky130_fd_sc_hd__clkbuf_1
X_188_ net4 net60 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame1_bit10.Q sky130_fd_sc_hd__dlxtp_1
X_309_ Inst_N_IO_switch_matrix.S2BEGb1 VGND VGND VPWR VPWR net181 sky130_fd_sc_hd__buf_1
X_111_ net41 net80 net96 net89 Inst_N_IO_ConfigMem.Inst_frame2_bit12.Q Inst_N_IO_ConfigMem.Inst_frame2_bit13.Q
+ VGND VGND VPWR VPWR Inst_N_IO_switch_matrix.S2BEGb5 sky130_fd_sc_hd__mux4_1
X_042_ Inst_N_IO_ConfigMem.Inst_frame0_bit23.Q Inst_N_IO_ConfigMem.Inst_frame0_bit24.Q
+ net42 VGND VGND VPWR VPWR _021_ sky130_fd_sc_hd__and3b_1
XFILLER_6_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_8 FrameStrobe[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput89 net106 VGND VGND VPWR VPWR A_config_C_bit0 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_2_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_290_ FrameStrobe[14] VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__clkbuf_1
XFILLER_4_391 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_342_ Inst_N_IO_switch_matrix.SS4BEG10 VGND VGND VPWR VPWR net205 sky130_fd_sc_hd__clkbuf_1
X_273_ net24 VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__clkbuf_2
Xoutput202 net219 VGND VGND VPWR VPWR SS4BEG[9] sky130_fd_sc_hd__buf_2
X_187_ net34 net61 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame1_bit9.Q sky130_fd_sc_hd__dlxtp_1
X_256_ net6 VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__clkbuf_1
X_325_ Inst_N_IO_switch_matrix.S4BEG9 VGND VGND VPWR VPWR net203 sky130_fd_sc_hd__clkbuf_1
XFILLER_11_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_041_ net71 net40 Inst_N_IO_ConfigMem.Inst_frame0_bit23.Q VGND VGND VPWR VPWR _020_
+ sky130_fd_sc_hd__mux2_1
X_110_ net40 net79 net95 net103 Inst_N_IO_ConfigMem.Inst_frame2_bit14.Q Inst_N_IO_ConfigMem.Inst_frame2_bit15.Q
+ VGND VGND VPWR VPWR Inst_N_IO_switch_matrix.S2BEGb6 sky130_fd_sc_hd__mux4_1
X_308_ Inst_N_IO_switch_matrix.S2BEGb0 VGND VGND VPWR VPWR net180 sky130_fd_sc_hd__clkbuf_1
X_239_ net24 net66 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame0_bit29.Q sky130_fd_sc_hd__dlxtp_1
XFILLER_4_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_9 net215 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_341_ Inst_N_IO_switch_matrix.SS4BEG9 VGND VGND VPWR VPWR net219 sky130_fd_sc_hd__clkbuf_1
X_272_ net23 VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_11_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput203 net220 VGND VGND VPWR VPWR UserCLKo sky130_fd_sc_hd__buf_1
X_186_ net33 net61 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame1_bit8.Q sky130_fd_sc_hd__dlxtp_1
X_324_ Inst_N_IO_switch_matrix.S4BEG8 VGND VGND VPWR VPWR net202 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_255_ net5 VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__clkbuf_1
XFILLER_9_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_040_ net38 net1 Inst_N_IO_ConfigMem.Inst_frame3_bit14.Q VGND VGND VPWR VPWR Inst_N_IO_switch_matrix.S1BEG0
+ sky130_fd_sc_hd__mux2_1
X_307_ Inst_N_IO_switch_matrix.S2BEG7 VGND VGND VPWR VPWR net179 sky130_fd_sc_hd__buf_1
X_169_ net18 net56 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame2_bit23.Q sky130_fd_sc_hd__dlxtp_1
X_238_ net23 net64 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame0_bit28.Q sky130_fd_sc_hd__dlxtp_1
XFILLER_8_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_11_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_340_ Inst_N_IO_switch_matrix.SS4BEG8 VGND VGND VPWR VPWR net218 sky130_fd_sc_hd__clkbuf_1
X_271_ net22 VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__clkbuf_2
X_323_ Inst_N_IO_switch_matrix.S4BEG7 VGND VGND VPWR VPWR net201 sky130_fd_sc_hd__buf_1
Xfanout60 net62 VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__buf_2
XFILLER_6_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_185_ net32 net60 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame1_bit7.Q sky130_fd_sc_hd__dlxtp_1
X_254_ net4 VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__clkbuf_1
X_099_ net35 net75 net91 Inst_B_IO_1_bidirectional_frame_config_pass.Q Inst_N_IO_ConfigMem.Inst_frame1_bit4.Q
+ Inst_N_IO_ConfigMem.Inst_frame1_bit5.Q VGND VGND VPWR VPWR Inst_N_IO_switch_matrix.S4BEG9
+ sky130_fd_sc_hd__mux4_1
XFILLER_6_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_168_ net17 net56 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame2_bit22.Q sky130_fd_sc_hd__dlxtp_1
X_306_ Inst_N_IO_switch_matrix.S2BEG6 VGND VGND VPWR VPWR net178 sky130_fd_sc_hd__clkbuf_1
X_237_ net22 net64 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame0_bit27.Q sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_270_ net21 VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__buf_1
XFILLER_4_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_322_ Inst_N_IO_switch_matrix.S4BEG6 VGND VGND VPWR VPWR net200 sky130_fd_sc_hd__clkbuf_1
Xfanout61 net62 VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__clkbuf_2
X_253_ net34 VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_9_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_184_ net31 net60 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame1_bit6.Q sky130_fd_sc_hd__dlxtp_1
XFILLER_10_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_167_ net16 net58 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame2_bit21.Q sky130_fd_sc_hd__dlxtp_1
X_305_ Inst_N_IO_switch_matrix.S2BEG5 VGND VGND VPWR VPWR net177 sky130_fd_sc_hd__clkbuf_1
X_236_ net21 net65 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame0_bit26.Q sky130_fd_sc_hd__dlxtp_1
X_098_ net87 net92 net103 Inst_A_IO_1_bidirectional_frame_config_pass.Q Inst_N_IO_ConfigMem.Inst_frame1_bit7.Q
+ Inst_N_IO_ConfigMem.Inst_frame1_bit6.Q VGND VGND VPWR VPWR Inst_N_IO_switch_matrix.S4BEG10
+ sky130_fd_sc_hd__mux4_1
X_219_ net34 net67 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame0_bit9.Q sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_11_Left_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_321_ Inst_N_IO_switch_matrix.S4BEG5 VGND VGND VPWR VPWR net199 sky130_fd_sc_hd__buf_1
X_252_ net33 VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_9_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_183_ net30 net62 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame1_bit5.Q sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_0_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout62 net63 VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__clkbuf_2
X_304_ Inst_N_IO_switch_matrix.S2BEG4 VGND VGND VPWR VPWR net176 sky130_fd_sc_hd__clkbuf_1
XFILLER_3_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_235_ net20 net64 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame0_bit25.Q sky130_fd_sc_hd__dlxtp_1
X_166_ net15 net58 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame2_bit20.Q sky130_fd_sc_hd__dlxtp_1
X_097_ net86 net91 net102 Inst_B_IO_1_bidirectional_frame_config_pass.Q Inst_N_IO_ConfigMem.Inst_frame1_bit9.Q
+ Inst_N_IO_ConfigMem.Inst_frame1_bit8.Q VGND VGND VPWR VPWR Inst_N_IO_switch_matrix.S4BEG11
+ sky130_fd_sc_hd__mux4_1
X_218_ net33 net67 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame0_bit8.Q sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_6_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_149_ net28 net59 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame2_bit3.Q sky130_fd_sc_hd__dlxtp_1
XFILLER_7_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_251_ net32 VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__buf_1
X_182_ net29 net62 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame1_bit4.Q sky130_fd_sc_hd__dlxtp_1
X_320_ Inst_N_IO_switch_matrix.S4BEG4 VGND VGND VPWR VPWR net198 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_0_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout63 FrameStrobe[1] VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__clkbuf_2
Xfanout52 net54 VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_9_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_234_ net19 net64 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame0_bit24.Q sky130_fd_sc_hd__dlxtp_1
X_165_ net13 net56 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame2_bit19.Q sky130_fd_sc_hd__dlxtp_1
X_303_ Inst_N_IO_switch_matrix.S2BEG3 VGND VGND VPWR VPWR net175 sky130_fd_sc_hd__buf_1
X_096_ net36 net99 net83 Inst_A_IO_1_bidirectional_frame_config_pass.Q Inst_N_IO_ConfigMem.Inst_frame1_bit11.Q
+ Inst_N_IO_ConfigMem.Inst_frame1_bit10.Q VGND VGND VPWR VPWR Inst_N_IO_switch_matrix.S4BEG12
+ sky130_fd_sc_hd__mux4_1
XFILLER_10_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_217_ net32 net67 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame0_bit7.Q sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_6_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_148_ net25 net59 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame2_bit2.Q sky130_fd_sc_hd__dlxtp_1
X_079_ net85 net87 net74 Inst_B_IO_1_bidirectional_frame_config_pass.Q Inst_N_IO_ConfigMem.Inst_frame0_bit12.Q
+ Inst_N_IO_ConfigMem.Inst_frame0_bit13.Q VGND VGND VPWR VPWR Inst_N_IO_switch_matrix.SS4BEG13
+ sky130_fd_sc_hd__mux4_1
XFILLER_8_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_250_ net31 VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__buf_1
XFILLER_6_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_181_ net28 net60 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame1_bit3.Q sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_0_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout64 net66 VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__clkbuf_2
Xfanout53 net54 VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__clkbuf_2
XFILLER_9_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_9_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_164_ net12 net56 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame2_bit18.Q sky130_fd_sc_hd__dlxtp_1
X_095_ net35 net98 net82 Inst_B_IO_1_bidirectional_frame_config_pass.Q Inst_N_IO_ConfigMem.Inst_frame1_bit13.Q
+ Inst_N_IO_ConfigMem.Inst_frame1_bit12.Q VGND VGND VPWR VPWR Inst_N_IO_switch_matrix.S4BEG13
+ sky130_fd_sc_hd__mux4_1
XFILLER_6_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_233_ net18 net65 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame0_bit23.Q sky130_fd_sc_hd__dlxtp_1
XFILLER_1_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_302_ Inst_N_IO_switch_matrix.S2BEG2 VGND VGND VPWR VPWR net174 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_6_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_216_ net31 net67 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame0_bit6.Q sky130_fd_sc_hd__dlxtp_1
X_147_ net14 net55 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame2_bit1.Q sky130_fd_sc_hd__dlxtp_1
X_078_ net47 net51 net49 net70 Inst_N_IO_ConfigMem.Inst_frame0_bit15.Q Inst_N_IO_ConfigMem.Inst_frame0_bit14.Q
+ VGND VGND VPWR VPWR Inst_N_IO_switch_matrix.SS4BEG14 sky130_fd_sc_hd__mux4_1
Xclkbuf_1_0__f_UserCLK_regs clknet_0_UserCLK_regs VGND VGND VPWR VPWR clknet_1_0__leaf_UserCLK_regs
+ sky130_fd_sc_hd__clkbuf_16
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout54 FrameStrobe[3] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__buf_2
X_180_ net25 net60 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame1_bit2.Q sky130_fd_sc_hd__dlxtp_1
Xfanout65 net66 VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_9_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_3_Left_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_163_ net11 net58 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame2_bit17.Q sky130_fd_sc_hd__dlxtp_1
XFILLER_10_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_301_ Inst_N_IO_switch_matrix.S2BEG1 VGND VGND VPWR VPWR net173 sky130_fd_sc_hd__buf_1
XFILLER_6_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_094_ net79 net95 net92 Inst_A_IO_1_bidirectional_frame_config_pass.Q Inst_N_IO_ConfigMem.Inst_frame1_bit14.Q
+ Inst_N_IO_ConfigMem.Inst_frame1_bit15.Q VGND VGND VPWR VPWR Inst_N_IO_switch_matrix.S4BEG14
+ sky130_fd_sc_hd__mux4_1
X_232_ net17 net64 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame0_bit22.Q sky130_fd_sc_hd__dlxtp_1
XFILLER_1_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_146_ net3 net55 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame2_bit0.Q sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_6_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_215_ net30 net68 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame0_bit5.Q sky130_fd_sc_hd__dlxtp_1
X_077_ net48 net69 net50 net71 Inst_N_IO_ConfigMem.Inst_frame0_bit17.Q Inst_N_IO_ConfigMem.Inst_frame0_bit16.Q
+ VGND VGND VPWR VPWR Inst_N_IO_switch_matrix.SS4BEG15 sky130_fd_sc_hd__mux4_1
XFILLER_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput80 NN4END[3] VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__buf_1
X_129_ net9 net54 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame3_bit15.Q sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_3_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout55 net59 VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_9_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout66 net68 VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_3_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_093_ net72 net88 net91 Inst_B_IO_1_bidirectional_frame_config_pass.Q Inst_N_IO_ConfigMem.Inst_frame1_bit16.Q
+ Inst_N_IO_ConfigMem.Inst_frame1_bit17.Q VGND VGND VPWR VPWR Inst_N_IO_switch_matrix.S4BEG15
+ sky130_fd_sc_hd__mux4_1
XFILLER_10_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_231_ net16 net64 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame0_bit21.Q sky130_fd_sc_hd__dlxtp_1
X_162_ net10 net58 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame2_bit16.Q sky130_fd_sc_hd__dlxtp_1
X_300_ Inst_N_IO_switch_matrix.S2BEG0 VGND VGND VPWR VPWR net172 sky130_fd_sc_hd__clkbuf_1
Xinput1 A_O_top VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__buf_2
X_076_ _014_ _016_ _019_ _003_ VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_6_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_145_ net27 net53 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame3_bit31.Q sky130_fd_sc_hd__dlxtp_1
X_214_ net29 net68 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame0_bit4.Q sky130_fd_sc_hd__dlxtp_1
Xclkbuf_1_0__f_UserCLK clknet_0_UserCLK VGND VGND VPWR VPWR clknet_1_0__leaf_UserCLK
+ sky130_fd_sc_hd__clkbuf_16
Xoutput190 net207 VGND VGND VPWR VPWR SS4BEG[12] sky130_fd_sc_hd__buf_2
XFILLER_11_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_128_ net8 net54 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame3_bit14.Q sky130_fd_sc_hd__dlxtp_1
X_059_ Inst_N_IO_ConfigMem.Inst_frame0_bit24.Q VGND VGND VPWR VPWR _004_ sky130_fd_sc_hd__inv_1
XFILLER_8_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput81 NN4END[4] VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_3_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput70 N4END[9] VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout56 net57 VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__clkbuf_2
Xfanout67 net68 VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_0_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_230_ net15 net65 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame0_bit20.Q sky130_fd_sc_hd__dlxtp_1
X_161_ net9 net56 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame2_bit15.Q sky130_fd_sc_hd__dlxtp_1
X_092_ net72 net80 net82 net1 Inst_N_IO_ConfigMem.Inst_frame1_bit18.Q Inst_N_IO_ConfigMem.Inst_frame1_bit19.Q
+ VGND VGND VPWR VPWR Inst_N_IO_switch_matrix.SS4BEG0 sky130_fd_sc_hd__mux4_1
Xinput2 B_O_top VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__buf_2
XFILLER_10_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_6_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_075_ _017_ _018_ Inst_N_IO_ConfigMem.Inst_frame0_bit20.Q VGND VGND VPWR VPWR _019_
+ sky130_fd_sc_hd__mux2_1
X_213_ net28 net67 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame0_bit3.Q sky130_fd_sc_hd__dlxtp_1
X_144_ net26 net53 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame3_bit30.Q sky130_fd_sc_hd__dlxtp_1
XFILLER_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput191 net208 VGND VGND VPWR VPWR SS4BEG[13] sky130_fd_sc_hd__buf_2
Xoutput180 net197 VGND VGND VPWR VPWR S4BEG[3] sky130_fd_sc_hd__buf_2
XFILLER_11_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_058_ Inst_N_IO_ConfigMem.Inst_frame0_bit21.Q VGND VGND VPWR VPWR _003_ sky130_fd_sc_hd__inv_2
X_127_ net7 net54 VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__dlxtp_1
XFILLER_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput71 NN4END[0] VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__buf_1
Xinput60 N4END[14] VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__buf_1
Xinput82 NN4END[5] VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_3_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout57 net58 VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__buf_1
XFILLER_6_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout68 FrameStrobe[0] VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__clkbuf_2
XFILLER_9_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_091_ net84 net86 net73 net2 Inst_N_IO_ConfigMem.Inst_frame1_bit20.Q Inst_N_IO_ConfigMem.Inst_frame1_bit21.Q
+ VGND VGND VPWR VPWR Inst_N_IO_switch_matrix.SS4BEG1 sky130_fd_sc_hd__mux4_1
Xclkbuf_regs_0_UserCLK UserCLK VGND VGND VPWR VPWR UserCLK_regs sky130_fd_sc_hd__clkbuf_16
X_160_ net8 net56 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame2_bit14.Q sky130_fd_sc_hd__dlxtp_1
Xinput3 FrameData[0] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_7_Left_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_289_ FrameStrobe[13] VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__clkbuf_1
XFILLER_10_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_212_ net25 net67 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame0_bit2.Q sky130_fd_sc_hd__dlxtp_1
X_143_ net24 net52 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame3_bit29.Q sky130_fd_sc_hd__dlxtp_1
X_074_ net51 net69 net70 net71 Inst_N_IO_ConfigMem.Inst_frame0_bit18.Q Inst_N_IO_ConfigMem.Inst_frame0_bit19.Q
+ VGND VGND VPWR VPWR _018_ sky130_fd_sc_hd__mux4_1
Xoutput170 net187 VGND VGND VPWR VPWR S2BEGb[7] sky130_fd_sc_hd__buf_2
Xoutput192 net209 VGND VGND VPWR VPWR SS4BEG[14] sky130_fd_sc_hd__buf_2
Xoutput181 net198 VGND VGND VPWR VPWR S4BEG[4] sky130_fd_sc_hd__buf_2
X_126_ net6 net53 VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__dlxtp_1
X_057_ Inst_N_IO_ConfigMem.Inst_frame0_bit20.Q VGND VGND VPWR VPWR _002_ sky130_fd_sc_hd__inv_1
Xinput61 N4END[15] VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__clkbuf_1
Xinput83 NN4END[6] VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__buf_1
Xinput72 NN4END[10] VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__buf_1
Xinput50 N2MID[3] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_109_ net39 net72 net88 net102 Inst_N_IO_ConfigMem.Inst_frame2_bit16.Q Inst_N_IO_ConfigMem.Inst_frame2_bit17.Q
+ VGND VGND VPWR VPWR Inst_N_IO_switch_matrix.S2BEGb7 sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_10_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout58 net59 VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_0_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_090_ net79 net81 net83 Inst_A_IO_1_bidirectional_frame_config_pass.Q Inst_N_IO_ConfigMem.Inst_frame1_bit22.Q
+ Inst_N_IO_ConfigMem.Inst_frame1_bit23.Q VGND VGND VPWR VPWR Inst_N_IO_switch_matrix.SS4BEG2
+ sky130_fd_sc_hd__mux4_1
Xclkbuf_0_UserCLK_regs UserCLK_regs VGND VGND VPWR VPWR clknet_0_UserCLK_regs sky130_fd_sc_hd__clkbuf_16
X_288_ FrameStrobe[12] VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__buf_1
Xinput4 FrameData[10] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_2
XFILLER_10_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_211_ net14 net64 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame0_bit1.Q sky130_fd_sc_hd__dlxtp_1
X_142_ net23 net54 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame3_bit28.Q sky130_fd_sc_hd__dlxtp_1
X_073_ net47 net48 net49 net50 Inst_N_IO_ConfigMem.Inst_frame0_bit18.Q Inst_N_IO_ConfigMem.Inst_frame0_bit19.Q
+ VGND VGND VPWR VPWR _017_ sky130_fd_sc_hd__mux4_1
XFILLER_2_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_125_ net5 net53 VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__dlxtp_1
Xoutput193 net210 VGND VGND VPWR VPWR SS4BEG[15] sky130_fd_sc_hd__buf_2
Xoutput182 net199 VGND VGND VPWR VPWR S4BEG[5] sky130_fd_sc_hd__buf_2
Xoutput160 net177 VGND VGND VPWR VPWR S2BEG[5] sky130_fd_sc_hd__buf_2
Xoutput171 net188 VGND VGND VPWR VPWR S4BEG[0] sky130_fd_sc_hd__buf_2
X_056_ Inst_N_IO_ConfigMem.Inst_frame0_bit28.Q VGND VGND VPWR VPWR _001_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_10_Left_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput51 N2MID[4] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_7_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput84 NN4END[7] VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__buf_1
Xinput73 NN4END[11] VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__buf_1
Xinput62 N4END[1] VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__clkbuf_2
Xinput40 N2END[1] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__buf_1
XFILLER_4_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_108_ net37 net78 net94 net1 Inst_N_IO_ConfigMem.Inst_frame2_bit18.Q Inst_N_IO_ConfigMem.Inst_frame2_bit19.Q
+ VGND VGND VPWR VPWR Inst_N_IO_switch_matrix.S4BEG0 sky130_fd_sc_hd__mux4_1
X_039_ net37 Inst_A_IO_1_bidirectional_frame_config_pass.Q Inst_N_IO_ConfigMem.Inst_frame3_bit15.Q
+ VGND VGND VPWR VPWR Inst_N_IO_switch_matrix.S1BEG1 sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_10_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout59 FrameStrobe[2] VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__clkbuf_2
XFILLER_9_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_287_ FrameStrobe[11] VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__clkbuf_1
Xinput5 FrameData[11] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_2
X_210_ net3 net64 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame0_bit0.Q sky130_fd_sc_hd__dlxtp_1
X_072_ _002_ _015_ Inst_N_IO_ConfigMem.Inst_frame0_bit21.Q VGND VGND VPWR VPWR _016_
+ sky130_fd_sc_hd__o21a_1
X_141_ net22 net53 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame3_bit27.Q sky130_fd_sc_hd__dlxtp_1
X_339_ Inst_N_IO_switch_matrix.SS4BEG7 VGND VGND VPWR VPWR net217 sky130_fd_sc_hd__buf_1
XANTENNA_10 net217 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput150 net167 VGND VGND VPWR VPWR FrameStrobe_O[9] sky130_fd_sc_hd__buf_2
X_055_ Inst_N_IO_ConfigMem.Inst_frame0_bit27.Q VGND VGND VPWR VPWR _000_ sky130_fd_sc_hd__inv_2
Xoutput194 net211 VGND VGND VPWR VPWR SS4BEG[1] sky130_fd_sc_hd__buf_2
Xoutput161 net178 VGND VGND VPWR VPWR S2BEG[6] sky130_fd_sc_hd__buf_2
Xoutput172 net189 VGND VGND VPWR VPWR S4BEG[10] sky130_fd_sc_hd__buf_2
Xoutput183 net200 VGND VGND VPWR VPWR S4BEG[6] sky130_fd_sc_hd__buf_2
X_124_ net4 net52 VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__dlxtp_1
Xinput85 NN4END[8] VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_7_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput74 NN4END[12] VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__clkbuf_2
Xinput63 N4END[2] VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput52 N2MID[5] VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput30 FrameData[5] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__clkbuf_2
Xinput41 N2END[2] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__buf_1
XFILLER_11_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_107_ net38 net77 net93 net2 Inst_N_IO_ConfigMem.Inst_frame2_bit20.Q Inst_N_IO_ConfigMem.Inst_frame2_bit21.Q
+ VGND VGND VPWR VPWR Inst_N_IO_switch_matrix.S4BEG1 sky130_fd_sc_hd__mux4_1
XFILLER_7_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_038_ net36 net2 Inst_N_IO_ConfigMem.Inst_frame3_bit16.Q VGND VGND VPWR VPWR Inst_N_IO_switch_matrix.S1BEG2
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_10_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_286_ FrameStrobe[10] VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__clkbuf_1
Xinput6 FrameData[12] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_2
XFILLER_2_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_140_ net21 net53 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame3_bit26.Q sky130_fd_sc_hd__dlxtp_1
X_071_ net43 net44 net45 net46 Inst_N_IO_ConfigMem.Inst_frame0_bit18.Q Inst_N_IO_ConfigMem.Inst_frame0_bit19.Q
+ VGND VGND VPWR VPWR _015_ sky130_fd_sc_hd__mux4_1
Xclkbuf_1_1__f_UserCLK_regs clknet_0_UserCLK_regs VGND VGND VPWR VPWR clknet_1_1__leaf_UserCLK_regs
+ sky130_fd_sc_hd__clkbuf_16
X_269_ net20 VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__clkbuf_2
X_338_ Inst_N_IO_switch_matrix.SS4BEG6 VGND VGND VPWR VPWR net216 sky130_fd_sc_hd__buf_1
Xoutput140 net157 VGND VGND VPWR VPWR FrameStrobe_O[18] sky130_fd_sc_hd__buf_2
XANTENNA_11 net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput184 net201 VGND VGND VPWR VPWR S4BEG[7] sky130_fd_sc_hd__buf_2
Xoutput162 net179 VGND VGND VPWR VPWR S2BEG[7] sky130_fd_sc_hd__buf_2
Xoutput173 net190 VGND VGND VPWR VPWR S4BEG[11] sky130_fd_sc_hd__buf_2
Xoutput195 net212 VGND VGND VPWR VPWR SS4BEG[2] sky130_fd_sc_hd__buf_2
Xoutput151 net168 VGND VGND VPWR VPWR S1BEG[0] sky130_fd_sc_hd__buf_2
XFILLER_11_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_123_ net34 net52 VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__dlxtp_1
Xinput20 FrameData[25] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_7_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput31 FrameData[6] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__clkbuf_2
X_054_ Inst_N_IO_ConfigMem.Inst_frame0_bit29.Q _029_ _030_ _031_ _028_ VGND VGND VPWR
+ VPWR net111 sky130_fd_sc_hd__a41o_1
Xinput42 N2END[3] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__buf_1
Xinput86 NN4END[9] VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__buf_1
Xinput75 NN4END[13] VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput64 N4END[3] VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__clkbuf_2
Xinput53 N2MID[6] VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__buf_1
X_037_ net35 Inst_B_IO_1_bidirectional_frame_config_pass.Q Inst_N_IO_ConfigMem.Inst_frame3_bit17.Q
+ VGND VGND VPWR VPWR Inst_N_IO_switch_matrix.S1BEG3 sky130_fd_sc_hd__mux2_1
X_106_ net74 net94 net90 net1 Inst_N_IO_ConfigMem.Inst_frame2_bit23.Q Inst_N_IO_ConfigMem.Inst_frame2_bit22.Q
+ VGND VGND VPWR VPWR Inst_N_IO_switch_matrix.S4BEG2 sky130_fd_sc_hd__mux4_1
XFILLER_8_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_285_ FrameStrobe[9] VGND VGND VPWR VPWR net167 sky130_fd_sc_hd__clkbuf_1
XFILLER_5_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput7 FrameData[13] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_2
X_070_ Inst_N_IO_ConfigMem.Inst_frame0_bit20.Q _013_ VGND VGND VPWR VPWR _014_ sky130_fd_sc_hd__or2_1
X_199_ net16 net62 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame1_bit21.Q sky130_fd_sc_hd__dlxtp_1
X_268_ net19 VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__clkbuf_2
X_337_ Inst_N_IO_switch_matrix.SS4BEG5 VGND VGND VPWR VPWR net215 sky130_fd_sc_hd__buf_1
Xoutput141 net158 VGND VGND VPWR VPWR FrameStrobe_O[19] sky130_fd_sc_hd__buf_2
Xoutput185 net202 VGND VGND VPWR VPWR S4BEG[8] sky130_fd_sc_hd__buf_2
Xoutput152 net169 VGND VGND VPWR VPWR S1BEG[1] sky130_fd_sc_hd__buf_2
Xoutput174 net191 VGND VGND VPWR VPWR S4BEG[12] sky130_fd_sc_hd__buf_2
XANTENNA_12 net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput196 net213 VGND VGND VPWR VPWR SS4BEG[3] sky130_fd_sc_hd__buf_2
Xoutput130 net147 VGND VGND VPWR VPWR FrameData_O[9] sky130_fd_sc_hd__buf_2
Xoutput163 net180 VGND VGND VPWR VPWR S2BEGb[0] sky130_fd_sc_hd__buf_2
XFILLER_11_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_122_ net33 net52 VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__dlxtp_1
XFILLER_7_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_7_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_053_ net43 Inst_N_IO_ConfigMem.Inst_frame0_bit30.Q VGND VGND VPWR VPWR _031_ sky130_fd_sc_hd__nand2_1
Xinput21 FrameData[26] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__clkbuf_2
Xinput76 NN4END[14] VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput54 N2MID[7] VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput32 FrameData[7] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__clkbuf_2
Xinput65 N4END[4] VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__clkbuf_2
Xinput10 FrameData[16] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__clkbuf_2
Xinput43 N2END[4] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__buf_1
X_105_ net73 net93 net89 net2 Inst_N_IO_ConfigMem.Inst_frame2_bit25.Q Inst_N_IO_ConfigMem.Inst_frame2_bit24.Q
+ VGND VGND VPWR VPWR Inst_N_IO_switch_matrix.S4BEG3 sky130_fd_sc_hd__mux4_1
XFILLER_4_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_036_ net71 net85 net101 net94 Inst_N_IO_ConfigMem.Inst_frame3_bit18.Q Inst_N_IO_ConfigMem.Inst_frame3_bit19.Q
+ VGND VGND VPWR VPWR Inst_N_IO_switch_matrix.S2BEG0 sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_10_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_4_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_284_ FrameStrobe[8] VGND VGND VPWR VPWR net166 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_1_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput8 FrameData[14] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_2_Left_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_198_ net15 net62 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame1_bit20.Q sky130_fd_sc_hd__dlxtp_1
X_336_ Inst_N_IO_switch_matrix.SS4BEG4 VGND VGND VPWR VPWR net214 sky130_fd_sc_hd__buf_1
X_267_ net18 VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__buf_1
Xoutput142 net159 VGND VGND VPWR VPWR FrameStrobe_O[1] sky130_fd_sc_hd__buf_2
Xoutput131 net148 VGND VGND VPWR VPWR FrameStrobe_O[0] sky130_fd_sc_hd__buf_2
Xoutput120 net137 VGND VGND VPWR VPWR FrameData_O[29] sky130_fd_sc_hd__buf_2
Xoutput175 net192 VGND VGND VPWR VPWR S4BEG[13] sky130_fd_sc_hd__buf_2
XFILLER_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_13 net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput153 net170 VGND VGND VPWR VPWR S1BEG[2] sky130_fd_sc_hd__buf_2
Xoutput197 net214 VGND VGND VPWR VPWR SS4BEG[4] sky130_fd_sc_hd__buf_2
Xoutput164 net181 VGND VGND VPWR VPWR S2BEGb[1] sky130_fd_sc_hd__buf_2
Xoutput186 net203 VGND VGND VPWR VPWR S4BEG[9] sky130_fd_sc_hd__buf_2
XFILLER_11_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_121_ net32 net52 VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__dlxtp_1
X_052_ net45 Inst_N_IO_ConfigMem.Inst_frame0_bit30.Q Inst_N_IO_ConfigMem.Inst_frame0_bit31.Q
+ VGND VGND VPWR VPWR _030_ sky130_fd_sc_hd__o21ai_1
Xinput22 FrameData[27] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__clkbuf_2
X_319_ Inst_N_IO_switch_matrix.S4BEG3 VGND VGND VPWR VPWR net197 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_7_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput11 FrameData[17] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__clkbuf_2
Xinput77 NN4END[15] VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__buf_1
Xinput66 N4END[5] VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__clkbuf_2
Xinput44 N2END[5] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput55 N4END[0] VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__clkbuf_2
Xinput33 FrameData[8] VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__clkbuf_2
XFILLER_11_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_035_ net70 net84 net100 net93 Inst_N_IO_ConfigMem.Inst_frame3_bit20.Q Inst_N_IO_ConfigMem.Inst_frame3_bit21.Q
+ VGND VGND VPWR VPWR Inst_N_IO_switch_matrix.S2BEG1 sky130_fd_sc_hd__mux4_1
X_104_ net37 net101 net85 net1 Inst_N_IO_ConfigMem.Inst_frame2_bit27.Q Inst_N_IO_ConfigMem.Inst_frame2_bit26.Q
+ VGND VGND VPWR VPWR Inst_N_IO_switch_matrix.S4BEG4 sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_10_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_283_ FrameStrobe[7] VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__buf_1
Xinput9 FrameData[15] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_2
XFILLER_5_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_1_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_197_ net13 net61 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame1_bit19.Q sky130_fd_sc_hd__dlxtp_1
X_335_ Inst_N_IO_switch_matrix.SS4BEG3 VGND VGND VPWR VPWR net213 sky130_fd_sc_hd__clkbuf_1
X_266_ net17 VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__buf_1
Xoutput132 net149 VGND VGND VPWR VPWR FrameStrobe_O[10] sky130_fd_sc_hd__buf_2
Xoutput143 net160 VGND VGND VPWR VPWR FrameStrobe_O[2] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput121 net138 VGND VGND VPWR VPWR FrameData_O[2] sky130_fd_sc_hd__buf_2
Xoutput110 net127 VGND VGND VPWR VPWR FrameData_O[1] sky130_fd_sc_hd__buf_2
XFILLER_11_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_120_ net31 net52 VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__dlxtp_1
Xoutput187 net204 VGND VGND VPWR VPWR SS4BEG[0] sky130_fd_sc_hd__buf_2
Xoutput165 net182 VGND VGND VPWR VPWR S2BEGb[2] sky130_fd_sc_hd__buf_2
X_051_ Inst_N_IO_ConfigMem.Inst_frame0_bit30.Q Inst_N_IO_ConfigMem.Inst_frame0_bit31.Q
+ net71 VGND VGND VPWR VPWR _029_ sky130_fd_sc_hd__or3b_1
Xoutput176 net193 VGND VGND VPWR VPWR S4BEG[14] sky130_fd_sc_hd__buf_2
Xoutput198 net215 VGND VGND VPWR VPWR SS4BEG[5] sky130_fd_sc_hd__buf_2
Xoutput154 net171 VGND VGND VPWR VPWR S1BEG[3] sky130_fd_sc_hd__buf_2
Xinput23 FrameData[28] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput12 FrameData[18] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput78 NN4END[1] VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_7_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput45 N2END[6] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__buf_1
X_318_ Inst_N_IO_switch_matrix.S4BEG2 VGND VGND VPWR VPWR net196 sky130_fd_sc_hd__clkbuf_1
Xinput56 N4END[10] VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput34 FrameData[9] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__clkbuf_2
Xinput67 N4END[6] VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__clkbuf_2
X_249_ net30 VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__clkbuf_2
XFILLER_4_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_103_ net38 net100 net84 net2 Inst_N_IO_ConfigMem.Inst_frame2_bit29.Q Inst_N_IO_ConfigMem.Inst_frame2_bit28.Q
+ VGND VGND VPWR VPWR Inst_N_IO_switch_matrix.S4BEG5 sky130_fd_sc_hd__mux4_1
X_034_ net69 net83 net99 net92 Inst_N_IO_ConfigMem.Inst_frame3_bit22.Q Inst_N_IO_ConfigMem.Inst_frame3_bit23.Q
+ VGND VGND VPWR VPWR Inst_N_IO_switch_matrix.S2BEG2 sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_4_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_282_ FrameStrobe[6] VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_1_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_334_ Inst_N_IO_switch_matrix.SS4BEG2 VGND VGND VPWR VPWR net212 sky130_fd_sc_hd__clkbuf_1
X_265_ net16 VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__clkbuf_2
X_196_ net12 net61 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame1_bit18.Q sky130_fd_sc_hd__dlxtp_1
Xoutput122 net139 VGND VGND VPWR VPWR FrameData_O[30] sky130_fd_sc_hd__buf_2
XFILLER_11_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput133 net150 VGND VGND VPWR VPWR FrameStrobe_O[11] sky130_fd_sc_hd__buf_2
Xoutput144 net161 VGND VGND VPWR VPWR FrameStrobe_O[3] sky130_fd_sc_hd__buf_2
XFILLER_11_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput111 net128 VGND VGND VPWR VPWR FrameData_O[20] sky130_fd_sc_hd__buf_2
XFILLER_7_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput155 net172 VGND VGND VPWR VPWR S2BEG[0] sky130_fd_sc_hd__buf_2
Xoutput166 net183 VGND VGND VPWR VPWR S2BEGb[3] sky130_fd_sc_hd__buf_2
Xoutput188 net205 VGND VGND VPWR VPWR SS4BEG[10] sky130_fd_sc_hd__buf_2
Xoutput177 net194 VGND VGND VPWR VPWR S4BEG[15] sky130_fd_sc_hd__buf_2
Xoutput199 net216 VGND VGND VPWR VPWR SS4BEG[6] sky130_fd_sc_hd__buf_2
Xoutput100 net117 VGND VGND VPWR VPWR FrameData_O[10] sky130_fd_sc_hd__buf_2
X_050_ _005_ _026_ _027_ Inst_N_IO_ConfigMem.Inst_frame0_bit29.Q VGND VGND VPWR VPWR
+ _028_ sky130_fd_sc_hd__a211oi_1
X_317_ Inst_N_IO_switch_matrix.S4BEG1 VGND VGND VPWR VPWR net195 sky130_fd_sc_hd__clkbuf_1
Xinput24 FrameData[29] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__clkbuf_2
X_248_ net29 VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__clkbuf_2
X_179_ net14 net60 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame1_bit1.Q sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_7_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput46 N2END[7] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__buf_1
Xinput13 FrameData[19] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput79 NN4END[2] VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__buf_1
Xinput68 N4END[7] VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__clkbuf_2
Xinput35 N1END[0] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__clkbuf_2
Xinput57 N4END[11] VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__buf_1
XFILLER_11_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_033_ net51 net82 net98 net91 Inst_N_IO_ConfigMem.Inst_frame3_bit24.Q Inst_N_IO_ConfigMem.Inst_frame3_bit25.Q
+ VGND VGND VPWR VPWR Inst_N_IO_switch_matrix.S2BEG3 sky130_fd_sc_hd__mux4_1
X_102_ net81 net97 net94 net1 Inst_N_IO_ConfigMem.Inst_frame2_bit30.Q Inst_N_IO_ConfigMem.Inst_frame2_bit31.Q
+ VGND VGND VPWR VPWR Inst_N_IO_switch_matrix.S4BEG6 sky130_fd_sc_hd__mux4_1
XFILLER_0_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_281_ FrameStrobe[5] VGND VGND VPWR VPWR net163 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_1_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_195_ net11 net61 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame1_bit17.Q sky130_fd_sc_hd__dlxtp_1
X_333_ Inst_N_IO_switch_matrix.SS4BEG1 VGND VGND VPWR VPWR net211 sky130_fd_sc_hd__clkbuf_1
X_264_ net15 VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__clkbuf_2
XFILLER_2_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput134 net151 VGND VGND VPWR VPWR FrameStrobe_O[12] sky130_fd_sc_hd__buf_2
Xoutput145 net162 VGND VGND VPWR VPWR FrameStrobe_O[4] sky130_fd_sc_hd__buf_2
Xoutput112 net129 VGND VGND VPWR VPWR FrameData_O[21] sky130_fd_sc_hd__buf_2
XFILLER_9_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput123 net140 VGND VGND VPWR VPWR FrameData_O[31] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_6_Left_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput156 net173 VGND VGND VPWR VPWR S2BEG[1] sky130_fd_sc_hd__buf_2
Xoutput167 net184 VGND VGND VPWR VPWR S2BEGb[4] sky130_fd_sc_hd__buf_2
Xoutput178 net195 VGND VGND VPWR VPWR S4BEG[1] sky130_fd_sc_hd__buf_2
Xoutput189 net206 VGND VGND VPWR VPWR SS4BEG[11] sky130_fd_sc_hd__buf_2
Xoutput101 net118 VGND VGND VPWR VPWR FrameData_O[11] sky130_fd_sc_hd__buf_2
XFILLER_11_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_316_ Inst_N_IO_switch_matrix.S4BEG0 VGND VGND VPWR VPWR net188 sky130_fd_sc_hd__clkbuf_1
Xinput14 FrameData[1] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__buf_1
X_247_ net28 VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__clkbuf_1
Xinput36 N1END[1] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__clkbuf_2
Xinput25 FrameData[2] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__clkbuf_2
X_178_ net3 net60 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame1_bit0.Q sky130_fd_sc_hd__dlxtp_1
XFILLER_10_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput47 N2MID[0] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__buf_1
Xinput69 N4END[8] VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput58 N4END[12] VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__buf_1
XFILLER_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_101_ net80 net96 net93 net2 Inst_N_IO_ConfigMem.Inst_frame1_bit0.Q Inst_N_IO_ConfigMem.Inst_frame1_bit1.Q
+ VGND VGND VPWR VPWR Inst_N_IO_switch_matrix.S4BEG7 sky130_fd_sc_hd__mux4_1
XFILLER_7_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_032_ net50 net81 net97 net90 Inst_N_IO_ConfigMem.Inst_frame3_bit26.Q Inst_N_IO_ConfigMem.Inst_frame3_bit27.Q
+ VGND VGND VPWR VPWR Inst_N_IO_switch_matrix.S2BEG4 sky130_fd_sc_hd__mux4_1
XFILLER_3_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_9_Left_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_280_ FrameStrobe[4] VGND VGND VPWR VPWR net162 sky130_fd_sc_hd__buf_1
XFILLER_5_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_332_ Inst_N_IO_switch_matrix.SS4BEG0 VGND VGND VPWR VPWR net204 sky130_fd_sc_hd__buf_1
X_194_ net10 net61 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame1_bit16.Q sky130_fd_sc_hd__dlxtp_1
X_263_ net13 VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__clkbuf_2
Xoutput135 net152 VGND VGND VPWR VPWR FrameStrobe_O[13] sky130_fd_sc_hd__buf_2
Xoutput146 net163 VGND VGND VPWR VPWR FrameStrobe_O[5] sky130_fd_sc_hd__buf_2
Xoutput113 net130 VGND VGND VPWR VPWR FrameData_O[22] sky130_fd_sc_hd__buf_2
Xoutput168 net185 VGND VGND VPWR VPWR S2BEGb[5] sky130_fd_sc_hd__buf_2
Xoutput124 net141 VGND VGND VPWR VPWR FrameData_O[3] sky130_fd_sc_hd__buf_2
Xoutput102 net119 VGND VGND VPWR VPWR FrameData_O[12] sky130_fd_sc_hd__buf_2
Xoutput157 net174 VGND VGND VPWR VPWR S2BEG[2] sky130_fd_sc_hd__buf_2
Xoutput179 net196 VGND VGND VPWR VPWR S4BEG[2] sky130_fd_sc_hd__buf_2
X_315_ Inst_N_IO_switch_matrix.S2BEGb7 VGND VGND VPWR VPWR net187 sky130_fd_sc_hd__buf_1
Xinput37 N1END[2] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__buf_1
Xinput26 FrameData[30] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__clkbuf_2
Xinput59 N4END[13] VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__buf_1
Xinput15 FrameData[20] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__clkbuf_2
X_246_ net25 VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__clkbuf_1
X_177_ net27 net56 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame2_bit31.Q sky130_fd_sc_hd__dlxtp_1
Xinput48 N2MID[1] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__buf_1
XFILLER_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_100_ net36 net76 net92 Inst_A_IO_1_bidirectional_frame_config_pass.Q Inst_N_IO_ConfigMem.Inst_frame1_bit2.Q
+ Inst_N_IO_ConfigMem.Inst_frame1_bit3.Q VGND VGND VPWR VPWR Inst_N_IO_switch_matrix.S4BEG8
+ sky130_fd_sc_hd__mux4_1
X_229_ net13 net65 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame0_bit19.Q sky130_fd_sc_hd__dlxtp_1
XFILLER_3_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_331_ Inst_N_IO_switch_matrix.S4BEG15 VGND VGND VPWR VPWR net194 sky130_fd_sc_hd__clkbuf_1
X_262_ net12 VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__clkbuf_2
X_193_ net9 net60 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame1_bit15.Q sky130_fd_sc_hd__dlxtp_1
Xoutput136 net153 VGND VGND VPWR VPWR FrameStrobe_O[14] sky130_fd_sc_hd__buf_2
Xoutput147 net164 VGND VGND VPWR VPWR FrameStrobe_O[6] sky130_fd_sc_hd__buf_2
Xoutput114 net131 VGND VGND VPWR VPWR FrameData_O[23] sky130_fd_sc_hd__buf_2
Xoutput103 net120 VGND VGND VPWR VPWR FrameData_O[13] sky130_fd_sc_hd__buf_2
Xoutput158 net175 VGND VGND VPWR VPWR S2BEG[3] sky130_fd_sc_hd__buf_2
Xoutput169 net186 VGND VGND VPWR VPWR S2BEGb[6] sky130_fd_sc_hd__buf_2
Xoutput125 net142 VGND VGND VPWR VPWR FrameData_O[4] sky130_fd_sc_hd__buf_2
XFILLER_11_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_245_ net14 VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__clkbuf_2
Xinput27 FrameData[31] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__clkbuf_2
XFILLER_10_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_314_ Inst_N_IO_switch_matrix.S2BEGb6 VGND VGND VPWR VPWR net186 sky130_fd_sc_hd__clkbuf_1
Xinput16 FrameData[21] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_176_ net26 net56 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame2_bit30.Q sky130_fd_sc_hd__dlxtp_1
Xinput38 N1END[3] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__clkbuf_2
Xinput49 N2MID[2] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__buf_1
XFILLER_8_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_228_ net12 net65 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame0_bit18.Q sky130_fd_sc_hd__dlxtp_1
X_159_ net7 net55 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame2_bit13.Q sky130_fd_sc_hd__dlxtp_1
XFILLER_6_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_390 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_261_ net11 VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__clkbuf_1
X_330_ Inst_N_IO_switch_matrix.S4BEG14 VGND VGND VPWR VPWR net193 sky130_fd_sc_hd__clkbuf_1
X_192_ net8 net60 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame1_bit14.Q sky130_fd_sc_hd__dlxtp_1
Xoutput115 net132 VGND VGND VPWR VPWR FrameData_O[24] sky130_fd_sc_hd__buf_2
Xoutput137 net154 VGND VGND VPWR VPWR FrameStrobe_O[15] sky130_fd_sc_hd__buf_2
Xoutput148 net165 VGND VGND VPWR VPWR FrameStrobe_O[7] sky130_fd_sc_hd__buf_2
XFILLER_9_374 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput126 net143 VGND VGND VPWR VPWR FrameData_O[5] sky130_fd_sc_hd__buf_2
Xoutput159 net176 VGND VGND VPWR VPWR S2BEG[4] sky130_fd_sc_hd__buf_2
Xoutput104 net121 VGND VGND VPWR VPWR FrameData_O[14] sky130_fd_sc_hd__buf_2
XFILLER_11_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_244_ net3 VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__clkbuf_2
Xinput17 FrameData[22] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__clkbuf_2
X_175_ net24 net56 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame2_bit29.Q sky130_fd_sc_hd__dlxtp_1
XFILLER_6_388 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_313_ Inst_N_IO_switch_matrix.S2BEGb5 VGND VGND VPWR VPWR net185 sky130_fd_sc_hd__clkbuf_1
Xinput39 N2END[0] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__clkbuf_2
Xinput28 FrameData[3] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__clkbuf_2
XFILLER_11_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_089_ net85 net87 net74 Inst_B_IO_1_bidirectional_frame_config_pass.Q Inst_N_IO_ConfigMem.Inst_frame1_bit24.Q
+ Inst_N_IO_ConfigMem.Inst_frame1_bit25.Q VGND VGND VPWR VPWR Inst_N_IO_switch_matrix.SS4BEG3
+ sky130_fd_sc_hd__mux4_1
X_158_ net6 net55 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame2_bit12.Q sky130_fd_sc_hd__dlxtp_1
X_227_ net11 net68 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame0_bit17.Q sky130_fd_sc_hd__dlxtp_1
XFILLER_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_260_ net10 VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__clkbuf_1
XFILLER_9_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_191_ net7 net61 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame1_bit13.Q sky130_fd_sc_hd__dlxtp_1
XFILLER_2_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput116 net133 VGND VGND VPWR VPWR FrameData_O[25] sky130_fd_sc_hd__buf_2
Xoutput138 net155 VGND VGND VPWR VPWR FrameStrobe_O[16] sky130_fd_sc_hd__buf_2
Xoutput149 net166 VGND VGND VPWR VPWR FrameStrobe_O[8] sky130_fd_sc_hd__buf_2
Xoutput105 net122 VGND VGND VPWR VPWR FrameData_O[15] sky130_fd_sc_hd__buf_2
Xoutput127 net144 VGND VGND VPWR VPWR FrameData_O[6] sky130_fd_sc_hd__buf_2
XFILLER_10_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput18 FrameData[23] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__clkbuf_2
X_174_ net23 net57 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame2_bit28.Q sky130_fd_sc_hd__dlxtp_1
X_243_ clknet_1_1__leaf_UserCLK_regs net2 VGND VGND VPWR VPWR Inst_B_IO_1_bidirectional_frame_config_pass.Q
+ sky130_fd_sc_hd__dfxtp_1
X_312_ Inst_N_IO_switch_matrix.S2BEGb4 VGND VGND VPWR VPWR net184 sky130_fd_sc_hd__clkbuf_1
Xinput29 FrameData[4] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__clkbuf_2
X_088_ net39 net41 net43 net45 Inst_N_IO_ConfigMem.Inst_frame1_bit26.Q Inst_N_IO_ConfigMem.Inst_frame1_bit27.Q
+ VGND VGND VPWR VPWR Inst_N_IO_switch_matrix.SS4BEG4 sky130_fd_sc_hd__mux4_1
X_157_ net5 net55 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame2_bit11.Q sky130_fd_sc_hd__dlxtp_1
X_226_ net10 net68 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame0_bit16.Q sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_8_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_209_ net27 net63 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame1_bit31.Q sky130_fd_sc_hd__dlxtp_1
XFILLER_8_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_1_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_190_ net6 net61 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame1_bit12.Q sky130_fd_sc_hd__dlxtp_1
Xoutput139 net156 VGND VGND VPWR VPWR FrameStrobe_O[17] sky130_fd_sc_hd__buf_2
Xoutput117 net134 VGND VGND VPWR VPWR FrameData_O[26] sky130_fd_sc_hd__buf_2
Xoutput106 net123 VGND VGND VPWR VPWR FrameData_O[16] sky130_fd_sc_hd__buf_2
Xoutput128 net145 VGND VGND VPWR VPWR FrameData_O[7] sky130_fd_sc_hd__buf_2
XFILLER_10_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput19 FrameData[24] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__clkbuf_2
X_311_ Inst_N_IO_switch_matrix.S2BEGb3 VGND VGND VPWR VPWR net183 sky130_fd_sc_hd__buf_1
X_173_ net22 net57 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame2_bit27.Q sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_1_Left_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_242_ clknet_1_0__leaf_UserCLK_regs net1 VGND VGND VPWR VPWR Inst_A_IO_1_bidirectional_frame_config_pass.Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_5_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_225_ net9 net64 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame0_bit15.Q sky130_fd_sc_hd__dlxtp_1
X_156_ net4 net55 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame2_bit10.Q sky130_fd_sc_hd__dlxtp_1
X_087_ net40 net42 net44 net46 Inst_N_IO_ConfigMem.Inst_frame1_bit28.Q Inst_N_IO_ConfigMem.Inst_frame1_bit29.Q
+ VGND VGND VPWR VPWR Inst_N_IO_switch_matrix.SS4BEG5 sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_8_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_139_ net20 net52 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame3_bit25.Q sky130_fd_sc_hd__dlxtp_1
X_208_ net26 net63 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame1_bit30.Q sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_5_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput118 net135 VGND VGND VPWR VPWR FrameData_O[27] sky130_fd_sc_hd__buf_2
Xoutput107 net124 VGND VGND VPWR VPWR FrameData_O[17] sky130_fd_sc_hd__buf_2
Xoutput129 net146 VGND VGND VPWR VPWR FrameData_O[8] sky130_fd_sc_hd__buf_2
X_310_ Inst_N_IO_switch_matrix.S2BEGb2 VGND VGND VPWR VPWR net182 sky130_fd_sc_hd__clkbuf_1
X_241_ net27 net66 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame0_bit31.Q sky130_fd_sc_hd__dlxtp_1
X_172_ net21 net57 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame2_bit26.Q sky130_fd_sc_hd__dlxtp_1
XFILLER_9_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_155_ net34 net55 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame2_bit9.Q sky130_fd_sc_hd__dlxtp_1
X_224_ net8 net64 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame0_bit14.Q sky130_fd_sc_hd__dlxtp_1
X_086_ net47 net51 net49 net70 Inst_N_IO_ConfigMem.Inst_frame1_bit31.Q Inst_N_IO_ConfigMem.Inst_frame1_bit30.Q
+ VGND VGND VPWR VPWR Inst_N_IO_switch_matrix.SS4BEG6 sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_8_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_069_ net39 net40 net41 net42 Inst_N_IO_ConfigMem.Inst_frame0_bit18.Q Inst_N_IO_ConfigMem.Inst_frame0_bit19.Q
+ VGND VGND VPWR VPWR _013_ sky130_fd_sc_hd__mux4_1
X_138_ net19 net52 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame3_bit24.Q sky130_fd_sc_hd__dlxtp_1
X_207_ net24 net63 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame1_bit29.Q sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput90 net107 VGND VGND VPWR VPWR A_config_C_bit1 sky130_fd_sc_hd__buf_2
Xoutput119 net136 VGND VGND VPWR VPWR FrameData_O[28] sky130_fd_sc_hd__buf_2
Xoutput108 net125 VGND VGND VPWR VPWR FrameData_O[18] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_2_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_171_ net20 net57 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame2_bit25.Q sky130_fd_sc_hd__dlxtp_1
X_240_ net26 net66 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame0_bit30.Q sky130_fd_sc_hd__dlxtp_1
XFILLER_11_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_223_ net7 net67 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame0_bit13.Q sky130_fd_sc_hd__dlxtp_1
X_154_ net33 net55 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame2_bit8.Q sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_8_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_085_ net48 net69 net50 net71 Inst_N_IO_ConfigMem.Inst_frame0_bit1.Q Inst_N_IO_ConfigMem.Inst_frame0_bit0.Q
+ VGND VGND VPWR VPWR Inst_N_IO_switch_matrix.SS4BEG7 sky130_fd_sc_hd__mux4_1
XFILLER_2_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_137_ net18 net53 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame3_bit23.Q sky130_fd_sc_hd__dlxtp_1
X_068_ _007_ _009_ _012_ _001_ VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__a22o_1
X_206_ net23 net63 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame1_bit28.Q sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_5_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput109 net126 VGND VGND VPWR VPWR FrameData_O[19] sky130_fd_sc_hd__buf_2
XFILLER_1_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput91 net108 VGND VGND VPWR VPWR A_config_C_bit2 sky130_fd_sc_hd__buf_2
XFILLER_11_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_170_ net19 net57 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame2_bit24.Q sky130_fd_sc_hd__dlxtp_1
X_299_ Inst_N_IO_switch_matrix.S1BEG3 VGND VGND VPWR VPWR net171 sky130_fd_sc_hd__buf_1
XFILLER_5_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_5_Left_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_084_ net82 net86 net84 net73 Inst_N_IO_ConfigMem.Inst_frame0_bit3.Q Inst_N_IO_ConfigMem.Inst_frame0_bit2.Q
+ VGND VGND VPWR VPWR Inst_N_IO_switch_matrix.SS4BEG8 sky130_fd_sc_hd__mux4_1
X_222_ net6 net67 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame0_bit12.Q sky130_fd_sc_hd__dlxtp_1
X_153_ net32 net59 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame2_bit7.Q sky130_fd_sc_hd__dlxtp_1
X_205_ net22 net63 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame1_bit27.Q sky130_fd_sc_hd__dlxtp_1
X_136_ net17 net53 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame3_bit22.Q sky130_fd_sc_hd__dlxtp_1
XFILLER_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_067_ _010_ _011_ _000_ VGND VGND VPWR VPWR _012_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_8_Left_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_119_ net49 net80 net96 net89 Inst_N_IO_ConfigMem.Inst_frame3_bit28.Q Inst_N_IO_ConfigMem.Inst_frame3_bit29.Q
+ VGND VGND VPWR VPWR Inst_N_IO_switch_matrix.S2BEG5 sky130_fd_sc_hd__mux4_1
XFILLER_9_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput92 net109 VGND VGND VPWR VPWR A_config_C_bit3 sky130_fd_sc_hd__buf_2
XFILLER_8_380 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_9_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_298_ Inst_N_IO_switch_matrix.S1BEG2 VGND VGND VPWR VPWR net170 sky130_fd_sc_hd__buf_1
X_152_ net31 net59 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame2_bit6.Q sky130_fd_sc_hd__dlxtp_1
X_221_ net5 net67 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame0_bit11.Q sky130_fd_sc_hd__dlxtp_1
X_083_ net79 net81 net83 net85 Inst_N_IO_ConfigMem.Inst_frame0_bit4.Q Inst_N_IO_ConfigMem.Inst_frame0_bit5.Q
+ VGND VGND VPWR VPWR Inst_N_IO_switch_matrix.SS4BEG9 sky130_fd_sc_hd__mux4_1
X_204_ net21 net63 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame1_bit26.Q sky130_fd_sc_hd__dlxtp_1
X_135_ net16 net52 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame3_bit21.Q sky130_fd_sc_hd__dlxtp_1
XFILLER_7_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_066_ net47 net48 net49 net50 Inst_N_IO_ConfigMem.Inst_frame0_bit25.Q Inst_N_IO_ConfigMem.Inst_frame0_bit26.Q
+ VGND VGND VPWR VPWR _011_ sky130_fd_sc_hd__mux4_1
XFILLER_8_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_118_ net48 net79 net95 net103 Inst_N_IO_ConfigMem.Inst_frame3_bit30.Q Inst_N_IO_ConfigMem.Inst_frame3_bit31.Q
+ VGND VGND VPWR VPWR Inst_N_IO_switch_matrix.S2BEG6 sky130_fd_sc_hd__mux4_1
X_049_ Inst_N_IO_ConfigMem.Inst_frame0_bit30.Q Inst_N_IO_ConfigMem.Inst_frame0_bit31.Q
+ net44 VGND VGND VPWR VPWR _027_ sky130_fd_sc_hd__and3b_1
XANTENNA_1 net129 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput93 net110 VGND VGND VPWR VPWR B_I_top sky130_fd_sc_hd__buf_2
XFILLER_8_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_297_ Inst_N_IO_switch_matrix.S1BEG1 VGND VGND VPWR VPWR net169 sky130_fd_sc_hd__clkbuf_1
X_082_ net72 net80 net82 net1 Inst_N_IO_ConfigMem.Inst_frame0_bit6.Q Inst_N_IO_ConfigMem.Inst_frame0_bit7.Q
+ VGND VGND VPWR VPWR Inst_N_IO_switch_matrix.SS4BEG10 sky130_fd_sc_hd__mux4_1
XFILLER_10_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_151_ net30 net55 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame2_bit5.Q sky130_fd_sc_hd__dlxtp_1
X_220_ net4 net67 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame0_bit10.Q sky130_fd_sc_hd__dlxtp_1
X_134_ net15 net52 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame3_bit20.Q sky130_fd_sc_hd__dlxtp_1
X_203_ net20 net61 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame1_bit25.Q sky130_fd_sc_hd__dlxtp_1
XFILLER_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_065_ net51 net69 net70 net71 Inst_N_IO_ConfigMem.Inst_frame0_bit25.Q Inst_N_IO_ConfigMem.Inst_frame0_bit26.Q
+ VGND VGND VPWR VPWR _010_ sky130_fd_sc_hd__mux4_1
XFILLER_9_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_UserCLK UserCLK VGND VGND VPWR VPWR clknet_0_UserCLK sky130_fd_sc_hd__clkbuf_16
X_117_ net47 net72 net88 net102 Inst_N_IO_ConfigMem.Inst_frame2_bit0.Q Inst_N_IO_ConfigMem.Inst_frame2_bit1.Q
+ VGND VGND VPWR VPWR Inst_N_IO_switch_matrix.S2BEG7 sky130_fd_sc_hd__mux4_1
X_048_ net70 net39 Inst_N_IO_ConfigMem.Inst_frame0_bit30.Q VGND VGND VPWR VPWR _026_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_2 net130 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput94 net111 VGND VGND VPWR VPWR B_T_top sky130_fd_sc_hd__buf_2
XFILLER_9_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_296_ Inst_N_IO_switch_matrix.S1BEG0 VGND VGND VPWR VPWR net168 sky130_fd_sc_hd__buf_1
X_150_ net29 net55 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame2_bit4.Q sky130_fd_sc_hd__dlxtp_1
X_081_ net84 net86 net73 net2 Inst_N_IO_ConfigMem.Inst_frame0_bit8.Q Inst_N_IO_ConfigMem.Inst_frame0_bit9.Q
+ VGND VGND VPWR VPWR Inst_N_IO_switch_matrix.SS4BEG11 sky130_fd_sc_hd__mux4_1
X_348_ clknet_1_0__leaf_UserCLK VGND VGND VPWR VPWR net220 sky130_fd_sc_hd__buf_2
X_279_ net54 VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__buf_1
X_202_ net19 net61 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame1_bit24.Q sky130_fd_sc_hd__dlxtp_1
X_133_ net13 net53 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame3_bit19.Q sky130_fd_sc_hd__dlxtp_1
X_064_ _000_ _008_ Inst_N_IO_ConfigMem.Inst_frame0_bit28.Q VGND VGND VPWR VPWR _009_
+ sky130_fd_sc_hd__o21a_1
X_116_ net46 net85 net101 net94 Inst_N_IO_ConfigMem.Inst_frame2_bit2.Q Inst_N_IO_ConfigMem.Inst_frame2_bit3.Q
+ VGND VGND VPWR VPWR Inst_N_IO_switch_matrix.S2BEGb0 sky130_fd_sc_hd__mux4_1
X_047_ Inst_N_IO_ConfigMem.Inst_frame0_bit22.Q _023_ _024_ _025_ _022_ VGND VGND VPWR
+ VPWR net105 sky130_fd_sc_hd__a41o_1
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_3 net131 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput95 net112 VGND VGND VPWR VPWR B_config_C_bit0 sky130_fd_sc_hd__buf_2
XFILLER_0_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_295_ FrameStrobe[19] VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__clkbuf_1
X_080_ net79 net81 net83 Inst_A_IO_1_bidirectional_frame_config_pass.Q Inst_N_IO_ConfigMem.Inst_frame0_bit10.Q
+ Inst_N_IO_ConfigMem.Inst_frame0_bit11.Q VGND VGND VPWR VPWR Inst_N_IO_switch_matrix.SS4BEG12
+ sky130_fd_sc_hd__mux4_1
X_278_ net56 VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_8_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_347_ Inst_N_IO_switch_matrix.SS4BEG15 VGND VGND VPWR VPWR net210 sky130_fd_sc_hd__buf_1
X_132_ net12 net53 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame3_bit18.Q sky130_fd_sc_hd__dlxtp_1
XFILLER_2_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_201_ net18 net62 VGND VGND VPWR VPWR Inst_N_IO_ConfigMem.Inst_frame1_bit23.Q sky130_fd_sc_hd__dlxtp_1
X_063_ net43 net44 net45 net46 Inst_N_IO_ConfigMem.Inst_frame0_bit25.Q Inst_N_IO_ConfigMem.Inst_frame0_bit26.Q
+ VGND VGND VPWR VPWR _008_ sky130_fd_sc_hd__mux4_1
XFILLER_9_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_115_ net45 net84 net100 net93 Inst_N_IO_ConfigMem.Inst_frame2_bit4.Q Inst_N_IO_ConfigMem.Inst_frame2_bit5.Q
+ VGND VGND VPWR VPWR Inst_N_IO_switch_matrix.S2BEGb1 sky130_fd_sc_hd__mux4_1
X_046_ net41 Inst_N_IO_ConfigMem.Inst_frame0_bit23.Q VGND VGND VPWR VPWR _025_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_5_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_4 net139 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput96 net113 VGND VGND VPWR VPWR B_config_C_bit1 sky130_fd_sc_hd__buf_2
.ends

