* NGSPICE file created from N_term_single.ext - technology: sky130A

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

.subckt N_term_single Ci FrameData[0] FrameData[10] FrameData[11] FrameData[12] FrameData[13]
+ FrameData[14] FrameData[15] FrameData[16] FrameData[17] FrameData[18] FrameData[19]
+ FrameData[1] FrameData[20] FrameData[21] FrameData[22] FrameData[23] FrameData[24]
+ FrameData[25] FrameData[26] FrameData[27] FrameData[28] FrameData[29] FrameData[2]
+ FrameData[30] FrameData[31] FrameData[3] FrameData[4] FrameData[5] FrameData[6]
+ FrameData[7] FrameData[8] FrameData[9] FrameData_O[0] FrameData_O[10] FrameData_O[11]
+ FrameData_O[12] FrameData_O[13] FrameData_O[14] FrameData_O[15] FrameData_O[16]
+ FrameData_O[17] FrameData_O[18] FrameData_O[19] FrameData_O[1] FrameData_O[20] FrameData_O[21]
+ FrameData_O[22] FrameData_O[23] FrameData_O[24] FrameData_O[25] FrameData_O[26]
+ FrameData_O[27] FrameData_O[28] FrameData_O[29] FrameData_O[2] FrameData_O[30] FrameData_O[31]
+ FrameData_O[3] FrameData_O[4] FrameData_O[5] FrameData_O[6] FrameData_O[7] FrameData_O[8]
+ FrameData_O[9] FrameStrobe[0] FrameStrobe[10] FrameStrobe[11] FrameStrobe[12] FrameStrobe[13]
+ FrameStrobe[14] FrameStrobe[15] FrameStrobe[16] FrameStrobe[17] FrameStrobe[18]
+ FrameStrobe[19] FrameStrobe[1] FrameStrobe[2] FrameStrobe[3] FrameStrobe[4] FrameStrobe[5]
+ FrameStrobe[6] FrameStrobe[7] FrameStrobe[8] FrameStrobe[9] FrameStrobe_O[0] FrameStrobe_O[10]
+ FrameStrobe_O[11] FrameStrobe_O[12] FrameStrobe_O[13] FrameStrobe_O[14] FrameStrobe_O[15]
+ FrameStrobe_O[16] FrameStrobe_O[17] FrameStrobe_O[18] FrameStrobe_O[19] FrameStrobe_O[1]
+ FrameStrobe_O[2] FrameStrobe_O[3] FrameStrobe_O[4] FrameStrobe_O[5] FrameStrobe_O[6]
+ FrameStrobe_O[7] FrameStrobe_O[8] FrameStrobe_O[9] N1END[0] N1END[1] N1END[2] N1END[3]
+ N2END[0] N2END[1] N2END[2] N2END[3] N2END[4] N2END[5] N2END[6] N2END[7] N2MID[0]
+ N2MID[1] N2MID[2] N2MID[3] N2MID[4] N2MID[5] N2MID[6] N2MID[7] N4END[0] N4END[10]
+ N4END[11] N4END[12] N4END[13] N4END[14] N4END[15] N4END[1] N4END[2] N4END[3] N4END[4]
+ N4END[5] N4END[6] N4END[7] N4END[8] N4END[9] NN4END[0] NN4END[10] NN4END[11] NN4END[12]
+ NN4END[13] NN4END[14] NN4END[15] NN4END[1] NN4END[2] NN4END[3] NN4END[4] NN4END[5]
+ NN4END[6] NN4END[7] NN4END[8] NN4END[9] S1BEG[0] S1BEG[1] S1BEG[2] S1BEG[3] S2BEG[0]
+ S2BEG[1] S2BEG[2] S2BEG[3] S2BEG[4] S2BEG[5] S2BEG[6] S2BEG[7] S2BEGb[0] S2BEGb[1]
+ S2BEGb[2] S2BEGb[3] S2BEGb[4] S2BEGb[5] S2BEGb[6] S2BEGb[7] S4BEG[0] S4BEG[10] S4BEG[11]
+ S4BEG[12] S4BEG[13] S4BEG[14] S4BEG[15] S4BEG[1] S4BEG[2] S4BEG[3] S4BEG[4] S4BEG[5]
+ S4BEG[6] S4BEG[7] S4BEG[8] S4BEG[9] SS4BEG[0] SS4BEG[10] SS4BEG[11] SS4BEG[12] SS4BEG[13]
+ SS4BEG[14] SS4BEG[15] SS4BEG[1] SS4BEG[2] SS4BEG[3] SS4BEG[4] SS4BEG[5] SS4BEG[6]
+ SS4BEG[7] SS4BEG[8] SS4BEG[9] UserCLK UserCLKo VGND VPWR
XFILLER_9_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_0_Left_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_11_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_062_ N2MID[1] VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__buf_1
XFILLER_7_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_045_ FrameStrobe[13] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__clkbuf_1
XFILLER_4_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_028_ FrameData[28] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__buf_1
XFILLER_6_89 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_5 FrameData[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput42 net42 VGND VGND VPWR VPWR FrameStrobe_O[18] sky130_fd_sc_hd__buf_2
Xoutput20 net20 VGND VGND VPWR VPWR FrameData_O[27] sky130_fd_sc_hd__buf_2
XFILLER_8_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput7 net7 VGND VGND VPWR VPWR FrameData_O[15] sky130_fd_sc_hd__buf_2
Xoutput64 net64 VGND VGND VPWR VPWR S2BEG[7] sky130_fd_sc_hd__buf_2
Xoutput53 net53 VGND VGND VPWR VPWR S1BEG[0] sky130_fd_sc_hd__buf_2
Xoutput86 net86 VGND VGND VPWR VPWR S4BEG[7] sky130_fd_sc_hd__buf_2
Xoutput75 net75 VGND VGND VPWR VPWR S4BEG[11] sky130_fd_sc_hd__buf_2
Xoutput97 net97 VGND VGND VPWR VPWR SS4BEG[2] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_2_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput31 net31 VGND VGND VPWR VPWR FrameData_O[8] sky130_fd_sc_hd__buf_2
XFILLER_10_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_11_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_196 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_061_ N2MID[2] VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__buf_1
XFILLER_0_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_044_ FrameStrobe[12] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__clkbuf_1
XFILLER_7_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_027_ FrameData[27] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__buf_1
XFILLER_3_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_6 FrameData[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput43 net43 VGND VGND VPWR VPWR FrameStrobe_O[19] sky130_fd_sc_hd__buf_2
Xoutput21 net21 VGND VGND VPWR VPWR FrameData_O[28] sky130_fd_sc_hd__buf_2
Xoutput8 net8 VGND VGND VPWR VPWR FrameData_O[16] sky130_fd_sc_hd__buf_2
Xoutput10 net10 VGND VGND VPWR VPWR FrameData_O[18] sky130_fd_sc_hd__buf_2
Xoutput65 net65 VGND VGND VPWR VPWR S2BEGb[0] sky130_fd_sc_hd__buf_2
Xoutput54 net54 VGND VGND VPWR VPWR S1BEG[1] sky130_fd_sc_hd__buf_2
Xoutput87 net87 VGND VGND VPWR VPWR S4BEG[8] sky130_fd_sc_hd__buf_2
Xoutput76 net76 VGND VGND VPWR VPWR S4BEG[12] sky130_fd_sc_hd__buf_2
Xoutput98 net98 VGND VGND VPWR VPWR SS4BEG[3] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_2_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput32 net32 VGND VGND VPWR VPWR FrameData_O[9] sky130_fd_sc_hd__buf_2
XFILLER_8_183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_060_ N2MID[3] VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__buf_1
XFILLER_0_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_043_ FrameStrobe[11] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__clkbuf_1
XFILLER_7_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_026_ FrameData[26] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__buf_1
XFILLER_6_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_7 FrameData[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput44 net44 VGND VGND VPWR VPWR FrameStrobe_O[1] sky130_fd_sc_hd__buf_2
Xoutput33 net33 VGND VGND VPWR VPWR FrameStrobe_O[0] sky130_fd_sc_hd__buf_2
Xoutput22 net22 VGND VGND VPWR VPWR FrameData_O[29] sky130_fd_sc_hd__buf_2
Xoutput11 net11 VGND VGND VPWR VPWR FrameData_O[19] sky130_fd_sc_hd__buf_2
Xoutput9 net9 VGND VGND VPWR VPWR FrameData_O[17] sky130_fd_sc_hd__buf_2
Xoutput66 net66 VGND VGND VPWR VPWR S2BEGb[1] sky130_fd_sc_hd__buf_2
Xoutput55 net55 VGND VGND VPWR VPWR S1BEG[2] sky130_fd_sc_hd__buf_2
Xoutput88 net88 VGND VGND VPWR VPWR S4BEG[9] sky130_fd_sc_hd__buf_2
Xoutput77 net77 VGND VGND VPWR VPWR S4BEG[13] sky130_fd_sc_hd__buf_2
Xoutput99 net99 VGND VGND VPWR VPWR SS4BEG[4] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_2_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_009_ FrameData[9] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__buf_1
XFILLER_10_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_4_Left_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_042_ FrameStrobe[10] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__clkbuf_1
XFILLER_7_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_025_ FrameData[25] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__buf_1
XANTENNA_8 FrameData[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput34 net34 VGND VGND VPWR VPWR FrameStrobe_O[10] sky130_fd_sc_hd__buf_2
Xoutput45 net45 VGND VGND VPWR VPWR FrameStrobe_O[2] sky130_fd_sc_hd__buf_2
Xoutput67 net67 VGND VGND VPWR VPWR S2BEGb[2] sky130_fd_sc_hd__buf_2
Xoutput56 net56 VGND VGND VPWR VPWR S1BEG[3] sky130_fd_sc_hd__buf_2
XFILLER_0_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput78 net78 VGND VGND VPWR VPWR S4BEG[14] sky130_fd_sc_hd__buf_2
Xoutput89 net89 VGND VGND VPWR VPWR SS4BEG[0] sky130_fd_sc_hd__buf_2
Xoutput12 net12 VGND VGND VPWR VPWR FrameData_O[1] sky130_fd_sc_hd__buf_2
Xoutput23 net23 VGND VGND VPWR VPWR FrameData_O[2] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_2_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_008_ FrameData[8] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__buf_1
XFILLER_3_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_391 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_041_ FrameStrobe[9] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__clkbuf_1
XFILLER_7_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_024_ FrameData[24] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__buf_1
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_9 FrameData[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput24 net24 VGND VGND VPWR VPWR FrameData_O[30] sky130_fd_sc_hd__buf_2
Xoutput35 net35 VGND VGND VPWR VPWR FrameStrobe_O[11] sky130_fd_sc_hd__buf_2
Xoutput46 net46 VGND VGND VPWR VPWR FrameStrobe_O[3] sky130_fd_sc_hd__buf_2
Xoutput13 net13 VGND VGND VPWR VPWR FrameData_O[20] sky130_fd_sc_hd__buf_2
Xoutput57 net57 VGND VGND VPWR VPWR S2BEG[0] sky130_fd_sc_hd__buf_2
XFILLER_8_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput68 net68 VGND VGND VPWR VPWR S2BEGb[3] sky130_fd_sc_hd__buf_2
XFILLER_0_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput79 net79 VGND VGND VPWR VPWR S4BEG[15] sky130_fd_sc_hd__buf_2
X_007_ FrameData[7] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__buf_1
XFILLER_7_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_236 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_040_ FrameStrobe[8] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__clkbuf_1
XFILLER_1_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_023_ FrameData[23] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__buf_1
Xoutput36 net36 VGND VGND VPWR VPWR FrameStrobe_O[12] sky130_fd_sc_hd__buf_2
Xoutput47 net47 VGND VGND VPWR VPWR FrameStrobe_O[4] sky130_fd_sc_hd__buf_2
Xoutput25 net25 VGND VGND VPWR VPWR FrameData_O[31] sky130_fd_sc_hd__buf_2
Xoutput14 net14 VGND VGND VPWR VPWR FrameData_O[21] sky130_fd_sc_hd__buf_2
XFILLER_8_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput69 net69 VGND VGND VPWR VPWR S2BEGb[4] sky130_fd_sc_hd__buf_2
Xoutput58 net58 VGND VGND VPWR VPWR S2BEG[1] sky130_fd_sc_hd__buf_2
X_006_ FrameData[6] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__buf_1
XFILLER_5_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_099_ NN4END[4] VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__clkbuf_1
XFILLER_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_022_ FrameData[22] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__buf_1
XFILLER_6_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput37 net37 VGND VGND VPWR VPWR FrameStrobe_O[13] sky130_fd_sc_hd__buf_2
Xoutput48 net48 VGND VGND VPWR VPWR FrameStrobe_O[5] sky130_fd_sc_hd__buf_2
Xoutput15 net15 VGND VGND VPWR VPWR FrameData_O[22] sky130_fd_sc_hd__buf_2
Xoutput59 net59 VGND VGND VPWR VPWR S2BEG[2] sky130_fd_sc_hd__buf_2
Xoutput26 net26 VGND VGND VPWR VPWR FrameData_O[3] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_005_ FrameData[5] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__buf_1
XFILLER_7_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_275 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_098_ NN4END[5] VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__clkbuf_1
XFILLER_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_021_ FrameData[21] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__buf_1
XFILLER_3_234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_256 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_11_Left_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput38 net38 VGND VGND VPWR VPWR FrameStrobe_O[14] sky130_fd_sc_hd__buf_2
Xoutput49 net49 VGND VGND VPWR VPWR FrameStrobe_O[6] sky130_fd_sc_hd__buf_2
Xoutput16 net16 VGND VGND VPWR VPWR FrameData_O[23] sky130_fd_sc_hd__buf_2
Xoutput27 net27 VGND VGND VPWR VPWR FrameData_O[4] sky130_fd_sc_hd__buf_2
X_004_ FrameData[4] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__buf_1
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_3_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_351 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_287 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_097_ NN4END[6] VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__clkbuf_1
X_020_ FrameData[20] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__buf_1
XFILLER_3_202 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput17 net17 VGND VGND VPWR VPWR FrameData_O[24] sky130_fd_sc_hd__buf_2
Xoutput39 net39 VGND VGND VPWR VPWR FrameStrobe_O[15] sky130_fd_sc_hd__buf_2
XFILLER_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput28 net28 VGND VGND VPWR VPWR FrameData_O[5] sky130_fd_sc_hd__buf_2
X_003_ FrameData[3] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__buf_1
XFILLER_7_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_171 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_096_ NN4END[7] VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__clkbuf_1
XFILLER_10_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput18 net18 VGND VGND VPWR VPWR FrameData_O[25] sky130_fd_sc_hd__buf_2
X_079_ N4END[8] VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__buf_1
Xoutput29 net29 VGND VGND VPWR VPWR FrameData_O[6] sky130_fd_sc_hd__buf_2
XFILLER_2_291 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_002_ FrameData[2] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__buf_1
XFILLER_7_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_54 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_095_ NN4END[8] VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__clkbuf_1
XFILLER_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_078_ N4END[9] VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__buf_1
Xoutput19 net19 VGND VGND VPWR VPWR FrameData_O[26] sky130_fd_sc_hd__buf_2
XFILLER_8_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_001_ FrameData[1] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__buf_1
XFILLER_7_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_87 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_3_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_66 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_3_Left_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_094_ NN4END[9] VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__clkbuf_1
XFILLER_10_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_077_ N4END[10] VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__buf_1
XFILLER_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_000_ FrameData[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__buf_1
XFILLER_7_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_99 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_3_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_093_ NN4END[10] VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__clkbuf_1
XFILLER_1_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_076_ N4END[11] VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__buf_1
XFILLER_8_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_059_ N2MID[4] VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_3_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_092_ NN4END[11] VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__clkbuf_1
XFILLER_5_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_6_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_075_ N4END[12] VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__buf_1
XANTENNA_40 NN4END[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_058_ N2MID[5] VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__buf_1
XFILLER_8_118 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_379 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_091_ NN4END[12] VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_7_Left_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_074_ N4END[13] VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__buf_1
XANTENNA_30 FrameStrobe[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_41 NN4END[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_057_ N2MID[6] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_090_ NN4END[13] VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__clkbuf_1
X_073_ N4END[14] VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__clkbuf_1
XFILLER_2_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_20 FrameData[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_31 FrameStrobe[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_42 NN4END[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_056_ N2MID[7] VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_10_Left_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_7_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_039_ FrameStrobe[7] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__buf_1
XFILLER_1_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_10_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_072_ N4END[15] VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__clkbuf_1
XANTENNA_21 FrameData[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_32 FrameStrobe[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_10 FrameData[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_43 NN4END[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_320 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_055_ N1END[0] VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__buf_1
XFILLER_11_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_7_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_038_ FrameStrobe[6] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__buf_1
XFILLER_7_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_10_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_071_ N2END[0] VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__buf_1
XFILLER_2_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_11 FrameData[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_33 N4END[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_22 FrameData[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_7_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_054_ N1END[1] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__buf_1
XFILLER_11_173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_037_ FrameStrobe[5] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__buf_1
XFILLER_7_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_4_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_1_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_070_ N2END[1] VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__buf_1
XFILLER_4_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_12 FrameData[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_23 FrameData[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_34 NN4END[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_053_ N1END[2] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__buf_1
XFILLER_11_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_152 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_036_ FrameStrobe[4] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__buf_1
XFILLER_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_019_ FrameData[19] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__buf_1
XFILLER_0_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_2_Left_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_202 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_279 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_13 FrameData[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_24 FrameData[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_35 NN4END[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_052_ N1END[3] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_7_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_035_ FrameStrobe[3] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__clkbuf_1
X_104_ UserCLK VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__buf_2
XFILLER_7_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_018_ FrameData[18] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__buf_1
XFILLER_0_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_14 FrameData[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_25 FrameData[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_36 NN4END[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_051_ FrameStrobe[19] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_7_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_034_ FrameStrobe[2] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__buf_1
XFILLER_7_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_103_ NN4END[0] VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__clkbuf_1
XFILLER_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_017_ FrameData[17] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__buf_1
XFILLER_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_15 FrameData[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_26 FrameData[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_37 NN4END[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_050_ FrameStrobe[18] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__clkbuf_1
Xoutput100 net100 VGND VGND VPWR VPWR SS4BEG[5] sky130_fd_sc_hd__buf_2
XFILLER_11_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_033_ FrameStrobe[1] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__buf_1
XFILLER_3_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_102_ NN4END[1] VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__clkbuf_1
XFILLER_8_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_016_ FrameData[16] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__buf_1
XFILLER_8_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_232 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_246 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_16 FrameData[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_6_Left_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput101 net101 VGND VGND VPWR VPWR SS4BEG[6] sky130_fd_sc_hd__buf_2
XANTENNA_27 FrameData[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_38 NN4END[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_032_ FrameStrobe[0] VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__buf_1
X_101_ NN4END[2] VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__clkbuf_1
XFILLER_8_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_9_Left_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_015_ FrameData[15] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__buf_1
XFILLER_0_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_258 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_17 FrameData[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput102 net102 VGND VGND VPWR VPWR SS4BEG[7] sky130_fd_sc_hd__buf_2
XANTENNA_28 FrameData[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_39 NN4END[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_031_ FrameData[31] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__buf_1
XFILLER_9_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_100_ NN4END[3] VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__clkbuf_1
XFILLER_8_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_014_ FrameData[14] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__buf_1
XFILLER_8_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_18 FrameData[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput103 net103 VGND VGND VPWR VPWR SS4BEG[8] sky130_fd_sc_hd__buf_2
XANTENNA_29 net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_030_ FrameData[30] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__buf_1
XFILLER_0_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_013_ FrameData[13] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__buf_1
XFILLER_3_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput104 net104 VGND VGND VPWR VPWR SS4BEG[9] sky130_fd_sc_hd__buf_2
XANTENNA_19 FrameData[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_89 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_089_ NN4END[14] VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__clkbuf_1
XFILLER_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_012_ FrameData[12] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__buf_1
XFILLER_5_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput105 net105 VGND VGND VPWR VPWR UserCLKo sky130_fd_sc_hd__buf_1
XFILLER_11_68 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_088_ NN4END[15] VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_8_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_011_ FrameData[11] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__buf_1
XFILLER_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_26 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_1_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_1_Left_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_087_ N4END[0] VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_8_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_010_ FrameData[10] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_5_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_38 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_086_ N4END[1] VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__clkbuf_1
XFILLER_3_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_8_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_069_ N2END[2] VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__buf_1
XFILLER_9_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput90 net90 VGND VGND VPWR VPWR SS4BEG[10] sky130_fd_sc_hd__buf_2
XFILLER_2_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_085_ N4END[2] VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__clkbuf_1
XFILLER_3_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_068_ N2END[3] VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__buf_1
XFILLER_9_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_5_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_302 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput1 net1 VGND VGND VPWR VPWR FrameData_O[0] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_2_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput80 net80 VGND VGND VPWR VPWR S4BEG[1] sky130_fd_sc_hd__buf_2
Xoutput91 net91 VGND VGND VPWR VPWR SS4BEG[11] sky130_fd_sc_hd__buf_2
XFILLER_10_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_5_Left_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_084_ N4END[3] VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__clkbuf_1
XFILLER_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_067_ N2END[4] VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__buf_1
XFILLER_0_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_8_Left_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_314 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput81 net81 VGND VGND VPWR VPWR S4BEG[2] sky130_fd_sc_hd__buf_2
Xoutput70 net70 VGND VGND VPWR VPWR S2BEGb[5] sky130_fd_sc_hd__buf_2
Xoutput92 net92 VGND VGND VPWR VPWR SS4BEG[12] sky130_fd_sc_hd__buf_2
Xoutput2 net2 VGND VGND VPWR VPWR FrameData_O[10] sky130_fd_sc_hd__buf_2
XFILLER_10_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_9_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_083_ N4END[4] VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__buf_1
XFILLER_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_066_ N2END[5] VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__buf_1
XFILLER_0_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_049_ FrameStrobe[17] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__clkbuf_1
XFILLER_4_223 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_1 FrameData[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput3 net3 VGND VGND VPWR VPWR FrameData_O[11] sky130_fd_sc_hd__buf_2
Xoutput82 net82 VGND VGND VPWR VPWR S4BEG[3] sky130_fd_sc_hd__buf_2
Xoutput71 net71 VGND VGND VPWR VPWR S2BEGb[6] sky130_fd_sc_hd__buf_2
Xoutput60 net60 VGND VGND VPWR VPWR S2BEG[3] sky130_fd_sc_hd__buf_2
Xoutput93 net93 VGND VGND VPWR VPWR SS4BEG[13] sky130_fd_sc_hd__buf_2
XFILLER_6_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_082_ N4END[5] VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__buf_1
XFILLER_2_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_065_ N2END[6] VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__buf_1
X_048_ FrameStrobe[16] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__clkbuf_1
XFILLER_4_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_2 FrameData[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput50 net50 VGND VGND VPWR VPWR FrameStrobe_O[7] sky130_fd_sc_hd__buf_2
XFILLER_9_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput4 net4 VGND VGND VPWR VPWR FrameData_O[12] sky130_fd_sc_hd__buf_2
Xoutput83 net83 VGND VGND VPWR VPWR S4BEG[4] sky130_fd_sc_hd__buf_2
Xoutput72 net72 VGND VGND VPWR VPWR S2BEGb[7] sky130_fd_sc_hd__buf_2
Xoutput61 net61 VGND VGND VPWR VPWR S2BEG[4] sky130_fd_sc_hd__buf_2
Xoutput94 net94 VGND VGND VPWR VPWR SS4BEG[14] sky130_fd_sc_hd__buf_2
XFILLER_9_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_081_ N4END[6] VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__buf_1
XFILLER_2_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_064_ N2END[7] VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__buf_1
XFILLER_2_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_047_ FrameStrobe[15] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_3 FrameData[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput40 net40 VGND VGND VPWR VPWR FrameStrobe_O[16] sky130_fd_sc_hd__buf_2
Xoutput51 net51 VGND VGND VPWR VPWR FrameStrobe_O[8] sky130_fd_sc_hd__buf_2
Xoutput5 net5 VGND VGND VPWR VPWR FrameData_O[13] sky130_fd_sc_hd__buf_2
Xoutput84 net84 VGND VGND VPWR VPWR S4BEG[5] sky130_fd_sc_hd__buf_2
Xoutput73 net73 VGND VGND VPWR VPWR S4BEG[0] sky130_fd_sc_hd__buf_2
Xoutput62 net62 VGND VGND VPWR VPWR S2BEG[5] sky130_fd_sc_hd__buf_2
Xoutput95 net95 VGND VGND VPWR VPWR SS4BEG[15] sky130_fd_sc_hd__buf_2
XFILLER_6_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_080_ N4END[7] VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_8_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_063_ N2MID[0] VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__buf_1
XFILLER_2_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_046_ FrameStrobe[14] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_029_ FrameData[29] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__clkbuf_1
XANTENNA_4 FrameData[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput41 net41 VGND VGND VPWR VPWR FrameStrobe_O[17] sky130_fd_sc_hd__buf_2
Xoutput52 net52 VGND VGND VPWR VPWR FrameStrobe_O[9] sky130_fd_sc_hd__buf_2
Xoutput6 net6 VGND VGND VPWR VPWR FrameData_O[14] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_2_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput30 net30 VGND VGND VPWR VPWR FrameData_O[7] sky130_fd_sc_hd__buf_2
Xoutput63 net63 VGND VGND VPWR VPWR S2BEG[6] sky130_fd_sc_hd__buf_2
Xoutput85 net85 VGND VGND VPWR VPWR S4BEG[6] sky130_fd_sc_hd__buf_2
Xoutput74 net74 VGND VGND VPWR VPWR S4BEG[10] sky130_fd_sc_hd__buf_2
Xoutput96 net96 VGND VGND VPWR VPWR SS4BEG[1] sky130_fd_sc_hd__buf_2
.ends

