module W_IO (A_I_top,
    A_O_top,
    A_T_top,
    A_config_C_bit0,
    A_config_C_bit1,
    A_config_C_bit2,
    A_config_C_bit3,
    B_I_top,
    B_O_top,
    B_T_top,
    B_config_C_bit0,
    B_config_C_bit1,
    B_config_C_bit2,
    B_config_C_bit3,
    UserCLK,
    UserCLKo,
    VPWR,
    VGND,
    E1BEG,
    E2BEG,
    E2BEGb,
    E6BEG,
    EE4BEG,
    FrameData,
    FrameData_O,
    FrameStrobe,
    FrameStrobe_O,
    W1END,
    W2END,
    W2MID,
    W6END,
    WW4END);
 output A_I_top;
 input A_O_top;
 output A_T_top;
 output A_config_C_bit0;
 output A_config_C_bit1;
 output A_config_C_bit2;
 output A_config_C_bit3;
 output B_I_top;
 input B_O_top;
 output B_T_top;
 output B_config_C_bit0;
 output B_config_C_bit1;
 output B_config_C_bit2;
 output B_config_C_bit3;
 input UserCLK;
 output UserCLKo;
 inout VPWR;
 inout VGND;
 output [3:0] E1BEG;
 output [7:0] E2BEG;
 output [7:0] E2BEGb;
 output [11:0] E6BEG;
 output [15:0] EE4BEG;
 input [31:0] FrameData;
 output [31:0] FrameData_O;
 input [19:0] FrameStrobe;
 output [19:0] FrameStrobe_O;
 input [3:0] W1END;
 input [7:0] W2END;
 input [7:0] W2MID;
 input [11:0] W6END;
 input [15:0] WW4END;

 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire \Inst_A_IO_1_bidirectional_frame_config_pass.Q ;
 wire \Inst_B_IO_1_bidirectional_frame_config_pass.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit0.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit1.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit10.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit11.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit12.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit13.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit14.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit15.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit16.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit17.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit18.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit19.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit2.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit20.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit21.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit22.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit23.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit24.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit25.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit26.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit27.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit28.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit29.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit3.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit30.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit31.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit4.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit5.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit6.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit7.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit8.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame0_bit9.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit0.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit1.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit10.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit11.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit12.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit13.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit14.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit15.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit16.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit17.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit18.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit19.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit2.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit20.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit21.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit22.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit23.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit24.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit25.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit26.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit27.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit28.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit29.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit3.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit30.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit31.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit4.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit5.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit6.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit7.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit8.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame1_bit9.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit0.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit1.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit10.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit11.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit12.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit13.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit14.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit15.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit16.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit17.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit18.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit19.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit2.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit20.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit21.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit22.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit23.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit24.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit25.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit26.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit27.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit28.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit29.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit3.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit30.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit31.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit4.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit5.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit6.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit7.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit8.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame2_bit9.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame3_bit22.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame3_bit23.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame3_bit24.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame3_bit25.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame3_bit26.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame3_bit27.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame3_bit28.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame3_bit29.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame3_bit30.Q ;
 wire \Inst_W_IO_ConfigMem.Inst_frame3_bit31.Q ;
 wire \Inst_W_IO_switch_matrix.E1BEG0 ;
 wire \Inst_W_IO_switch_matrix.E1BEG1 ;
 wire \Inst_W_IO_switch_matrix.E1BEG2 ;
 wire \Inst_W_IO_switch_matrix.E1BEG3 ;
 wire \Inst_W_IO_switch_matrix.E2BEG0 ;
 wire \Inst_W_IO_switch_matrix.E2BEG1 ;
 wire \Inst_W_IO_switch_matrix.E2BEG2 ;
 wire \Inst_W_IO_switch_matrix.E2BEG3 ;
 wire \Inst_W_IO_switch_matrix.E2BEG4 ;
 wire \Inst_W_IO_switch_matrix.E2BEG5 ;
 wire \Inst_W_IO_switch_matrix.E2BEG6 ;
 wire \Inst_W_IO_switch_matrix.E2BEG7 ;
 wire \Inst_W_IO_switch_matrix.E2BEGb0 ;
 wire \Inst_W_IO_switch_matrix.E2BEGb1 ;
 wire \Inst_W_IO_switch_matrix.E2BEGb2 ;
 wire \Inst_W_IO_switch_matrix.E2BEGb3 ;
 wire \Inst_W_IO_switch_matrix.E2BEGb4 ;
 wire \Inst_W_IO_switch_matrix.E2BEGb5 ;
 wire \Inst_W_IO_switch_matrix.E2BEGb6 ;
 wire \Inst_W_IO_switch_matrix.E2BEGb7 ;
 wire \Inst_W_IO_switch_matrix.E6BEG0 ;
 wire \Inst_W_IO_switch_matrix.E6BEG1 ;
 wire \Inst_W_IO_switch_matrix.E6BEG10 ;
 wire \Inst_W_IO_switch_matrix.E6BEG11 ;
 wire \Inst_W_IO_switch_matrix.E6BEG2 ;
 wire \Inst_W_IO_switch_matrix.E6BEG3 ;
 wire \Inst_W_IO_switch_matrix.E6BEG4 ;
 wire \Inst_W_IO_switch_matrix.E6BEG5 ;
 wire \Inst_W_IO_switch_matrix.E6BEG6 ;
 wire \Inst_W_IO_switch_matrix.E6BEG7 ;
 wire \Inst_W_IO_switch_matrix.E6BEG8 ;
 wire \Inst_W_IO_switch_matrix.E6BEG9 ;
 wire \Inst_W_IO_switch_matrix.EE4BEG0 ;
 wire \Inst_W_IO_switch_matrix.EE4BEG1 ;
 wire \Inst_W_IO_switch_matrix.EE4BEG10 ;
 wire \Inst_W_IO_switch_matrix.EE4BEG11 ;
 wire \Inst_W_IO_switch_matrix.EE4BEG12 ;
 wire \Inst_W_IO_switch_matrix.EE4BEG13 ;
 wire \Inst_W_IO_switch_matrix.EE4BEG14 ;
 wire \Inst_W_IO_switch_matrix.EE4BEG15 ;
 wire \Inst_W_IO_switch_matrix.EE4BEG2 ;
 wire \Inst_W_IO_switch_matrix.EE4BEG3 ;
 wire \Inst_W_IO_switch_matrix.EE4BEG4 ;
 wire \Inst_W_IO_switch_matrix.EE4BEG5 ;
 wire \Inst_W_IO_switch_matrix.EE4BEG6 ;
 wire \Inst_W_IO_switch_matrix.EE4BEG7 ;
 wire \Inst_W_IO_switch_matrix.EE4BEG8 ;
 wire \Inst_W_IO_switch_matrix.EE4BEG9 ;
 wire net218;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire net220;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net219;

 sg13g2_inv_1 _049_ (.VDD(VPWR),
    .Y(_000_),
    .A(net40),
    .VSS(VGND));
 sg13g2_inv_1 _050_ (.VDD(VPWR),
    .Y(_001_),
    .A(\Inst_W_IO_ConfigMem.Inst_frame0_bit24.Q ),
    .VSS(VGND));
 sg13g2_mux2_1 _051_ (.A0(net41),
    .A1(net42),
    .S(\Inst_W_IO_ConfigMem.Inst_frame0_bit25.Q ),
    .X(_002_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _052_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_003_),
    .B(net39),
    .A(net66));
 sg13g2_a21oi_1 _053_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net66),
    .A2(_000_),
    .Y(_004_),
    .B1(\Inst_W_IO_ConfigMem.Inst_frame0_bit26.Q ));
 sg13g2_a221oi_1 _054_ (.VSS(VGND),
    .VDD(VPWR),
    .B2(_004_),
    .C1(\Inst_W_IO_ConfigMem.Inst_frame0_bit27.Q ),
    .B1(_003_),
    .A1(\Inst_W_IO_ConfigMem.Inst_frame0_bit26.Q ),
    .Y(_005_),
    .A2(_002_));
 sg13g2_nand2_1 _055_ (.Y(_006_),
    .A(net66),
    .B(net44),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _056_ (.Y(_007_),
    .B(net43),
    .A_N(net66),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _057_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_006_),
    .A2(_007_),
    .Y(_008_),
    .B1(\Inst_W_IO_ConfigMem.Inst_frame0_bit26.Q ));
 sg13g2_nor2b_1 _058_ (.A(net46),
    .B_N(net66),
    .Y(_009_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _059_ (.B1(\Inst_W_IO_ConfigMem.Inst_frame0_bit26.Q ),
    .VDD(VPWR),
    .Y(_010_),
    .VSS(VGND),
    .A1(net66),
    .A2(net45));
 sg13g2_o21ai_1 _060_ (.B1(\Inst_W_IO_ConfigMem.Inst_frame0_bit27.Q ),
    .VDD(VPWR),
    .Y(_011_),
    .VSS(VGND),
    .A1(_009_),
    .A2(_010_));
 sg13g2_o21ai_1 _061_ (.B1(\Inst_W_IO_ConfigMem.Inst_frame0_bit28.Q ),
    .VDD(VPWR),
    .Y(_012_),
    .VSS(VGND),
    .A1(_008_),
    .A2(_011_));
 sg13g2_mux4_1 _062_ (.S0(net66),
    .A0(net47),
    .A1(net48),
    .A2(net49),
    .A3(net50),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame0_bit26.Q ),
    .X(_013_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _063_ (.S0(net66),
    .A0(net51),
    .A1(net52),
    .A2(net53),
    .A3(net54),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame0_bit26.Q ),
    .X(_014_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _064_ (.A0(_013_),
    .A1(_014_),
    .S(\Inst_W_IO_ConfigMem.Inst_frame0_bit27.Q ),
    .X(_015_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _065_ (.Y(_016_),
    .B(_015_),
    .A_N(\Inst_W_IO_ConfigMem.Inst_frame0_bit28.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _066_ (.B1(_016_),
    .VDD(VPWR),
    .Y(net112),
    .VSS(VGND),
    .A1(_005_),
    .A2(_012_));
 sg13g2_mux2_1 _067_ (.A0(net41),
    .A1(net42),
    .S(net67),
    .X(_017_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _068_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_018_),
    .B(net67),
    .A(net39));
 sg13g2_a21oi_1 _069_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_000_),
    .A2(net67),
    .Y(_019_),
    .B1(\Inst_W_IO_ConfigMem.Inst_frame0_bit19.Q ));
 sg13g2_a221oi_1 _070_ (.VSS(VGND),
    .VDD(VPWR),
    .B2(_019_),
    .C1(\Inst_W_IO_ConfigMem.Inst_frame0_bit20.Q ),
    .B1(_018_),
    .A1(\Inst_W_IO_ConfigMem.Inst_frame0_bit19.Q ),
    .Y(_020_),
    .A2(_017_));
 sg13g2_nand2_1 _071_ (.Y(_021_),
    .A(net44),
    .B(net67),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _072_ (.Y(_022_),
    .B(net43),
    .A_N(net67),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _073_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_021_),
    .A2(_022_),
    .Y(_023_),
    .B1(\Inst_W_IO_ConfigMem.Inst_frame0_bit19.Q ));
 sg13g2_nor2b_1 _074_ (.A(net46),
    .B_N(net67),
    .Y(_024_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _075_ (.B1(\Inst_W_IO_ConfigMem.Inst_frame0_bit19.Q ),
    .VDD(VPWR),
    .Y(_025_),
    .VSS(VGND),
    .A1(net45),
    .A2(net67));
 sg13g2_o21ai_1 _076_ (.B1(\Inst_W_IO_ConfigMem.Inst_frame0_bit20.Q ),
    .VDD(VPWR),
    .Y(_026_),
    .VSS(VGND),
    .A1(_024_),
    .A2(_025_));
 sg13g2_o21ai_1 _077_ (.B1(\Inst_W_IO_ConfigMem.Inst_frame0_bit21.Q ),
    .VDD(VPWR),
    .Y(_027_),
    .VSS(VGND),
    .A1(_023_),
    .A2(_026_));
 sg13g2_mux4_1 _078_ (.S0(\Inst_W_IO_ConfigMem.Inst_frame0_bit18.Q ),
    .A0(net47),
    .A1(net48),
    .A2(net49),
    .A3(net50),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame0_bit19.Q ),
    .X(_028_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _079_ (.S0(net67),
    .A0(net51),
    .A1(net52),
    .A2(net53),
    .A3(net54),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame0_bit19.Q ),
    .X(_029_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _080_ (.A0(_028_),
    .A1(_029_),
    .S(\Inst_W_IO_ConfigMem.Inst_frame0_bit20.Q ),
    .X(_030_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _081_ (.Y(_031_),
    .B(_030_),
    .A_N(\Inst_W_IO_ConfigMem.Inst_frame0_bit21.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _082_ (.B1(_031_),
    .VDD(VPWR),
    .Y(net106),
    .VSS(VGND),
    .A1(_020_),
    .A2(_027_));
 sg13g2_mux4_1 _083_ (.S0(\Inst_W_IO_ConfigMem.Inst_frame0_bit16.Q ),
    .A0(net35),
    .A1(net90),
    .A2(net55),
    .A3(\Inst_B_IO_1_bidirectional_frame_config_pass.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame0_bit17.Q ),
    .X(\Inst_W_IO_switch_matrix.E6BEG11 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _084_ (.S0(\Inst_W_IO_ConfigMem.Inst_frame0_bit14.Q ),
    .A0(net36),
    .A1(net97),
    .A2(net58),
    .A3(\Inst_A_IO_1_bidirectional_frame_config_pass.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame0_bit15.Q ),
    .X(\Inst_W_IO_switch_matrix.E6BEG10 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _085_ (.S0(\Inst_W_IO_ConfigMem.Inst_frame0_bit12.Q ),
    .A0(net100),
    .A1(net93),
    .A2(net61),
    .A3(\Inst_B_IO_1_bidirectional_frame_config_pass.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame0_bit13.Q ),
    .X(\Inst_W_IO_switch_matrix.E6BEG9 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _086_ (.S0(\Inst_W_IO_ConfigMem.Inst_frame0_bit10.Q ),
    .A0(net101),
    .A1(net94),
    .A2(net62),
    .A3(\Inst_A_IO_1_bidirectional_frame_config_pass.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame0_bit11.Q ),
    .X(\Inst_W_IO_switch_matrix.E6BEG8 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _087_ (.S0(\Inst_W_IO_ConfigMem.Inst_frame0_bit8.Q ),
    .A0(net35),
    .A1(net104),
    .A2(net65),
    .A3(\Inst_B_IO_1_bidirectional_frame_config_pass.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame0_bit9.Q ),
    .X(\Inst_W_IO_switch_matrix.E6BEG7 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _088_ (.S0(\Inst_W_IO_ConfigMem.Inst_frame0_bit6.Q ),
    .A0(net36),
    .A1(net105),
    .A2(net89),
    .A3(\Inst_A_IO_1_bidirectional_frame_config_pass.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame0_bit7.Q ),
    .X(\Inst_W_IO_switch_matrix.E6BEG6 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _089_ (.S0(\Inst_W_IO_ConfigMem.Inst_frame0_bit4.Q ),
    .A0(net38),
    .A1(net98),
    .A2(net59),
    .A3(net2),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame0_bit5.Q ),
    .X(\Inst_W_IO_switch_matrix.E6BEG5 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _090_ (.S0(\Inst_W_IO_ConfigMem.Inst_frame0_bit2.Q ),
    .A0(net37),
    .A1(net99),
    .A2(net60),
    .A3(net1),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame0_bit3.Q ),
    .X(\Inst_W_IO_switch_matrix.E6BEG4 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _091_ (.S0(\Inst_W_IO_ConfigMem.Inst_frame0_bit0.Q ),
    .A0(net102),
    .A1(net95),
    .A2(net63),
    .A3(net2),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame0_bit1.Q ),
    .X(\Inst_W_IO_switch_matrix.E6BEG3 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _092_ (.S0(\Inst_W_IO_ConfigMem.Inst_frame1_bit30.Q ),
    .A0(net103),
    .A1(net96),
    .A2(net64),
    .A3(net1),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame1_bit31.Q ),
    .X(\Inst_W_IO_switch_matrix.E6BEG2 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _093_ (.S0(\Inst_W_IO_ConfigMem.Inst_frame1_bit28.Q ),
    .A0(net38),
    .A1(net91),
    .A2(net56),
    .A3(net2),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame1_bit29.Q ),
    .X(\Inst_W_IO_switch_matrix.E6BEG1 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _094_ (.S0(\Inst_W_IO_ConfigMem.Inst_frame1_bit26.Q ),
    .A0(net37),
    .A1(net92),
    .A2(net57),
    .A3(net1),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame1_bit27.Q ),
    .X(\Inst_W_IO_switch_matrix.E6BEG0 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _095_ (.S0(\Inst_W_IO_ConfigMem.Inst_frame1_bit25.Q ),
    .A0(net48),
    .A1(net52),
    .A2(net50),
    .A3(net54),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame1_bit24.Q ),
    .X(\Inst_W_IO_switch_matrix.EE4BEG15 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _096_ (.S0(\Inst_W_IO_ConfigMem.Inst_frame1_bit23.Q ),
    .A0(net47),
    .A1(net51),
    .A2(net49),
    .A3(net53),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame1_bit22.Q ),
    .X(\Inst_W_IO_switch_matrix.EE4BEG14 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _097_ (.S0(\Inst_W_IO_ConfigMem.Inst_frame1_bit21.Q ),
    .A0(net64),
    .A1(net57),
    .A2(net89),
    .A3(\Inst_B_IO_1_bidirectional_frame_config_pass.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame1_bit20.Q ),
    .X(\Inst_W_IO_switch_matrix.EE4BEG13 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _098_ (.S0(\Inst_W_IO_ConfigMem.Inst_frame1_bit19.Q ),
    .A0(net58),
    .A1(net62),
    .A2(net60),
    .A3(\Inst_A_IO_1_bidirectional_frame_config_pass.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame1_bit18.Q ),
    .X(\Inst_W_IO_switch_matrix.EE4BEG12 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _099_ (.S0(\Inst_W_IO_ConfigMem.Inst_frame1_bit17.Q ),
    .A0(net63),
    .A1(net56),
    .A2(net65),
    .A3(net2),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame1_bit16.Q ),
    .X(\Inst_W_IO_switch_matrix.EE4BEG11 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _100_ (.S0(\Inst_W_IO_ConfigMem.Inst_frame1_bit15.Q ),
    .A0(net55),
    .A1(net61),
    .A2(net59),
    .A3(net1),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame1_bit14.Q ),
    .X(\Inst_W_IO_switch_matrix.EE4BEG10 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _101_ (.S0(\Inst_W_IO_ConfigMem.Inst_frame1_bit13.Q ),
    .A0(net58),
    .A1(net62),
    .A2(net60),
    .A3(net64),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame1_bit12.Q ),
    .X(\Inst_W_IO_switch_matrix.EE4BEG9 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _102_ (.S0(\Inst_W_IO_ConfigMem.Inst_frame1_bit11.Q ),
    .A0(net61),
    .A1(net65),
    .A2(net63),
    .A3(net56),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame1_bit10.Q ),
    .X(\Inst_W_IO_switch_matrix.EE4BEG8 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _103_ (.S0(\Inst_W_IO_ConfigMem.Inst_frame1_bit9.Q ),
    .A0(net48),
    .A1(net52),
    .A2(net50),
    .A3(net54),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame1_bit8.Q ),
    .X(\Inst_W_IO_switch_matrix.EE4BEG7 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _104_ (.S0(\Inst_W_IO_ConfigMem.Inst_frame1_bit7.Q ),
    .A0(net47),
    .A1(net51),
    .A2(net49),
    .A3(net53),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame1_bit6.Q ),
    .X(\Inst_W_IO_switch_matrix.EE4BEG6 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _105_ (.S0(\Inst_W_IO_ConfigMem.Inst_frame1_bit4.Q ),
    .A0(net40),
    .A1(net42),
    .A2(net44),
    .A3(net46),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame1_bit5.Q ),
    .X(\Inst_W_IO_switch_matrix.EE4BEG5 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _106_ (.S0(\Inst_W_IO_ConfigMem.Inst_frame1_bit2.Q ),
    .A0(net39),
    .A1(net41),
    .A2(net43),
    .A3(net45),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame1_bit3.Q ),
    .X(\Inst_W_IO_switch_matrix.EE4BEG4 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _107_ (.S0(\Inst_W_IO_ConfigMem.Inst_frame1_bit1.Q ),
    .A0(net64),
    .A1(net57),
    .A2(net89),
    .A3(\Inst_B_IO_1_bidirectional_frame_config_pass.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame1_bit0.Q ),
    .X(\Inst_W_IO_switch_matrix.EE4BEG3 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _108_ (.S0(\Inst_W_IO_ConfigMem.Inst_frame2_bit31.Q ),
    .A0(net58),
    .A1(net62),
    .A2(net60),
    .A3(\Inst_A_IO_1_bidirectional_frame_config_pass.Q ),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame2_bit30.Q ),
    .X(\Inst_W_IO_switch_matrix.EE4BEG2 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _109_ (.S0(\Inst_W_IO_ConfigMem.Inst_frame2_bit29.Q ),
    .A0(net63),
    .A1(net56),
    .A2(net65),
    .A3(net2),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame2_bit28.Q ),
    .X(\Inst_W_IO_switch_matrix.EE4BEG1 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _110_ (.S0(\Inst_W_IO_ConfigMem.Inst_frame2_bit27.Q ),
    .A0(net55),
    .A1(net61),
    .A2(net59),
    .A3(net1),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame2_bit26.Q ),
    .X(\Inst_W_IO_switch_matrix.EE4BEG0 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _111_ (.S0(\Inst_W_IO_ConfigMem.Inst_frame2_bit24.Q ),
    .A0(net39),
    .A1(net90),
    .A2(net104),
    .A3(net55),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame2_bit25.Q ),
    .X(\Inst_W_IO_switch_matrix.E2BEGb7 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _112_ (.S0(\Inst_W_IO_ConfigMem.Inst_frame2_bit22.Q ),
    .A0(net40),
    .A1(net97),
    .A2(net105),
    .A3(net58),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame2_bit23.Q ),
    .X(\Inst_W_IO_switch_matrix.E2BEGb6 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _113_ (.S0(\Inst_W_IO_ConfigMem.Inst_frame2_bit20.Q ),
    .A0(net41),
    .A1(net98),
    .A2(net91),
    .A3(net59),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame2_bit21.Q ),
    .X(\Inst_W_IO_switch_matrix.E2BEGb5 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _114_ (.S0(\Inst_W_IO_ConfigMem.Inst_frame2_bit18.Q ),
    .A0(net42),
    .A1(net99),
    .A2(net92),
    .A3(net60),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame2_bit19.Q ),
    .X(\Inst_W_IO_switch_matrix.E2BEGb4 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _115_ (.S0(\Inst_W_IO_ConfigMem.Inst_frame2_bit16.Q ),
    .A0(net43),
    .A1(net100),
    .A2(net93),
    .A3(net61),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame2_bit17.Q ),
    .X(\Inst_W_IO_switch_matrix.E2BEGb3 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _116_ (.S0(\Inst_W_IO_ConfigMem.Inst_frame2_bit14.Q ),
    .A0(net44),
    .A1(net101),
    .A2(net94),
    .A3(net62),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame2_bit15.Q ),
    .X(\Inst_W_IO_switch_matrix.E2BEGb2 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _117_ (.S0(\Inst_W_IO_ConfigMem.Inst_frame2_bit12.Q ),
    .A0(net45),
    .A1(net102),
    .A2(net95),
    .A3(net63),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame2_bit13.Q ),
    .X(\Inst_W_IO_switch_matrix.E2BEGb1 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _118_ (.S0(\Inst_W_IO_ConfigMem.Inst_frame2_bit10.Q ),
    .A0(net46),
    .A1(net103),
    .A2(net96),
    .A3(net64),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame2_bit11.Q ),
    .X(\Inst_W_IO_switch_matrix.E2BEGb0 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _119_ (.S0(\Inst_W_IO_ConfigMem.Inst_frame2_bit8.Q ),
    .A0(net47),
    .A1(net90),
    .A2(net104),
    .A3(net55),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame2_bit9.Q ),
    .X(\Inst_W_IO_switch_matrix.E2BEG7 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _120_ (.S0(\Inst_W_IO_ConfigMem.Inst_frame2_bit6.Q ),
    .A0(net48),
    .A1(net97),
    .A2(net105),
    .A3(net58),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame2_bit7.Q ),
    .X(\Inst_W_IO_switch_matrix.E2BEG6 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _121_ (.S0(\Inst_W_IO_ConfigMem.Inst_frame2_bit4.Q ),
    .A0(net49),
    .A1(net98),
    .A2(net91),
    .A3(net59),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame2_bit5.Q ),
    .X(\Inst_W_IO_switch_matrix.E2BEG5 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _122_ (.S0(\Inst_W_IO_ConfigMem.Inst_frame2_bit2.Q ),
    .A0(net50),
    .A1(net99),
    .A2(net92),
    .A3(net60),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame2_bit3.Q ),
    .X(\Inst_W_IO_switch_matrix.E2BEG4 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _123_ (.S0(\Inst_W_IO_ConfigMem.Inst_frame2_bit0.Q ),
    .A0(net51),
    .A1(net100),
    .A2(net93),
    .A3(net61),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame2_bit1.Q ),
    .X(\Inst_W_IO_switch_matrix.E2BEG3 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _124_ (.S0(\Inst_W_IO_ConfigMem.Inst_frame3_bit30.Q ),
    .A0(net52),
    .A1(net101),
    .A2(net94),
    .A3(net62),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame3_bit31.Q ),
    .X(\Inst_W_IO_switch_matrix.E2BEG2 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _125_ (.S0(\Inst_W_IO_ConfigMem.Inst_frame3_bit28.Q ),
    .A0(net53),
    .A1(net102),
    .A2(net95),
    .A3(net63),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame3_bit29.Q ),
    .X(\Inst_W_IO_switch_matrix.E2BEG1 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _126_ (.S0(\Inst_W_IO_ConfigMem.Inst_frame3_bit26.Q ),
    .A0(net54),
    .A1(net103),
    .A2(net96),
    .A3(net64),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame3_bit27.Q ),
    .X(\Inst_W_IO_switch_matrix.E2BEG0 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _127_ (.A0(net35),
    .A1(\Inst_B_IO_1_bidirectional_frame_config_pass.Q ),
    .S(\Inst_W_IO_ConfigMem.Inst_frame3_bit25.Q ),
    .X(\Inst_W_IO_switch_matrix.E1BEG3 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _128_ (.A0(net36),
    .A1(net2),
    .S(\Inst_W_IO_ConfigMem.Inst_frame3_bit24.Q ),
    .X(\Inst_W_IO_switch_matrix.E1BEG2 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _129_ (.A0(net37),
    .A1(\Inst_A_IO_1_bidirectional_frame_config_pass.Q ),
    .S(\Inst_W_IO_ConfigMem.Inst_frame3_bit23.Q ),
    .X(\Inst_W_IO_switch_matrix.E1BEG1 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _130_ (.A0(net38),
    .A1(net1),
    .S(\Inst_W_IO_ConfigMem.Inst_frame3_bit22.Q ),
    .X(\Inst_W_IO_switch_matrix.E1BEG0 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _131_ (.Y(_032_),
    .B(\Inst_W_IO_ConfigMem.Inst_frame0_bit24.Q ),
    .A_N(net42),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _132_ (.B1(_032_),
    .VDD(VPWR),
    .Y(_033_),
    .VSS(VGND),
    .A1(net54),
    .A2(\Inst_W_IO_ConfigMem.Inst_frame0_bit24.Q ));
 sg13g2_nand3_1 _133_ (.B(\Inst_W_IO_ConfigMem.Inst_frame0_bit23.Q ),
    .C(_001_),
    .A(net40),
    .Y(_034_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _134_ (.B1(_034_),
    .VDD(VPWR),
    .Y(_035_),
    .VSS(VGND),
    .A1(\Inst_W_IO_ConfigMem.Inst_frame0_bit23.Q ),
    .A2(_033_));
 sg13g2_nand3b_1 _135_ (.B(_001_),
    .C(net39),
    .Y(_036_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(\Inst_W_IO_ConfigMem.Inst_frame0_bit23.Q ));
 sg13g2_o21ai_1 _136_ (.B1(\Inst_W_IO_ConfigMem.Inst_frame0_bit23.Q ),
    .VDD(VPWR),
    .Y(_037_),
    .VSS(VGND),
    .A1(net41),
    .A2(\Inst_W_IO_ConfigMem.Inst_frame0_bit24.Q ));
 sg13g2_nand2_1 _137_ (.Y(_038_),
    .A(net43),
    .B(\Inst_W_IO_ConfigMem.Inst_frame0_bit24.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _138_ (.B(_036_),
    .C(_037_),
    .A(\Inst_W_IO_ConfigMem.Inst_frame0_bit22.Q ),
    .Y(_039_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_038_));
 sg13g2_o21ai_1 _139_ (.B1(_039_),
    .VDD(VPWR),
    .Y(net107),
    .VSS(VGND),
    .A1(\Inst_W_IO_ConfigMem.Inst_frame0_bit22.Q ),
    .A2(_035_));
 sg13g2_nand2b_1 _140_ (.Y(_040_),
    .B(net44),
    .A_N(\Inst_W_IO_ConfigMem.Inst_frame0_bit30.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _141_ (.S0(\Inst_W_IO_ConfigMem.Inst_frame0_bit29.Q ),
    .A0(net53),
    .A1(net54),
    .A2(net39),
    .A3(net43),
    .S1(\Inst_W_IO_ConfigMem.Inst_frame0_bit30.Q ),
    .X(_041_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _142_ (.B1(\Inst_W_IO_ConfigMem.Inst_frame0_bit29.Q ),
    .VDD(VPWR),
    .Y(_042_),
    .VSS(VGND),
    .A1(net45),
    .A2(\Inst_W_IO_ConfigMem.Inst_frame0_bit30.Q ));
 sg13g2_o21ai_1 _143_ (.B1(\Inst_W_IO_ConfigMem.Inst_frame0_bit31.Q ),
    .VDD(VPWR),
    .Y(_043_),
    .VSS(VGND),
    .A1(\Inst_W_IO_ConfigMem.Inst_frame0_bit29.Q ),
    .A2(_040_));
 sg13g2_nand2b_1 _144_ (.Y(_044_),
    .B(_042_),
    .A_N(_043_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _145_ (.B1(_044_),
    .VDD(VPWR),
    .Y(net113),
    .VSS(VGND),
    .A1(\Inst_W_IO_ConfigMem.Inst_frame0_bit31.Q ),
    .A2(_041_));
 sg13g2_dlhq_1 _146_ (.D(net8),
    .GATE(net68),
    .Q(net108),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _147_ (.D(net9),
    .GATE(net68),
    .Q(net109),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _148_ (.D(net10),
    .GATE(net68),
    .Q(net110),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _149_ (.D(net11),
    .GATE(net68),
    .Q(net111),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _150_ (.D(net12),
    .GATE(net68),
    .Q(net114),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _151_ (.D(net13),
    .GATE(net68),
    .Q(net115),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _152_ (.D(net15),
    .GATE(net68),
    .Q(net116),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _153_ (.D(net16),
    .GATE(net68),
    .Q(net117),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _154_ (.D(net17),
    .GATE(net69),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame3_bit22.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _155_ (.D(net18),
    .GATE(net71),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame3_bit23.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _156_ (.D(net19),
    .GATE(net69),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame3_bit24.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _157_ (.D(net20),
    .GATE(net71),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame3_bit25.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _158_ (.D(net21),
    .GATE(net69),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame3_bit26.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _159_ (.D(net22),
    .GATE(net69),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame3_bit27.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _160_ (.D(net23),
    .GATE(net70),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame3_bit28.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _161_ (.D(net24),
    .GATE(net70),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame3_bit29.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _162_ (.D(net26),
    .GATE(net70),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame3_bit30.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _163_ (.D(net27),
    .GATE(net70),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame3_bit31.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _164_ (.D(net3),
    .GATE(net75),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit0.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _165_ (.D(net14),
    .GATE(net74),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit1.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _166_ (.D(net25),
    .GATE(net75),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit2.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _167_ (.D(net28),
    .GATE(net74),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit3.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _168_ (.D(net29),
    .GATE(net73),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit4.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _169_ (.D(net30),
    .GATE(net73),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit5.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _170_ (.D(net31),
    .GATE(net73),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit6.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _171_ (.D(net32),
    .GATE(net73),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit7.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _172_ (.D(net33),
    .GATE(net74),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit8.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _173_ (.D(net34),
    .GATE(net74),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit9.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _174_ (.D(net4),
    .GATE(net76),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit10.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _175_ (.D(net5),
    .GATE(net76),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit11.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _176_ (.D(net6),
    .GATE(net76),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit12.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _177_ (.D(net7),
    .GATE(net76),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit13.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _178_ (.D(net8),
    .GATE(net74),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit14.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _179_ (.D(net9),
    .GATE(net74),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit15.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _180_ (.D(net10),
    .GATE(net74),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit16.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _181_ (.D(net11),
    .GATE(net74),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit17.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _182_ (.D(net12),
    .GATE(net72),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit18.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _183_ (.D(net13),
    .GATE(net72),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit19.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _184_ (.D(net15),
    .GATE(net72),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit20.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _185_ (.D(net16),
    .GATE(net72),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit21.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _186_ (.D(net17),
    .GATE(net72),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit22.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _187_ (.D(net18),
    .GATE(net72),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit23.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _188_ (.D(net19),
    .GATE(net72),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit24.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _189_ (.D(net20),
    .GATE(net72),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit25.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _190_ (.D(net21),
    .GATE(net76),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit26.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _191_ (.D(net22),
    .GATE(net76),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit27.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _192_ (.D(net23),
    .GATE(net76),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit28.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _193_ (.D(net24),
    .GATE(net76),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit29.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _194_ (.D(net26),
    .GATE(net77),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit30.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _195_ (.D(net27),
    .GATE(net77),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame2_bit31.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _196_ (.D(net3),
    .GATE(net80),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit0.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _197_ (.D(net14),
    .GATE(net82),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit1.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _198_ (.D(net25),
    .GATE(net82),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit2.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _199_ (.D(net28),
    .GATE(net78),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit3.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _200_ (.D(net29),
    .GATE(net79),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit4.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _201_ (.D(net30),
    .GATE(net79),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit5.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _202_ (.D(net31),
    .GATE(net78),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit6.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _203_ (.D(net32),
    .GATE(net78),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit7.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _204_ (.D(net33),
    .GATE(net78),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit8.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _205_ (.D(net34),
    .GATE(net78),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit9.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _206_ (.D(net4),
    .GATE(net81),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit10.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _207_ (.D(net5),
    .GATE(net81),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit11.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _208_ (.D(net6),
    .GATE(net80),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit12.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _209_ (.D(net7),
    .GATE(net80),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit13.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _210_ (.D(net8),
    .GATE(net81),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit14.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _211_ (.D(net9),
    .GATE(net81),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit15.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _212_ (.D(net10),
    .GATE(net81),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit16.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _213_ (.D(net11),
    .GATE(net81),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit17.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _214_ (.D(net12),
    .GATE(net80),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit18.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _215_ (.D(net13),
    .GATE(net80),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit19.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _216_ (.D(net15),
    .GATE(net80),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit20.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _217_ (.D(net16),
    .GATE(net80),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit21.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _218_ (.D(net17),
    .GATE(net79),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit22.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _219_ (.D(net18),
    .GATE(net79),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit23.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _220_ (.D(net19),
    .GATE(net79),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit24.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _221_ (.D(net20),
    .GATE(net79),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit25.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _222_ (.D(net21),
    .GATE(net81),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit26.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _223_ (.D(net22),
    .GATE(net81),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit27.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _224_ (.D(net23),
    .GATE(net78),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit28.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _225_ (.D(net24),
    .GATE(net79),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit29.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _226_ (.D(net26),
    .GATE(net78),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit30.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _227_ (.D(net27),
    .GATE(net78),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame1_bit31.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _228_ (.D(net3),
    .GATE(net85),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit0.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _229_ (.D(net14),
    .GATE(net85),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit1.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _230_ (.D(net25),
    .GATE(net85),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit2.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _231_ (.D(net28),
    .GATE(net85),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit3.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _232_ (.D(net29),
    .GATE(net88),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit4.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _233_ (.D(net30),
    .GATE(net88),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit5.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _234_ (.D(net31),
    .GATE(net87),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit6.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _235_ (.D(net32),
    .GATE(net87),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit7.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _236_ (.D(net33),
    .GATE(net86),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit8.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _237_ (.D(net34),
    .GATE(net86),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit9.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _238_ (.D(net4),
    .GATE(net85),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit10.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _239_ (.D(net5),
    .GATE(net85),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit11.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _240_ (.D(net6),
    .GATE(net85),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit12.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _241_ (.D(net7),
    .GATE(net85),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit13.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _242_ (.D(net8),
    .GATE(net87),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit14.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _243_ (.D(net9),
    .GATE(net87),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit15.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _244_ (.D(net10),
    .GATE(net86),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit16.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _245_ (.D(net11),
    .GATE(net86),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit17.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _246_ (.D(net12),
    .GATE(net83),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit18.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _247_ (.D(net13),
    .GATE(net84),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit19.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _248_ (.D(net15),
    .GATE(net84),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit20.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _249_ (.D(net16),
    .GATE(net83),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit21.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _250_ (.D(net17),
    .GATE(net83),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit22.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _251_ (.D(net18),
    .GATE(net83),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit23.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _252_ (.D(net19),
    .GATE(net83),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit24.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _253_ (.D(net20),
    .GATE(net83),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit25.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _254_ (.D(net21),
    .GATE(net84),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit26.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _255_ (.D(net22),
    .GATE(net83),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit27.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _256_ (.D(net23),
    .GATE(net83),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit28.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _257_ (.D(net24),
    .GATE(net84),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit29.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _258_ (.D(net26),
    .GATE(net84),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit30.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _259_ (.D(net27),
    .GATE(net84),
    .Q(\Inst_W_IO_ConfigMem.Inst_frame0_bit31.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dfrbp_1 _260_ (.CLK(UserCLK),
    .RESET_B(net219),
    .D(net1),
    .Q_N(_046_),
    .Q(\Inst_A_IO_1_bidirectional_frame_config_pass.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dfrbp_1 _261_ (.CLK(UserCLK),
    .RESET_B(net220),
    .D(net2),
    .Q_N(_045_),
    .Q(\Inst_B_IO_1_bidirectional_frame_config_pass.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_tiehi _261__197 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net220));
 sg13g2_decap_8 FILLER_0_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _264_ (.A(\Inst_W_IO_switch_matrix.E2BEG2 ),
    .X(net124),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _265_ (.A(\Inst_W_IO_switch_matrix.E2BEG3 ),
    .X(net125),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _266_ (.A(\Inst_W_IO_switch_matrix.E2BEG4 ),
    .X(net126),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _267_ (.A(\Inst_W_IO_switch_matrix.E2BEG5 ),
    .X(net127),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _268_ (.A(\Inst_W_IO_switch_matrix.E2BEG6 ),
    .X(net128),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _269_ (.A(\Inst_W_IO_switch_matrix.E2BEG7 ),
    .X(net129),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _270_ (.A(\Inst_W_IO_switch_matrix.E2BEGb0 ),
    .X(net130),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _271_ (.A(\Inst_W_IO_switch_matrix.E2BEGb1 ),
    .X(net131),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _272_ (.A(\Inst_W_IO_switch_matrix.E2BEGb2 ),
    .X(net132),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _273_ (.A(\Inst_W_IO_switch_matrix.E2BEGb3 ),
    .X(net133),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _274_ (.A(\Inst_W_IO_switch_matrix.E2BEGb4 ),
    .X(net134),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _275_ (.A(\Inst_W_IO_switch_matrix.E2BEGb5 ),
    .X(net135),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _276_ (.A(\Inst_W_IO_switch_matrix.E2BEGb6 ),
    .X(net136),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _277_ (.A(\Inst_W_IO_switch_matrix.E2BEGb7 ),
    .X(net137),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _278_ (.A(\Inst_W_IO_switch_matrix.E6BEG0 ),
    .X(net138),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _279_ (.A(\Inst_W_IO_switch_matrix.E6BEG1 ),
    .X(net141),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _280_ (.A(\Inst_W_IO_switch_matrix.E6BEG2 ),
    .X(net142),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _281_ (.A(\Inst_W_IO_switch_matrix.E6BEG3 ),
    .X(net143),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _282_ (.A(\Inst_W_IO_switch_matrix.E6BEG4 ),
    .X(net144),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _283_ (.A(\Inst_W_IO_switch_matrix.E6BEG5 ),
    .X(net145),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _284_ (.A(\Inst_W_IO_switch_matrix.E6BEG6 ),
    .X(net146),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _285_ (.A(\Inst_W_IO_switch_matrix.E6BEG7 ),
    .X(net147),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _286_ (.A(\Inst_W_IO_switch_matrix.E6BEG8 ),
    .X(net148),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _287_ (.A(\Inst_W_IO_switch_matrix.E6BEG9 ),
    .X(net149),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _288_ (.A(\Inst_W_IO_switch_matrix.E6BEG10 ),
    .X(net139),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _289_ (.A(\Inst_W_IO_switch_matrix.E6BEG11 ),
    .X(net140),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _290_ (.A(\Inst_W_IO_switch_matrix.EE4BEG0 ),
    .X(net150),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _291_ (.A(\Inst_W_IO_switch_matrix.EE4BEG1 ),
    .X(net157),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _292_ (.A(\Inst_W_IO_switch_matrix.EE4BEG2 ),
    .X(net158),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _293_ (.A(\Inst_W_IO_switch_matrix.EE4BEG3 ),
    .X(net159),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _294_ (.A(\Inst_W_IO_switch_matrix.EE4BEG4 ),
    .X(net160),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _295_ (.A(\Inst_W_IO_switch_matrix.EE4BEG5 ),
    .X(net161),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _296_ (.A(\Inst_W_IO_switch_matrix.EE4BEG6 ),
    .X(net162),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _297_ (.A(\Inst_W_IO_switch_matrix.EE4BEG7 ),
    .X(net163),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _298_ (.A(\Inst_W_IO_switch_matrix.EE4BEG8 ),
    .X(net164),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _299_ (.A(\Inst_W_IO_switch_matrix.EE4BEG9 ),
    .X(net165),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _300_ (.A(\Inst_W_IO_switch_matrix.EE4BEG10 ),
    .X(net151),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _301_ (.A(\Inst_W_IO_switch_matrix.EE4BEG11 ),
    .X(net152),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _302_ (.A(\Inst_W_IO_switch_matrix.EE4BEG12 ),
    .X(net153),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _303_ (.A(\Inst_W_IO_switch_matrix.EE4BEG13 ),
    .X(net154),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _304_ (.A(\Inst_W_IO_switch_matrix.EE4BEG14 ),
    .X(net155),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _305_ (.A(\Inst_W_IO_switch_matrix.EE4BEG15 ),
    .X(net156),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _306_ (.A(net3),
    .X(net166),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _307_ (.A(net14),
    .X(net177),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _308_ (.A(net25),
    .X(net188),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _309_ (.A(net28),
    .X(net191),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _310_ (.A(net29),
    .X(net192),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _311_ (.A(net30),
    .X(net193),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _312_ (.A(net31),
    .X(net194),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _313_ (.A(net32),
    .X(net195),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _314_ (.A(net33),
    .X(net196),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _315_ (.A(net34),
    .X(net197),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _316_ (.A(net4),
    .X(net167),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _317_ (.A(net5),
    .X(net168),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _318_ (.A(net6),
    .X(net169),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _319_ (.A(net7),
    .X(net170),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _320_ (.A(net8),
    .X(net171),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _321_ (.A(net9),
    .X(net172),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _322_ (.A(net10),
    .X(net173),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _323_ (.A(net11),
    .X(net174),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _324_ (.A(net12),
    .X(net175),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _325_ (.A(net13),
    .X(net176),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _326_ (.A(net15),
    .X(net178),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _327_ (.A(net16),
    .X(net179),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _328_ (.A(net17),
    .X(net180),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _329_ (.A(net18),
    .X(net181),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _330_ (.A(net19),
    .X(net182),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _331_ (.A(net20),
    .X(net183),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _332_ (.A(net21),
    .X(net184),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _333_ (.A(net22),
    .X(net185),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _334_ (.A(net23),
    .X(net186),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _335_ (.A(net24),
    .X(net187),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _336_ (.A(net26),
    .X(net189),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _337_ (.A(net27),
    .X(net190),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _338_ (.A(net87),
    .X(net198),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _339_ (.A(net80),
    .X(net209),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _340_ (.A(net77),
    .X(net210),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _341_ (.A(net71),
    .X(net211),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _342_ (.A(FrameStrobe[4]),
    .X(net212),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _343_ (.A(FrameStrobe[5]),
    .X(net213),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _344_ (.A(FrameStrobe[6]),
    .X(net214),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _345_ (.A(FrameStrobe[7]),
    .X(net215),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _346_ (.A(FrameStrobe[8]),
    .X(net216),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _347_ (.A(FrameStrobe[9]),
    .X(net217),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _348_ (.A(FrameStrobe[10]),
    .X(net199),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _349_ (.A(FrameStrobe[11]),
    .X(net200),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _350_ (.A(FrameStrobe[12]),
    .X(net201),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _351_ (.A(FrameStrobe[13]),
    .X(net202),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _352_ (.A(FrameStrobe[14]),
    .X(net203),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _353_ (.A(FrameStrobe[15]),
    .X(net204),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _354_ (.A(FrameStrobe[16]),
    .X(net205),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _355_ (.A(FrameStrobe[17]),
    .X(net206),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _356_ (.A(FrameStrobe[18]),
    .X(net207),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _357_ (.A(FrameStrobe[19]),
    .X(net208),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _358_ (.A(UserCLK),
    .X(net218),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _359_ (.A(\Inst_W_IO_switch_matrix.E1BEG0 ),
    .X(net118),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _360_ (.A(\Inst_W_IO_switch_matrix.E1BEG1 ),
    .X(net119),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _361_ (.A(\Inst_W_IO_switch_matrix.E1BEG2 ),
    .X(net120),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _362_ (.A(\Inst_W_IO_switch_matrix.E1BEG3 ),
    .X(net121),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _363_ (.A(\Inst_W_IO_switch_matrix.E2BEG0 ),
    .X(net122),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _364_ (.A(\Inst_W_IO_switch_matrix.E2BEG1 ),
    .X(net123),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout66 (.A(\Inst_W_IO_ConfigMem.Inst_frame0_bit25.Q ),
    .X(net66),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout67 (.A(\Inst_W_IO_ConfigMem.Inst_frame0_bit18.Q ),
    .X(net67),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout68 (.A(net70),
    .X(net68),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout69 (.A(net70),
    .X(net69),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout70 (.A(net71),
    .X(net70),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout71 (.A(FrameStrobe[3]),
    .X(net71),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout72 (.A(net75),
    .X(net72),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout73 (.A(net75),
    .X(net73),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout74 (.A(net75),
    .X(net74),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout75 (.A(net77),
    .X(net75),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout76 (.A(net77),
    .X(net76),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout77 (.A(FrameStrobe[2]),
    .X(net77),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout78 (.A(net79),
    .X(net78),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout79 (.A(net82),
    .X(net79),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout80 (.A(net82),
    .X(net80),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout81 (.A(net82),
    .X(net81),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout82 (.A(FrameStrobe[1]),
    .X(net82),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout83 (.A(net84),
    .X(net83),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout84 (.A(net88),
    .X(net84),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout85 (.A(net87),
    .X(net85),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout86 (.A(net87),
    .X(net86),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout87 (.A(net88),
    .X(net87),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout88 (.A(FrameStrobe[0]),
    .X(net88),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input1 (.A(A_O_top),
    .X(net1),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input2 (.A(B_O_top),
    .X(net2),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input3 (.A(FrameData[0]),
    .X(net3),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input4 (.A(FrameData[10]),
    .X(net4),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input5 (.A(FrameData[11]),
    .X(net5),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input6 (.A(FrameData[12]),
    .X(net6),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input7 (.A(FrameData[13]),
    .X(net7),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input8 (.A(FrameData[14]),
    .X(net8),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input9 (.A(FrameData[15]),
    .X(net9),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input10 (.A(FrameData[16]),
    .X(net10),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input11 (.A(FrameData[17]),
    .X(net11),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input12 (.A(FrameData[18]),
    .X(net12),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input13 (.A(FrameData[19]),
    .X(net13),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input14 (.A(FrameData[1]),
    .X(net14),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input15 (.A(FrameData[20]),
    .X(net15),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input16 (.A(FrameData[21]),
    .X(net16),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input17 (.A(FrameData[22]),
    .X(net17),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input18 (.A(FrameData[23]),
    .X(net18),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input19 (.A(FrameData[24]),
    .X(net19),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input20 (.A(FrameData[25]),
    .X(net20),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input21 (.A(FrameData[26]),
    .X(net21),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input22 (.A(FrameData[27]),
    .X(net22),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input23 (.A(FrameData[28]),
    .X(net23),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input24 (.A(FrameData[29]),
    .X(net24),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input25 (.A(FrameData[2]),
    .X(net25),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input26 (.A(FrameData[30]),
    .X(net26),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input27 (.A(FrameData[31]),
    .X(net27),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input28 (.A(FrameData[3]),
    .X(net28),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input29 (.A(FrameData[4]),
    .X(net29),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input30 (.A(FrameData[5]),
    .X(net30),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input31 (.A(FrameData[6]),
    .X(net31),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input32 (.A(FrameData[7]),
    .X(net32),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input33 (.A(FrameData[8]),
    .X(net33),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input34 (.A(FrameData[9]),
    .X(net34),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input35 (.A(W1END[0]),
    .X(net35),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input36 (.A(W1END[1]),
    .X(net36),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input37 (.A(W1END[2]),
    .X(net37),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input38 (.A(W1END[3]),
    .X(net38),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input39 (.A(W2END[0]),
    .X(net39),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input40 (.A(W2END[1]),
    .X(net40),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input41 (.A(W2END[2]),
    .X(net41),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input42 (.A(W2END[3]),
    .X(net42),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input43 (.A(W2END[4]),
    .X(net43),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input44 (.A(W2END[5]),
    .X(net44),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input45 (.A(W2END[6]),
    .X(net45),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input46 (.A(W2END[7]),
    .X(net46),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input47 (.A(W2MID[0]),
    .X(net47),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input48 (.A(W2MID[1]),
    .X(net48),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input49 (.A(W2MID[2]),
    .X(net49),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input50 (.A(W2MID[3]),
    .X(net50),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input51 (.A(W2MID[4]),
    .X(net51),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input52 (.A(W2MID[5]),
    .X(net52),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input53 (.A(W2MID[6]),
    .X(net53),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input54 (.A(W2MID[7]),
    .X(net54),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input55 (.A(W6END[0]),
    .X(net55),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input56 (.A(W6END[10]),
    .X(net56),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input57 (.A(W6END[11]),
    .X(net57),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input58 (.A(W6END[1]),
    .X(net58),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input59 (.A(W6END[2]),
    .X(net59),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input60 (.A(W6END[3]),
    .X(net60),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input61 (.A(W6END[4]),
    .X(net61),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input62 (.A(W6END[5]),
    .X(net62),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input63 (.A(W6END[6]),
    .X(net63),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input64 (.A(W6END[7]),
    .X(net64),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input65 (.A(W6END[8]),
    .X(net65),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input66 (.A(W6END[9]),
    .X(net89),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input67 (.A(WW4END[0]),
    .X(net90),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input68 (.A(WW4END[10]),
    .X(net91),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input69 (.A(WW4END[11]),
    .X(net92),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input70 (.A(WW4END[12]),
    .X(net93),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input71 (.A(WW4END[13]),
    .X(net94),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input72 (.A(WW4END[14]),
    .X(net95),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input73 (.A(WW4END[15]),
    .X(net96),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input74 (.A(WW4END[1]),
    .X(net97),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input75 (.A(WW4END[2]),
    .X(net98),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input76 (.A(WW4END[3]),
    .X(net99),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input77 (.A(WW4END[4]),
    .X(net100),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input78 (.A(WW4END[5]),
    .X(net101),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input79 (.A(WW4END[6]),
    .X(net102),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input80 (.A(WW4END[7]),
    .X(net103),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input81 (.A(WW4END[8]),
    .X(net104),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input82 (.A(WW4END[9]),
    .X(net105),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output83 (.A(net106),
    .X(A_I_top),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output84 (.A(net107),
    .X(A_T_top),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output85 (.A(net108),
    .X(A_config_C_bit0),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output86 (.A(net109),
    .X(A_config_C_bit1),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output87 (.A(net110),
    .X(A_config_C_bit2),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output88 (.A(net111),
    .X(A_config_C_bit3),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output89 (.A(net112),
    .X(B_I_top),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output90 (.A(net113),
    .X(B_T_top),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output91 (.A(net114),
    .X(B_config_C_bit0),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output92 (.A(net115),
    .X(B_config_C_bit1),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output93 (.A(net116),
    .X(B_config_C_bit2),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output94 (.A(net117),
    .X(B_config_C_bit3),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output95 (.A(net118),
    .X(E1BEG[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output96 (.A(net119),
    .X(E1BEG[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output97 (.A(net120),
    .X(E1BEG[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output98 (.A(net121),
    .X(E1BEG[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output99 (.A(net122),
    .X(E2BEG[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output100 (.A(net123),
    .X(E2BEG[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output101 (.A(net124),
    .X(E2BEG[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output102 (.A(net125),
    .X(E2BEG[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output103 (.A(net126),
    .X(E2BEG[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output104 (.A(net127),
    .X(E2BEG[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output105 (.A(net128),
    .X(E2BEG[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output106 (.A(net129),
    .X(E2BEG[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output107 (.A(net130),
    .X(E2BEGb[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output108 (.A(net131),
    .X(E2BEGb[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output109 (.A(net132),
    .X(E2BEGb[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output110 (.A(net133),
    .X(E2BEGb[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output111 (.A(net134),
    .X(E2BEGb[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output112 (.A(net135),
    .X(E2BEGb[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output113 (.A(net136),
    .X(E2BEGb[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output114 (.A(net137),
    .X(E2BEGb[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output115 (.A(net138),
    .X(E6BEG[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output116 (.A(net139),
    .X(E6BEG[10]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output117 (.A(net140),
    .X(E6BEG[11]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output118 (.A(net141),
    .X(E6BEG[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output119 (.A(net142),
    .X(E6BEG[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output120 (.A(net143),
    .X(E6BEG[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output121 (.A(net144),
    .X(E6BEG[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output122 (.A(net145),
    .X(E6BEG[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output123 (.A(net146),
    .X(E6BEG[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output124 (.A(net147),
    .X(E6BEG[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output125 (.A(net148),
    .X(E6BEG[8]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output126 (.A(net149),
    .X(E6BEG[9]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output127 (.A(net150),
    .X(EE4BEG[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output128 (.A(net151),
    .X(EE4BEG[10]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output129 (.A(net152),
    .X(EE4BEG[11]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output130 (.A(net153),
    .X(EE4BEG[12]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output131 (.A(net154),
    .X(EE4BEG[13]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output132 (.A(net155),
    .X(EE4BEG[14]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output133 (.A(net156),
    .X(EE4BEG[15]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output134 (.A(net157),
    .X(EE4BEG[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output135 (.A(net158),
    .X(EE4BEG[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output136 (.A(net159),
    .X(EE4BEG[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output137 (.A(net160),
    .X(EE4BEG[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output138 (.A(net161),
    .X(EE4BEG[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output139 (.A(net162),
    .X(EE4BEG[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output140 (.A(net163),
    .X(EE4BEG[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output141 (.A(net164),
    .X(EE4BEG[8]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output142 (.A(net165),
    .X(EE4BEG[9]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output143 (.A(net166),
    .X(FrameData_O[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output144 (.A(net167),
    .X(FrameData_O[10]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output145 (.A(net168),
    .X(FrameData_O[11]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output146 (.A(net169),
    .X(FrameData_O[12]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output147 (.A(net170),
    .X(FrameData_O[13]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output148 (.A(net171),
    .X(FrameData_O[14]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output149 (.A(net172),
    .X(FrameData_O[15]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output150 (.A(net173),
    .X(FrameData_O[16]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output151 (.A(net174),
    .X(FrameData_O[17]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output152 (.A(net175),
    .X(FrameData_O[18]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output153 (.A(net176),
    .X(FrameData_O[19]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output154 (.A(net177),
    .X(FrameData_O[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output155 (.A(net178),
    .X(FrameData_O[20]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output156 (.A(net179),
    .X(FrameData_O[21]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output157 (.A(net180),
    .X(FrameData_O[22]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output158 (.A(net181),
    .X(FrameData_O[23]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output159 (.A(net182),
    .X(FrameData_O[24]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output160 (.A(net183),
    .X(FrameData_O[25]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output161 (.A(net184),
    .X(FrameData_O[26]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output162 (.A(net185),
    .X(FrameData_O[27]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output163 (.A(net186),
    .X(FrameData_O[28]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output164 (.A(net187),
    .X(FrameData_O[29]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output165 (.A(net188),
    .X(FrameData_O[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output166 (.A(net189),
    .X(FrameData_O[30]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output167 (.A(net190),
    .X(FrameData_O[31]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output168 (.A(net191),
    .X(FrameData_O[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output169 (.A(net192),
    .X(FrameData_O[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output170 (.A(net193),
    .X(FrameData_O[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output171 (.A(net194),
    .X(FrameData_O[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output172 (.A(net195),
    .X(FrameData_O[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output173 (.A(net196),
    .X(FrameData_O[8]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output174 (.A(net197),
    .X(FrameData_O[9]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output175 (.A(net198),
    .X(FrameStrobe_O[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output176 (.A(net199),
    .X(FrameStrobe_O[10]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output177 (.A(net200),
    .X(FrameStrobe_O[11]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output178 (.A(net201),
    .X(FrameStrobe_O[12]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output179 (.A(net202),
    .X(FrameStrobe_O[13]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output180 (.A(net203),
    .X(FrameStrobe_O[14]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output181 (.A(net204),
    .X(FrameStrobe_O[15]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output182 (.A(net205),
    .X(FrameStrobe_O[16]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output183 (.A(net206),
    .X(FrameStrobe_O[17]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output184 (.A(net207),
    .X(FrameStrobe_O[18]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output185 (.A(net208),
    .X(FrameStrobe_O[19]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output186 (.A(net209),
    .X(FrameStrobe_O[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output187 (.A(net210),
    .X(FrameStrobe_O[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output188 (.A(net211),
    .X(FrameStrobe_O[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output189 (.A(net212),
    .X(FrameStrobe_O[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output190 (.A(net213),
    .X(FrameStrobe_O[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output191 (.A(net214),
    .X(FrameStrobe_O[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output192 (.A(net215),
    .X(FrameStrobe_O[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output193 (.A(net216),
    .X(FrameStrobe_O[8]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output194 (.A(net217),
    .X(FrameStrobe_O[9]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output195 (.A(net218),
    .X(UserCLKo),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_tiehi _260__196 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net219));
 sg13g2_decap_8 FILLER_0_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_45 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_52 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_59 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_64 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_64 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_66 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_92 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_43 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_50 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_90 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_97 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_29 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_52 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_78 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_36 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_86 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_20 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_66 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_73 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_114 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_30 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_37 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_55 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_62 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_22 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_26 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_50 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_90 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_92 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_114 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_37 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_48 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_50 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_73 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_30 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_79 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_6 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_41 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_43 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_90 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_114 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_37 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_34 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_36 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_41 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_43 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_24 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_55 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_27 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_34 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_41 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_48 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_55 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_90 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_34 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_58 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_64 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_65 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_79 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_79 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_15 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_55 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_62 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_29 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_64 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_9 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_27 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_38 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_45 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_52 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_15 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_86 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_38 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_86 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_13 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_31 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_38 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_45 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_52 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_16 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_37 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_41 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_51 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_15 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_64 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_65 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_27 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_29 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_59 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_66 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_73 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_80 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_114 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_71 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_78 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_29 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_90 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_50_97 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_50_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_51_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_51_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_52_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_52_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_53_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_54_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_54_114 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_55_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_79 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_86 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_55_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_55_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_56_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_56_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_57_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_37 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_48 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_55 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_62 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_69 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_57_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_57_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_57_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_57_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_57_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_15 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_22 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_29 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_36 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_43 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_50 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_64 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_71 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_78 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_58_92 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_58_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_59_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_59_9 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_59_15 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_59_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_59_27 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_59_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_59_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_59_45 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_59_51 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_59_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_59_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_59_69 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_59_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_59_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_59_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_59_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_59_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_59_105 (.VDD(VPWR),
    .VSS(VGND));
endmodule
