module S_CPU_IRQ (Co,
    IRQ_top0,
    IRQ_top1,
    IRQ_top2,
    IRQ_top3,
    UserCLK,
    UserCLKo,
    FrameData,
    FrameData_O,
    FrameStrobe,
    FrameStrobe_O,
    N1BEG,
    N2BEG,
    N2BEGb,
    N4BEG,
    NN4BEG,
    S1END,
    S2END,
    S2MID,
    S4END,
    SS4END);
 output Co;
 output IRQ_top0;
 output IRQ_top1;
 output IRQ_top2;
 output IRQ_top3;
 input UserCLK;
 output UserCLKo;
 input [31:0] FrameData;
 output [31:0] FrameData_O;
 input [19:0] FrameStrobe;
 output [19:0] FrameStrobe_O;
 output [3:0] N1BEG;
 output [7:0] N2BEG;
 output [7:0] N2BEGb;
 output [15:0] N4BEG;
 output [15:0] NN4BEG;
 input [3:0] S1END;
 input [7:0] S2END;
 input [7:0] S2MID;
 input [15:0] S4END;
 input [15:0] SS4END;

 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire \Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit20.Q ;
 wire \Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit21.Q ;
 wire \Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit22.Q ;
 wire \Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit23.Q ;
 wire \Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit24.Q ;
 wire \Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit25.Q ;
 wire \Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit26.Q ;
 wire \Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit27.Q ;
 wire \Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit28.Q ;
 wire \Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit29.Q ;
 wire \Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit30.Q ;
 wire \Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit31.Q ;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire net3;
 wire net1;
 wire net2;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net156;

 sky130_fd_sc_hd__inv_2 _024_ (.A(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit31.Q ),
    .Y(_000_));
 sky130_fd_sc_hd__inv_2 _025_ (.A(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit28.Q ),
    .Y(_001_));
 sky130_fd_sc_hd__inv_2 _026_ (.A(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit25.Q ),
    .Y(_002_));
 sky130_fd_sc_hd__inv_2 _027_ (.A(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit22.Q ),
    .Y(_003_));
 sky130_fd_sc_hd__mux4_1 _028_ (.A0(net34),
    .A1(net38),
    .A2(net42),
    .A3(net46),
    .S0(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit29.Q ),
    .S1(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit30.Q ),
    .X(_004_));
 sky130_fd_sc_hd__nand2b_1 _029_ (.A_N(net30),
    .B(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit29.Q ),
    .Y(_005_));
 sky130_fd_sc_hd__o21ba_1 _030_ (.A1(net18),
    .A2(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit29.Q ),
    .B1_N(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit30.Q ),
    .X(_006_));
 sky130_fd_sc_hd__mux2_1 _031_ (.A0(net22),
    .A1(net26),
    .S(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit29.Q ),
    .X(_007_));
 sky130_fd_sc_hd__a221o_1 _032_ (.A1(_005_),
    .A2(_006_),
    .B1(_007_),
    .B2(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit30.Q ),
    .C1(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit31.Q ),
    .X(_008_));
 sky130_fd_sc_hd__o21a_1 _033_ (.A1(_000_),
    .A2(_004_),
    .B1(_008_),
    .X(net102));
 sky130_fd_sc_hd__mux4_1 _034_ (.A0(net33),
    .A1(net37),
    .A2(net41),
    .A3(net45),
    .S0(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit26.Q ),
    .S1(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit27.Q ),
    .X(_009_));
 sky130_fd_sc_hd__nand2b_1 _035_ (.A_N(net29),
    .B(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit26.Q ),
    .Y(_010_));
 sky130_fd_sc_hd__o21ba_1 _036_ (.A1(net17),
    .A2(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit26.Q ),
    .B1_N(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit27.Q ),
    .X(_011_));
 sky130_fd_sc_hd__mux2_1 _037_ (.A0(net21),
    .A1(net25),
    .S(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit26.Q ),
    .X(_012_));
 sky130_fd_sc_hd__a221o_1 _038_ (.A1(_010_),
    .A2(_011_),
    .B1(_012_),
    .B2(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit27.Q ),
    .C1(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit28.Q ),
    .X(_013_));
 sky130_fd_sc_hd__o21a_1 _039_ (.A1(_001_),
    .A2(_009_),
    .B1(_013_),
    .X(net101));
 sky130_fd_sc_hd__mux4_1 _040_ (.A0(net32),
    .A1(net36),
    .A2(net40),
    .A3(net44),
    .S0(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit23.Q ),
    .S1(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit24.Q ),
    .X(_014_));
 sky130_fd_sc_hd__nand2b_1 _041_ (.A_N(net28),
    .B(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit23.Q ),
    .Y(_015_));
 sky130_fd_sc_hd__o21ba_1 _042_ (.A1(net16),
    .A2(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit23.Q ),
    .B1_N(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit24.Q ),
    .X(_016_));
 sky130_fd_sc_hd__mux2_1 _043_ (.A0(net20),
    .A1(net24),
    .S(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit23.Q ),
    .X(_017_));
 sky130_fd_sc_hd__a221o_1 _044_ (.A1(_015_),
    .A2(_016_),
    .B1(_017_),
    .B2(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit24.Q ),
    .C1(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit25.Q ),
    .X(_018_));
 sky130_fd_sc_hd__o21a_1 _045_ (.A1(_002_),
    .A2(_014_),
    .B1(_018_),
    .X(net100));
 sky130_fd_sc_hd__mux4_1 _046_ (.A0(net31),
    .A1(net35),
    .A2(net39),
    .A3(net43),
    .S0(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit20.Q ),
    .S1(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit21.Q ),
    .X(_019_));
 sky130_fd_sc_hd__nand2b_1 _047_ (.A_N(net27),
    .B(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit20.Q ),
    .Y(_020_));
 sky130_fd_sc_hd__o21ba_1 _048_ (.A1(net15),
    .A2(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit20.Q ),
    .B1_N(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit21.Q ),
    .X(_021_));
 sky130_fd_sc_hd__mux2_1 _049_ (.A0(net19),
    .A1(net23),
    .S(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit20.Q ),
    .X(_022_));
 sky130_fd_sc_hd__a221o_1 _050_ (.A1(_020_),
    .A2(_021_),
    .B1(_022_),
    .B2(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit21.Q ),
    .C1(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit22.Q ),
    .X(_023_));
 sky130_fd_sc_hd__o21a_1 _051_ (.A1(_003_),
    .A2(_019_),
    .B1(_023_),
    .X(net99));
 sky130_fd_sc_hd__dlxtp_1 _052_ (.D(net1),
    .GATE(net3),
    .Q(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _053_ (.D(net2),
    .GATE(net3),
    .Q(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _054_ (.D(net4),
    .GATE(net3),
    .Q(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _055_ (.D(net5),
    .GATE(net3),
    .Q(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _056_ (.D(net6),
    .GATE(net3),
    .Q(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _057_ (.D(net7),
    .GATE(net3),
    .Q(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _058_ (.D(net8),
    .GATE(net3),
    .Q(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _059_ (.D(net9),
    .GATE(net3),
    .Q(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _060_ (.D(net10),
    .GATE(net3),
    .Q(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _061_ (.D(net11),
    .GATE(net3),
    .Q(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _062_ (.D(net12),
    .GATE(net14),
    .Q(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _063_ (.D(net13),
    .GATE(net14),
    .Q(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit31.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(FrameData[0]));
 sky130_fd_sc_hd__clkbuf_1 _065_ (.A(FrameData[0]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_2 _066_ (.A(FrameData[1]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_1 _067_ (.A(FrameData[2]),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_1 _068_ (.A(FrameData[3]),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_1 _069_ (.A(FrameData[4]),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_2 _070_ (.A(FrameData[5]),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_2 _071_ (.A(FrameData[6]),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_2 _072_ (.A(FrameData[7]),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_2 _073_ (.A(FrameData[8]),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_2 _074_ (.A(FrameData[9]),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_2 _075_ (.A(FrameData[10]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_2 _076_ (.A(FrameData[11]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_1 _077_ (.A(FrameData[12]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_2 _078_ (.A(FrameData[13]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_1 _079_ (.A(FrameData[14]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_1 _080_ (.A(FrameData[15]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_2 _081_ (.A(FrameData[16]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_2 _082_ (.A(FrameData[17]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_2 _083_ (.A(FrameData[18]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_1 _084_ (.A(FrameData[19]),
    .X(net57));
 sky130_fd_sc_hd__buf_1 _085_ (.A(net1),
    .X(net59));
 sky130_fd_sc_hd__buf_1 _086_ (.A(net2),
    .X(net60));
 sky130_fd_sc_hd__buf_1 _087_ (.A(net4),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_2 _088_ (.A(net5),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_2 _089_ (.A(net6),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_2 _090_ (.A(net7),
    .X(net64));
 sky130_fd_sc_hd__buf_1 _091_ (.A(net8),
    .X(net65));
 sky130_fd_sc_hd__buf_1 _092_ (.A(net9),
    .X(net66));
 sky130_fd_sc_hd__buf_1 _093_ (.A(net10),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_2 _094_ (.A(net11),
    .X(net68));
 sky130_fd_sc_hd__buf_1 _095_ (.A(net12),
    .X(net70));
 sky130_fd_sc_hd__buf_1 _096_ (.A(net13),
    .X(net71));
 sky130_fd_sc_hd__buf_1 _097_ (.A(net14),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_1 _098_ (.A(FrameStrobe[1]),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_1 _099_ (.A(FrameStrobe[2]),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_1 _100_ (.A(FrameStrobe[3]),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_1 _101_ (.A(FrameStrobe[4]),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_1 _102_ (.A(FrameStrobe[5]),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_1 _103_ (.A(FrameStrobe[6]),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_1 _104_ (.A(FrameStrobe[7]),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_1 _105_ (.A(FrameStrobe[8]),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_1 _106_ (.A(FrameStrobe[9]),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_1 _107_ (.A(FrameStrobe[10]),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_1 _108_ (.A(FrameStrobe[11]),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_1 _109_ (.A(FrameStrobe[12]),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_1 _110_ (.A(FrameStrobe[13]),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_1 _111_ (.A(FrameStrobe[14]),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_1 _112_ (.A(FrameStrobe[15]),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_1 _113_ (.A(FrameStrobe[16]),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_1 _114_ (.A(FrameStrobe[17]),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_1 _115_ (.A(FrameStrobe[18]),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_1 _116_ (.A(FrameStrobe[19]),
    .X(net89));
 sky130_fd_sc_hd__buf_1 _117_ (.A(net18),
    .X(net103));
 sky130_fd_sc_hd__buf_1 _118_ (.A(net17),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_1 _119_ (.A(net16),
    .X(net105));
 sky130_fd_sc_hd__buf_1 _120_ (.A(net15),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_1 _121_ (.A(S2MID[7]),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_1 _122_ (.A(S2MID[6]),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_1 _123_ (.A(S2MID[5]),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_1 _124_ (.A(S2MID[4]),
    .X(net110));
 sky130_fd_sc_hd__buf_1 _125_ (.A(net30),
    .X(net111));
 sky130_fd_sc_hd__buf_1 _126_ (.A(net29),
    .X(net112));
 sky130_fd_sc_hd__clkbuf_1 _127_ (.A(net28),
    .X(net113));
 sky130_fd_sc_hd__buf_1 _128_ (.A(net27),
    .X(net114));
 sky130_fd_sc_hd__buf_1 _129_ (.A(net26),
    .X(net115));
 sky130_fd_sc_hd__buf_1 _130_ (.A(net25),
    .X(net116));
 sky130_fd_sc_hd__clkbuf_1 _131_ (.A(net24),
    .X(net117));
 sky130_fd_sc_hd__clkbuf_1 _132_ (.A(net23),
    .X(net118));
 sky130_fd_sc_hd__buf_1 _133_ (.A(net22),
    .X(net119));
 sky130_fd_sc_hd__clkbuf_1 _134_ (.A(net21),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_1 _135_ (.A(net20),
    .X(net121));
 sky130_fd_sc_hd__buf_1 _136_ (.A(net19),
    .X(net122));
 sky130_fd_sc_hd__buf_1 _137_ (.A(S4END[15]),
    .X(net123));
 sky130_fd_sc_hd__buf_1 _138_ (.A(S4END[14]),
    .X(net130));
 sky130_fd_sc_hd__buf_1 _139_ (.A(S4END[13]),
    .X(net131));
 sky130_fd_sc_hd__buf_1 _140_ (.A(S4END[12]),
    .X(net132));
 sky130_fd_sc_hd__buf_1 _141_ (.A(S4END[11]),
    .X(net133));
 sky130_fd_sc_hd__buf_1 _142_ (.A(S4END[10]),
    .X(net134));
 sky130_fd_sc_hd__buf_1 _143_ (.A(S4END[9]),
    .X(net135));
 sky130_fd_sc_hd__buf_1 _144_ (.A(S4END[8]),
    .X(net136));
 sky130_fd_sc_hd__buf_1 _145_ (.A(net38),
    .X(net137));
 sky130_fd_sc_hd__clkbuf_1 _146_ (.A(net37),
    .X(net138));
 sky130_fd_sc_hd__clkbuf_1 _147_ (.A(net36),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_1 _148_ (.A(net35),
    .X(net125));
 sky130_fd_sc_hd__buf_1 _149_ (.A(net34),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_1 _150_ (.A(net33),
    .X(net127));
 sky130_fd_sc_hd__clkbuf_1 _151_ (.A(net32),
    .X(net128));
 sky130_fd_sc_hd__clkbuf_1 _152_ (.A(net31),
    .X(net129));
 sky130_fd_sc_hd__buf_1 _153_ (.A(SS4END[15]),
    .X(net139));
 sky130_fd_sc_hd__buf_1 _154_ (.A(SS4END[14]),
    .X(net146));
 sky130_fd_sc_hd__buf_1 _155_ (.A(SS4END[13]),
    .X(net147));
 sky130_fd_sc_hd__buf_1 _156_ (.A(SS4END[12]),
    .X(net148));
 sky130_fd_sc_hd__buf_1 _157_ (.A(SS4END[11]),
    .X(net149));
 sky130_fd_sc_hd__buf_1 _158_ (.A(SS4END[10]),
    .X(net150));
 sky130_fd_sc_hd__buf_1 _159_ (.A(SS4END[9]),
    .X(net151));
 sky130_fd_sc_hd__buf_1 _160_ (.A(SS4END[8]),
    .X(net152));
 sky130_fd_sc_hd__clkbuf_1 _161_ (.A(net46),
    .X(net153));
 sky130_fd_sc_hd__clkbuf_1 _162_ (.A(net45),
    .X(net154));
 sky130_fd_sc_hd__buf_1 _163_ (.A(net44),
    .X(net140));
 sky130_fd_sc_hd__clkbuf_1 _164_ (.A(net43),
    .X(net141));
 sky130_fd_sc_hd__clkbuf_1 _165_ (.A(net42),
    .X(net142));
 sky130_fd_sc_hd__clkbuf_1 _166_ (.A(net41),
    .X(net143));
 sky130_fd_sc_hd__buf_1 _167_ (.A(net40),
    .X(net144));
 sky130_fd_sc_hd__clkbuf_1 _168_ (.A(net39),
    .X(net145));
 sky130_fd_sc_hd__buf_2 _169_ (.A(UserCLK),
    .X(net155));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_121 ();
 sky130_fd_sc_hd__clkbuf_2 fanout3 (.A(net14),
    .X(net3));
 sky130_fd_sc_hd__buf_1 input1 (.A(FrameData[20]),
    .X(net1));
 sky130_fd_sc_hd__buf_1 input2 (.A(FrameData[21]),
    .X(net2));
 sky130_fd_sc_hd__buf_1 input3 (.A(FrameData[22]),
    .X(net4));
 sky130_fd_sc_hd__buf_1 input4 (.A(FrameData[23]),
    .X(net5));
 sky130_fd_sc_hd__buf_1 input5 (.A(FrameData[24]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(FrameData[25]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(FrameData[26]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(FrameData[27]),
    .X(net9));
 sky130_fd_sc_hd__buf_1 input9 (.A(FrameData[28]),
    .X(net10));
 sky130_fd_sc_hd__buf_1 input10 (.A(FrameData[29]),
    .X(net11));
 sky130_fd_sc_hd__buf_1 input11 (.A(FrameData[30]),
    .X(net12));
 sky130_fd_sc_hd__buf_1 input12 (.A(FrameData[31]),
    .X(net13));
 sky130_fd_sc_hd__dlymetal6s2s_1 input13 (.A(FrameStrobe[0]),
    .X(net14));
 sky130_fd_sc_hd__buf_1 input14 (.A(S1END[0]),
    .X(net15));
 sky130_fd_sc_hd__buf_1 input15 (.A(S1END[1]),
    .X(net16));
 sky130_fd_sc_hd__buf_1 input16 (.A(S1END[2]),
    .X(net17));
 sky130_fd_sc_hd__buf_1 input17 (.A(S1END[3]),
    .X(net18));
 sky130_fd_sc_hd__buf_1 input18 (.A(S2END[0]),
    .X(net19));
 sky130_fd_sc_hd__buf_1 input19 (.A(S2END[1]),
    .X(net20));
 sky130_fd_sc_hd__buf_1 input20 (.A(S2END[2]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(S2END[3]),
    .X(net22));
 sky130_fd_sc_hd__buf_1 input22 (.A(S2END[4]),
    .X(net23));
 sky130_fd_sc_hd__buf_1 input23 (.A(S2END[5]),
    .X(net24));
 sky130_fd_sc_hd__buf_1 input24 (.A(S2END[6]),
    .X(net25));
 sky130_fd_sc_hd__buf_1 input25 (.A(S2END[7]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(S2MID[0]),
    .X(net27));
 sky130_fd_sc_hd__buf_1 input27 (.A(S2MID[1]),
    .X(net28));
 sky130_fd_sc_hd__buf_1 input28 (.A(S2MID[2]),
    .X(net29));
 sky130_fd_sc_hd__buf_1 input29 (.A(S2MID[3]),
    .X(net30));
 sky130_fd_sc_hd__buf_1 input30 (.A(S4END[0]),
    .X(net31));
 sky130_fd_sc_hd__buf_1 input31 (.A(S4END[1]),
    .X(net32));
 sky130_fd_sc_hd__buf_1 input32 (.A(S4END[2]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 input33 (.A(S4END[3]),
    .X(net34));
 sky130_fd_sc_hd__buf_1 input34 (.A(S4END[4]),
    .X(net35));
 sky130_fd_sc_hd__buf_1 input35 (.A(S4END[5]),
    .X(net36));
 sky130_fd_sc_hd__buf_1 input36 (.A(S4END[6]),
    .X(net37));
 sky130_fd_sc_hd__buf_1 input37 (.A(S4END[7]),
    .X(net38));
 sky130_fd_sc_hd__buf_1 input38 (.A(SS4END[0]),
    .X(net39));
 sky130_fd_sc_hd__dlymetal6s2s_1 input39 (.A(SS4END[1]),
    .X(net40));
 sky130_fd_sc_hd__buf_1 input40 (.A(SS4END[2]),
    .X(net41));
 sky130_fd_sc_hd__buf_1 input41 (.A(SS4END[3]),
    .X(net42));
 sky130_fd_sc_hd__buf_1 input42 (.A(SS4END[4]),
    .X(net43));
 sky130_fd_sc_hd__dlymetal6s2s_1 input43 (.A(SS4END[5]),
    .X(net44));
 sky130_fd_sc_hd__buf_1 input44 (.A(SS4END[6]),
    .X(net45));
 sky130_fd_sc_hd__buf_1 input45 (.A(SS4END[7]),
    .X(net46));
 sky130_fd_sc_hd__buf_2 output46 (.A(net47),
    .X(FrameData_O[0]));
 sky130_fd_sc_hd__buf_2 output47 (.A(net48),
    .X(FrameData_O[10]));
 sky130_fd_sc_hd__buf_2 output48 (.A(net49),
    .X(FrameData_O[11]));
 sky130_fd_sc_hd__buf_2 output49 (.A(net50),
    .X(FrameData_O[12]));
 sky130_fd_sc_hd__buf_2 output50 (.A(net51),
    .X(FrameData_O[13]));
 sky130_fd_sc_hd__buf_2 output51 (.A(net52),
    .X(FrameData_O[14]));
 sky130_fd_sc_hd__buf_2 output52 (.A(net53),
    .X(FrameData_O[15]));
 sky130_fd_sc_hd__buf_2 output53 (.A(net54),
    .X(FrameData_O[16]));
 sky130_fd_sc_hd__buf_2 output54 (.A(net55),
    .X(FrameData_O[17]));
 sky130_fd_sc_hd__buf_2 output55 (.A(net56),
    .X(FrameData_O[18]));
 sky130_fd_sc_hd__buf_2 output56 (.A(net57),
    .X(FrameData_O[19]));
 sky130_fd_sc_hd__buf_2 output57 (.A(net58),
    .X(FrameData_O[1]));
 sky130_fd_sc_hd__buf_2 output58 (.A(net59),
    .X(FrameData_O[20]));
 sky130_fd_sc_hd__buf_2 output59 (.A(net60),
    .X(FrameData_O[21]));
 sky130_fd_sc_hd__buf_2 output60 (.A(net61),
    .X(FrameData_O[22]));
 sky130_fd_sc_hd__buf_2 output61 (.A(net62),
    .X(FrameData_O[23]));
 sky130_fd_sc_hd__buf_2 output62 (.A(net63),
    .X(FrameData_O[24]));
 sky130_fd_sc_hd__buf_2 output63 (.A(net64),
    .X(FrameData_O[25]));
 sky130_fd_sc_hd__buf_2 output64 (.A(net65),
    .X(FrameData_O[26]));
 sky130_fd_sc_hd__buf_2 output65 (.A(net66),
    .X(FrameData_O[27]));
 sky130_fd_sc_hd__buf_2 output66 (.A(net67),
    .X(FrameData_O[28]));
 sky130_fd_sc_hd__buf_2 output67 (.A(net68),
    .X(FrameData_O[29]));
 sky130_fd_sc_hd__buf_2 output68 (.A(net69),
    .X(FrameData_O[2]));
 sky130_fd_sc_hd__buf_2 output69 (.A(net70),
    .X(FrameData_O[30]));
 sky130_fd_sc_hd__buf_2 output70 (.A(net71),
    .X(FrameData_O[31]));
 sky130_fd_sc_hd__buf_2 output71 (.A(net72),
    .X(FrameData_O[3]));
 sky130_fd_sc_hd__buf_2 output72 (.A(net73),
    .X(FrameData_O[4]));
 sky130_fd_sc_hd__buf_2 output73 (.A(net74),
    .X(FrameData_O[5]));
 sky130_fd_sc_hd__buf_2 output74 (.A(net75),
    .X(FrameData_O[6]));
 sky130_fd_sc_hd__buf_2 output75 (.A(net76),
    .X(FrameData_O[7]));
 sky130_fd_sc_hd__buf_2 output76 (.A(net77),
    .X(FrameData_O[8]));
 sky130_fd_sc_hd__buf_2 output77 (.A(net78),
    .X(FrameData_O[9]));
 sky130_fd_sc_hd__buf_2 output78 (.A(net79),
    .X(FrameStrobe_O[0]));
 sky130_fd_sc_hd__buf_2 output79 (.A(net80),
    .X(FrameStrobe_O[10]));
 sky130_fd_sc_hd__buf_2 output80 (.A(net81),
    .X(FrameStrobe_O[11]));
 sky130_fd_sc_hd__buf_2 output81 (.A(net82),
    .X(FrameStrobe_O[12]));
 sky130_fd_sc_hd__buf_2 output82 (.A(net83),
    .X(FrameStrobe_O[13]));
 sky130_fd_sc_hd__buf_2 output83 (.A(net84),
    .X(FrameStrobe_O[14]));
 sky130_fd_sc_hd__buf_2 output84 (.A(net85),
    .X(FrameStrobe_O[15]));
 sky130_fd_sc_hd__buf_2 output85 (.A(net86),
    .X(FrameStrobe_O[16]));
 sky130_fd_sc_hd__buf_2 output86 (.A(net87),
    .X(FrameStrobe_O[17]));
 sky130_fd_sc_hd__buf_2 output87 (.A(net88),
    .X(FrameStrobe_O[18]));
 sky130_fd_sc_hd__buf_2 output88 (.A(net89),
    .X(FrameStrobe_O[19]));
 sky130_fd_sc_hd__buf_2 output89 (.A(net90),
    .X(FrameStrobe_O[1]));
 sky130_fd_sc_hd__buf_2 output90 (.A(net91),
    .X(FrameStrobe_O[2]));
 sky130_fd_sc_hd__buf_2 output91 (.A(net92),
    .X(FrameStrobe_O[3]));
 sky130_fd_sc_hd__buf_2 output92 (.A(net93),
    .X(FrameStrobe_O[4]));
 sky130_fd_sc_hd__buf_2 output93 (.A(net94),
    .X(FrameStrobe_O[5]));
 sky130_fd_sc_hd__buf_2 output94 (.A(net95),
    .X(FrameStrobe_O[6]));
 sky130_fd_sc_hd__buf_2 output95 (.A(net96),
    .X(FrameStrobe_O[7]));
 sky130_fd_sc_hd__buf_2 output96 (.A(net97),
    .X(FrameStrobe_O[8]));
 sky130_fd_sc_hd__buf_2 output97 (.A(net98),
    .X(FrameStrobe_O[9]));
 sky130_fd_sc_hd__buf_2 output98 (.A(net99),
    .X(IRQ_top0));
 sky130_fd_sc_hd__buf_2 output99 (.A(net100),
    .X(IRQ_top1));
 sky130_fd_sc_hd__buf_2 output100 (.A(net101),
    .X(IRQ_top2));
 sky130_fd_sc_hd__buf_2 output101 (.A(net102),
    .X(IRQ_top3));
 sky130_fd_sc_hd__buf_2 output102 (.A(net103),
    .X(N1BEG[0]));
 sky130_fd_sc_hd__buf_2 output103 (.A(net104),
    .X(N1BEG[1]));
 sky130_fd_sc_hd__buf_2 output104 (.A(net105),
    .X(N1BEG[2]));
 sky130_fd_sc_hd__buf_2 output105 (.A(net106),
    .X(N1BEG[3]));
 sky130_fd_sc_hd__buf_2 output106 (.A(net107),
    .X(N2BEG[0]));
 sky130_fd_sc_hd__buf_2 output107 (.A(net108),
    .X(N2BEG[1]));
 sky130_fd_sc_hd__buf_2 output108 (.A(net109),
    .X(N2BEG[2]));
 sky130_fd_sc_hd__buf_2 output109 (.A(net110),
    .X(N2BEG[3]));
 sky130_fd_sc_hd__buf_2 output110 (.A(net111),
    .X(N2BEG[4]));
 sky130_fd_sc_hd__buf_2 output111 (.A(net112),
    .X(N2BEG[5]));
 sky130_fd_sc_hd__buf_2 output112 (.A(net113),
    .X(N2BEG[6]));
 sky130_fd_sc_hd__buf_2 output113 (.A(net114),
    .X(N2BEG[7]));
 sky130_fd_sc_hd__buf_2 output114 (.A(net115),
    .X(N2BEGb[0]));
 sky130_fd_sc_hd__buf_2 output115 (.A(net116),
    .X(N2BEGb[1]));
 sky130_fd_sc_hd__buf_2 output116 (.A(net117),
    .X(N2BEGb[2]));
 sky130_fd_sc_hd__buf_2 output117 (.A(net118),
    .X(N2BEGb[3]));
 sky130_fd_sc_hd__buf_2 output118 (.A(net119),
    .X(N2BEGb[4]));
 sky130_fd_sc_hd__buf_2 output119 (.A(net120),
    .X(N2BEGb[5]));
 sky130_fd_sc_hd__buf_2 output120 (.A(net121),
    .X(N2BEGb[6]));
 sky130_fd_sc_hd__buf_2 output121 (.A(net122),
    .X(N2BEGb[7]));
 sky130_fd_sc_hd__buf_2 output122 (.A(net123),
    .X(N4BEG[0]));
 sky130_fd_sc_hd__buf_2 output123 (.A(net124),
    .X(N4BEG[10]));
 sky130_fd_sc_hd__buf_2 output124 (.A(net125),
    .X(N4BEG[11]));
 sky130_fd_sc_hd__buf_2 output125 (.A(net126),
    .X(N4BEG[12]));
 sky130_fd_sc_hd__buf_2 output126 (.A(net127),
    .X(N4BEG[13]));
 sky130_fd_sc_hd__buf_2 output127 (.A(net128),
    .X(N4BEG[14]));
 sky130_fd_sc_hd__buf_2 output128 (.A(net129),
    .X(N4BEG[15]));
 sky130_fd_sc_hd__buf_2 output129 (.A(net130),
    .X(N4BEG[1]));
 sky130_fd_sc_hd__buf_2 output130 (.A(net131),
    .X(N4BEG[2]));
 sky130_fd_sc_hd__buf_2 output131 (.A(net132),
    .X(N4BEG[3]));
 sky130_fd_sc_hd__buf_2 output132 (.A(net133),
    .X(N4BEG[4]));
 sky130_fd_sc_hd__buf_2 output133 (.A(net134),
    .X(N4BEG[5]));
 sky130_fd_sc_hd__buf_2 output134 (.A(net135),
    .X(N4BEG[6]));
 sky130_fd_sc_hd__buf_2 output135 (.A(net136),
    .X(N4BEG[7]));
 sky130_fd_sc_hd__buf_2 output136 (.A(net137),
    .X(N4BEG[8]));
 sky130_fd_sc_hd__buf_2 output137 (.A(net138),
    .X(N4BEG[9]));
 sky130_fd_sc_hd__buf_2 output138 (.A(net139),
    .X(NN4BEG[0]));
 sky130_fd_sc_hd__buf_2 output139 (.A(net140),
    .X(NN4BEG[10]));
 sky130_fd_sc_hd__buf_2 output140 (.A(net141),
    .X(NN4BEG[11]));
 sky130_fd_sc_hd__buf_2 output141 (.A(net142),
    .X(NN4BEG[12]));
 sky130_fd_sc_hd__buf_2 output142 (.A(net143),
    .X(NN4BEG[13]));
 sky130_fd_sc_hd__buf_2 output143 (.A(net144),
    .X(NN4BEG[14]));
 sky130_fd_sc_hd__buf_2 output144 (.A(net145),
    .X(NN4BEG[15]));
 sky130_fd_sc_hd__buf_2 output145 (.A(net146),
    .X(NN4BEG[1]));
 sky130_fd_sc_hd__buf_2 output146 (.A(net147),
    .X(NN4BEG[2]));
 sky130_fd_sc_hd__buf_2 output147 (.A(net148),
    .X(NN4BEG[3]));
 sky130_fd_sc_hd__buf_2 output148 (.A(net149),
    .X(NN4BEG[4]));
 sky130_fd_sc_hd__buf_2 output149 (.A(net150),
    .X(NN4BEG[5]));
 sky130_fd_sc_hd__buf_2 output150 (.A(net151),
    .X(NN4BEG[6]));
 sky130_fd_sc_hd__buf_2 output151 (.A(net152),
    .X(NN4BEG[7]));
 sky130_fd_sc_hd__buf_2 output152 (.A(net153),
    .X(NN4BEG[8]));
 sky130_fd_sc_hd__buf_2 output153 (.A(net154),
    .X(NN4BEG[9]));
 sky130_fd_sc_hd__buf_1 output154 (.A(net155),
    .X(UserCLKo));
 sky130_fd_sc_hd__conb_1 S_CPU_IRQ_155 (.LO(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(FrameData[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(FrameData[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(FrameData[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(FrameData[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(FrameData[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(FrameData[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(FrameStrobe[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(FrameStrobe[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(FrameStrobe[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(FrameStrobe[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(S2MID[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(FrameStrobe[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(net148));
 sky130_fd_sc_hd__fill_2 FILLER_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_144 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_56 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_409 ();
 assign Co = net156;
endmodule
