* NGSPICE file created from S_EF_DAC8.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlxtp_1 abstract view
.subckt sky130_fd_sc_hd__dlxtp_1 D GATE VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

.subckt S_EF_DAC8 Co FrameData[0] FrameData[10] FrameData[11] FrameData[12] FrameData[13]
+ FrameData[14] FrameData[15] FrameData[16] FrameData[17] FrameData[18] FrameData[19]
+ FrameData[1] FrameData[20] FrameData[21] FrameData[22] FrameData[23] FrameData[24]
+ FrameData[25] FrameData[26] FrameData[27] FrameData[28] FrameData[29] FrameData[2]
+ FrameData[30] FrameData[31] FrameData[3] FrameData[4] FrameData[5] FrameData[6]
+ FrameData[7] FrameData[8] FrameData[9] FrameData_O[0] FrameData_O[10] FrameData_O[11]
+ FrameData_O[12] FrameData_O[13] FrameData_O[14] FrameData_O[15] FrameData_O[16]
+ FrameData_O[17] FrameData_O[18] FrameData_O[19] FrameData_O[1] FrameData_O[20] FrameData_O[21]
+ FrameData_O[22] FrameData_O[23] FrameData_O[24] FrameData_O[25] FrameData_O[26]
+ FrameData_O[27] FrameData_O[28] FrameData_O[29] FrameData_O[2] FrameData_O[30] FrameData_O[31]
+ FrameData_O[3] FrameData_O[4] FrameData_O[5] FrameData_O[6] FrameData_O[7] FrameData_O[8]
+ FrameData_O[9] FrameStrobe[0] FrameStrobe[10] FrameStrobe[11] FrameStrobe[12] FrameStrobe[13]
+ FrameStrobe[14] FrameStrobe[15] FrameStrobe[16] FrameStrobe[17] FrameStrobe[18]
+ FrameStrobe[19] FrameStrobe[1] FrameStrobe[2] FrameStrobe[3] FrameStrobe[4] FrameStrobe[5]
+ FrameStrobe[6] FrameStrobe[7] FrameStrobe[8] FrameStrobe[9] FrameStrobe_O[0] FrameStrobe_O[10]
+ FrameStrobe_O[11] FrameStrobe_O[12] FrameStrobe_O[13] FrameStrobe_O[14] FrameStrobe_O[15]
+ FrameStrobe_O[16] FrameStrobe_O[17] FrameStrobe_O[18] FrameStrobe_O[19] FrameStrobe_O[1]
+ FrameStrobe_O[2] FrameStrobe_O[3] FrameStrobe_O[4] FrameStrobe_O[5] FrameStrobe_O[6]
+ FrameStrobe_O[7] FrameStrobe_O[8] FrameStrobe_O[9] N1BEG[0] N1BEG[1] N1BEG[2] N1BEG[3]
+ N2BEG[0] N2BEG[1] N2BEG[2] N2BEG[3] N2BEG[4] N2BEG[5] N2BEG[6] N2BEG[7] N2BEGb[0]
+ N2BEGb[1] N2BEGb[2] N2BEGb[3] N2BEGb[4] N2BEGb[5] N2BEGb[6] N2BEGb[7] N4BEG[0] N4BEG[10]
+ N4BEG[11] N4BEG[12] N4BEG[13] N4BEG[14] N4BEG[15] N4BEG[1] N4BEG[2] N4BEG[3] N4BEG[4]
+ N4BEG[5] N4BEG[6] N4BEG[7] N4BEG[8] N4BEG[9] NN4BEG[0] NN4BEG[10] NN4BEG[11] NN4BEG[12]
+ NN4BEG[13] NN4BEG[14] NN4BEG[15] NN4BEG[1] NN4BEG[2] NN4BEG[3] NN4BEG[4] NN4BEG[5]
+ NN4BEG[6] NN4BEG[7] NN4BEG[8] NN4BEG[9] S1END[0] S1END[1] S1END[2] S1END[3] S2END[0]
+ S2END[1] S2END[2] S2END[3] S2END[4] S2END[5] S2END[6] S2END[7] S2MID[0] S2MID[1]
+ S2MID[2] S2MID[3] S2MID[4] S2MID[5] S2MID[6] S2MID[7] S4END[0] S4END[10] S4END[11]
+ S4END[12] S4END[13] S4END[14] S4END[15] S4END[1] S4END[2] S4END[3] S4END[4] S4END[5]
+ S4END[6] S4END[7] S4END[8] S4END[9] SS4END[0] SS4END[10] SS4END[11] SS4END[12] SS4END[13]
+ SS4END[14] SS4END[15] SS4END[1] SS4END[2] SS4END[3] SS4END[4] SS4END[5] SS4END[6]
+ SS4END[7] SS4END[8] SS4END[9] UserCLK UserCLKo VALUE_top0 VALUE_top1 VALUE_top2
+ VALUE_top3 VALUE_top4 VALUE_top5 VALUE_top6 VALUE_top7 VGND VPWR
XFILLER_10_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_0_Left_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_11_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_062_ net21 net15 VGND VGND VPWR VPWR Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
X_131_ Inst_S_EF_DAC8_switch_matrix.N2BEG2 VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__clkbuf_1
XFILLER_9_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_114_ FrameStrobe[9] VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__clkbuf_1
X_045_ net34 net16 VGND VGND VPWR VPWR Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_5_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_12 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_028_ net19 net13 VGND VGND VPWR VPWR Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XANTENNA_5 FrameStrobe[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput97 net103 VGND VGND VPWR VPWR FrameData_O[28] sky130_fd_sc_hd__buf_2
XFILLER_8_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput86 net92 VGND VGND VPWR VPWR FrameData_O[18] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_2_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_130_ Inst_S_EF_DAC8_switch_matrix.N2BEG1 VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__clkbuf_2
XFILLER_9_23 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_061_ net20 net18 VGND VGND VPWR VPWR Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_4_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_044_ net33 net16 VGND VGND VPWR VPWR Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
X_113_ FrameStrobe[8] VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_5_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_6 FrameStrobe[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_027_ net11 net14 VGND VGND VPWR VPWR Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput98 net104 VGND VGND VPWR VPWR FrameData_O[29] sky130_fd_sc_hd__buf_2
Xoutput87 net93 VGND VGND VPWR VPWR FrameData_O[19] sky130_fd_sc_hd__buf_2
XFILLER_0_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_123 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_060_ net19 net17 VGND VGND VPWR VPWR Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_9_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_5_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_112_ FrameStrobe[7] VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__clkbuf_1
X_043_ net32 net17 VGND VGND VPWR VPWR Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
XANTENNA_7 net136 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_026_ net10 net14 VGND VGND VPWR VPWR Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput99 net105 VGND VGND VPWR VPWR FrameData_O[2] sky130_fd_sc_hd__buf_2
Xoutput88 net94 VGND VGND VPWR VPWR FrameData_O[1] sky130_fd_sc_hd__buf_2
Xoutput77 net83 VGND VGND VPWR VPWR FrameData_O[0] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_2_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_009_ net44 net60 net74 net82 Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit12.Q Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit13.Q
+ VGND VGND VPWR VPWR Inst_S_EF_DAC8_switch_matrix.N2BEGb6 sky130_fd_sc_hd__mux4_1
XFILLER_9_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_11_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_4_Left_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_042_ net29 net17 VGND VGND VPWR VPWR Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
X_111_ FrameStrobe[6] VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__clkbuf_1
XANTENNA_8 net146 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_025_ net9 net14 VGND VGND VPWR VPWR Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_3_252 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput89 net95 VGND VGND VPWR VPWR FrameData_O[20] sky130_fd_sc_hd__buf_2
XFILLER_0_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_2_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput78 net84 VGND VGND VPWR VPWR FrameData_O[10] sky130_fd_sc_hd__buf_2
XFILLER_8_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_008_ net43 net59 net67 net81 Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit14.Q Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit15.Q
+ VGND VGND VPWR VPWR Inst_S_EF_DAC8_switch_matrix.N2BEGb7 sky130_fd_sc_hd__mux4_1
XFILLER_7_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_041_ net12 net15 VGND VGND VPWR VPWR Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_7_228 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_110_ FrameStrobe[5] VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__clkbuf_1
XFILLER_10_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_283 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_9 net155 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_024_ net8 net13 VGND VGND VPWR VPWR Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_3_264 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_007_ net51 net47 net59 net67 Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit16.Q Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit17.Q
+ VGND VGND VPWR VPWR net188 sky130_fd_sc_hd__mux4_2
Xoutput79 net85 VGND VGND VPWR VPWR FrameData_O[11] sky130_fd_sc_hd__buf_2
XFILLER_5_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_040_ net1 net15 VGND VGND VPWR VPWR Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
X_169_ net80 VGND VGND VPWR VPWR net185 sky130_fd_sc_hd__clkbuf_1
XFILLER_6_295 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_023_ net58 net80 net66 net73 Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit17.Q Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit16.Q
+ VGND VGND VPWR VPWR Inst_S_EF_DAC8_switch_matrix.N2BEG0 sky130_fd_sc_hd__mux4_1
XFILLER_3_210 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_006_ net52 net48 net60 net74 Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit18.Q Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit19.Q
+ VGND VGND VPWR VPWR net189 sky130_fd_sc_hd__mux4_1
XFILLER_5_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_168_ net81 VGND VGND VPWR VPWR net184 sky130_fd_sc_hd__buf_1
X_099_ net25 VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__clkbuf_2
XFILLER_1_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_022_ net57 net79 net65 net72 Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit19.Q Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit18.Q
+ VGND VGND VPWR VPWR Inst_S_EF_DAC8_switch_matrix.N2BEG1 sky130_fd_sc_hd__mux4_1
XFILLER_0_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_005_ net53 net49 net61 net75 Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit20.Q Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit21.Q
+ VGND VGND VPWR VPWR net190 sky130_fd_sc_hd__mux4_2
XFILLER_7_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_350 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_098_ net24 VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__clkbuf_2
X_167_ net82 VGND VGND VPWR VPWR net183 sky130_fd_sc_hd__clkbuf_1
X_021_ net56 net78 net64 net71 Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit21.Q Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit20.Q
+ VGND VGND VPWR VPWR Inst_S_EF_DAC8_switch_matrix.N2BEG2 sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_11_Left_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_004_ net54 net50 net62 net76 Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit22.Q Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit23.Q
+ VGND VGND VPWR VPWR net191 sky130_fd_sc_hd__mux4_1
XFILLER_5_307 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_097_ net23 VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__clkbuf_2
XFILLER_1_31 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_166_ net68 VGND VGND VPWR VPWR net182 sky130_fd_sc_hd__buf_1
X_020_ net55 net77 net63 net70 Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit23.Q Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit22.Q
+ VGND VGND VPWR VPWR Inst_S_EF_DAC8_switch_matrix.N2BEG3 sky130_fd_sc_hd__mux4_1
XFILLER_10_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_149_ S4END[11] VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_6_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_003_ net39 net43 net63 net77 Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit24.Q Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit25.Q
+ VGND VGND VPWR VPWR net192 sky130_fd_sc_hd__mux4_1
XFILLER_7_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_319 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_311 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_196 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_165_ net69 VGND VGND VPWR VPWR net181 sky130_fd_sc_hd__clkbuf_1
X_096_ net22 VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__buf_1
XFILLER_1_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_148_ S4END[12] VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_6_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_079_ net35 VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__buf_1
XFILLER_2_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_239 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_002_ net40 net44 net64 net78 Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit26.Q Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit27.Q
+ VGND VGND VPWR VPWR net193 sky130_fd_sc_hd__mux4_1
XFILLER_7_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_323 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_164_ net70 VGND VGND VPWR VPWR net180 sky130_fd_sc_hd__clkbuf_1
X_095_ net21 VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__buf_1
XFILLER_6_212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_6_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_147_ S4END[13] VGND VGND VPWR VPWR net163 sky130_fd_sc_hd__clkbuf_2
X_078_ net34 VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__clkbuf_2
X_001_ net41 net45 net65 net79 Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit28.Q Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit29.Q
+ VGND VGND VPWR VPWR net194 sky130_fd_sc_hd__mux4_2
XFILLER_7_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_3_Left_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_224 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_094_ net20 VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__clkbuf_2
X_163_ net71 VGND VGND VPWR VPWR net179 sky130_fd_sc_hd__buf_1
XFILLER_10_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_146_ S4END[14] VGND VGND VPWR VPWR net162 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_6_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_077_ net33 VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__clkbuf_2
X_000_ net42 net46 net66 net80 Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit30.Q Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit31.Q
+ VGND VGND VPWR VPWR net195 sky130_fd_sc_hd__mux4_1
XFILLER_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_129_ Inst_S_EF_DAC8_switch_matrix.N2BEG0 VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__buf_1
XFILLER_7_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_236 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_093_ net19 VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__buf_1
X_162_ net72 VGND VGND VPWR VPWR net178 sky130_fd_sc_hd__buf_1
Xinput1 FrameData[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__buf_1
X_145_ S4END[15] VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_6_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_076_ net32 VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_128_ net39 VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__buf_1
X_059_ net11 net16 VGND VGND VPWR VPWR Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput70 SS4END[3] VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_3_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_161_ net73 VGND VGND VPWR VPWR net171 sky130_fd_sc_hd__clkbuf_1
XFILLER_6_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_092_ net11 VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__clkbuf_2
XFILLER_5_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput2 FrameData[10] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__buf_1
X_144_ Inst_S_EF_DAC8_switch_matrix.N2BEGb7 VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_6_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_075_ net29 VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__clkbuf_1
Xoutput180 net186 VGND VGND VPWR VPWR NN4BEG[9] sky130_fd_sc_hd__buf_2
XFILLER_7_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_058_ net10 net16 VGND VGND VPWR VPWR Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
X_127_ net40 VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__clkbuf_1
Xinput60 S4END[7] VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__buf_1
Xinput71 SS4END[4] VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_3_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout13 FrameStrobe[1] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__clkbuf_2
XFILLER_10_278 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_160_ net59 VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__buf_1
X_091_ net10 VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_7_Left_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput3 FrameData[11] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__buf_1
XFILLER_10_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_074_ net12 VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__clkbuf_2
X_143_ Inst_S_EF_DAC8_switch_matrix.N2BEGb6 VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__clkbuf_1
Xoutput170 net176 VGND VGND VPWR VPWR NN4BEG[14] sky130_fd_sc_hd__buf_2
Xoutput181 net187 VGND VGND VPWR VPWR UserCLKo sky130_fd_sc_hd__buf_1
XFILLER_11_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_057_ net9 net15 VGND VGND VPWR VPWR Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_7_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_25 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_126_ net41 VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__clkbuf_2
Xinput72 SS4END[5] VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__clkbuf_2
Xinput61 SS4END[0] VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__buf_1
Xinput50 S2MID[5] VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_314 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_109_ FrameStrobe[4] VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__clkbuf_1
XFILLER_3_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout14 FrameStrobe[1] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_9_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_090_ net9 VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__buf_1
XFILLER_5_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput4 FrameData[12] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_1
XFILLER_10_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_142_ Inst_S_EF_DAC8_switch_matrix.N2BEGb5 VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__buf_1
X_073_ net1 VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__clkbuf_2
Xoutput171 net177 VGND VGND VPWR VPWR NN4BEG[15] sky130_fd_sc_hd__buf_2
Xoutput160 net166 VGND VGND VPWR VPWR N4BEG[5] sky130_fd_sc_hd__buf_2
X_125_ net42 VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__buf_1
X_056_ net8 net18 VGND VGND VPWR VPWR Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_7_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput182 net188 VGND VGND VPWR VPWR VALUE_top0 sky130_fd_sc_hd__buf_2
Xinput40 S2END[3] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__buf_1
Xinput51 S2MID[6] VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__clkbuf_1
Xinput73 SS4END[6] VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__buf_1
Xinput62 SS4END[10] VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_10_Left_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_7_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_326 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_039_ net31 net14 VGND VGND VPWR VPWR Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
X_108_ FrameStrobe[3] VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_10_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout15 net18 VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__clkbuf_2
XFILLER_9_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput5 FrameData[13] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_1
XFILLER_10_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_141_ Inst_S_EF_DAC8_switch_matrix.N2BEGb4 VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__clkbuf_1
XANTENNA_10 net162 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput150 net156 VGND VGND VPWR VPWR N4BEG[10] sky130_fd_sc_hd__buf_2
Xoutput172 net178 VGND VGND VPWR VPWR NN4BEG[1] sky130_fd_sc_hd__buf_2
Xoutput161 net167 VGND VGND VPWR VPWR N4BEG[6] sky130_fd_sc_hd__buf_2
X_124_ FrameStrobe[19] VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__clkbuf_1
XFILLER_7_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_055_ net7 net15 VGND VGND VPWR VPWR Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_7_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput183 net189 VGND VGND VPWR VPWR VALUE_top1 sky130_fd_sc_hd__buf_2
Xinput41 S2END[4] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__buf_1
Xinput52 S2MID[7] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__clkbuf_1
Xinput74 SS4END[7] VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__buf_1
Xinput63 SS4END[11] VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_7_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput30 FrameData[7] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__buf_1
XFILLER_4_338 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_038_ net30 net14 VGND VGND VPWR VPWR Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
X_107_ FrameStrobe[2] VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__clkbuf_1
XFILLER_3_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout16 net18 VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_4_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput6 FrameData[14] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__buf_1
X_071_ net31 net17 VGND VGND VPWR VPWR Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
X_140_ Inst_S_EF_DAC8_switch_matrix.N2BEGb3 VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__clkbuf_1
Xoutput173 net179 VGND VGND VPWR VPWR NN4BEG[2] sky130_fd_sc_hd__buf_2
Xoutput162 net168 VGND VGND VPWR VPWR N4BEG[7] sky130_fd_sc_hd__buf_2
XANTENNA_11 net164 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput140 net146 VGND VGND VPWR VPWR N2BEG[7] sky130_fd_sc_hd__buf_2
Xoutput151 net157 VGND VGND VPWR VPWR N4BEG[11] sky130_fd_sc_hd__buf_2
Xoutput184 net190 VGND VGND VPWR VPWR VALUE_top2 sky130_fd_sc_hd__buf_2
Xinput20 FrameData[27] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__buf_1
X_123_ FrameStrobe[18] VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__clkbuf_1
X_054_ net6 net15 VGND VGND VPWR VPWR Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_7_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput31 FrameData[8] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__buf_1
Xinput64 SS4END[12] VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__buf_1
Xinput53 S4END[0] VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__buf_1
Xinput42 S2END[5] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__buf_1
Xinput75 SS4END[8] VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__buf_1
X_037_ net28 net13 VGND VGND VPWR VPWR Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_3_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_106_ net13 VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout17 net18 VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__clkbuf_2
XFILLER_10_216 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput7 FrameData[15] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_1_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_070_ net30 net17 VGND VGND VPWR VPWR Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_2_256 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput174 net180 VGND VGND VPWR VPWR NN4BEG[3] sky130_fd_sc_hd__buf_2
Xoutput152 net158 VGND VGND VPWR VPWR N4BEG[12] sky130_fd_sc_hd__buf_2
Xoutput163 net169 VGND VGND VPWR VPWR N4BEG[8] sky130_fd_sc_hd__buf_2
XANTENNA_12 net165 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput130 net136 VGND VGND VPWR VPWR N1BEG[1] sky130_fd_sc_hd__buf_2
Xoutput141 net147 VGND VGND VPWR VPWR N2BEGb[0] sky130_fd_sc_hd__buf_2
Xoutput185 net191 VGND VGND VPWR VPWR VALUE_top3 sky130_fd_sc_hd__buf_2
X_122_ FrameStrobe[17] VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__clkbuf_1
XFILLER_7_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_053_ net5 net16 VGND VGND VPWR VPWR Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput65 SS4END[13] VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__clkbuf_2
Xinput76 SS4END[9] VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput54 S4END[1] VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput43 S2END[6] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__buf_1
Xinput21 FrameData[28] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__clkbuf_2
Xinput10 FrameData[18] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__buf_1
Xinput32 FrameData[9] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__buf_1
XFILLER_11_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_105_ net17 VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__clkbuf_1
XFILLER_4_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_036_ net27 net13 VGND VGND VPWR VPWR Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_3_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_019_ net54 net62 net76 net69 Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit24.Q Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit25.Q
+ VGND VGND VPWR VPWR Inst_S_EF_DAC8_switch_matrix.N2BEG4 sky130_fd_sc_hd__mux4_1
XFILLER_0_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout18 FrameStrobe[0] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__clkbuf_2
XFILLER_8_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_228 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput8 FrameData[16] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_1_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_2_Left_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput120 net126 VGND VGND VPWR VPWR FrameStrobe_O[1] sky130_fd_sc_hd__buf_2
Xoutput153 net159 VGND VGND VPWR VPWR N4BEG[13] sky130_fd_sc_hd__buf_2
Xoutput142 net148 VGND VGND VPWR VPWR N2BEGb[1] sky130_fd_sc_hd__buf_2
Xoutput131 net137 VGND VGND VPWR VPWR N1BEG[2] sky130_fd_sc_hd__buf_2
Xoutput175 net181 VGND VGND VPWR VPWR NN4BEG[4] sky130_fd_sc_hd__buf_2
Xoutput164 net170 VGND VGND VPWR VPWR N4BEG[9] sky130_fd_sc_hd__buf_2
XANTENNA_13 S4END[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput186 net192 VGND VGND VPWR VPWR VALUE_top4 sky130_fd_sc_hd__buf_2
XFILLER_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_121_ FrameStrobe[16] VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__clkbuf_1
XFILLER_7_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_052_ net4 net16 VGND VGND VPWR VPWR Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput55 S4END[2] VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__buf_1
Xinput44 S2END[7] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__buf_1
Xinput66 SS4END[14] VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__buf_1
Xinput33 S1END[0] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__clkbuf_1
Xinput22 FrameData[29] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__clkbuf_2
Xinput11 FrameData[19] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_7_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_104_ net31 VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__buf_1
XFILLER_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_035_ net26 net14 VGND VGND VPWR VPWR Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_3_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_018_ net53 net61 net75 net68 Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit26.Q Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit27.Q
+ VGND VGND VPWR VPWR Inst_S_EF_DAC8_switch_matrix.N2BEG5 sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_4_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput9 FrameData[17] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_5_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput110 net116 VGND VGND VPWR VPWR FrameStrobe_O[10] sky130_fd_sc_hd__buf_2
Xoutput121 net127 VGND VGND VPWR VPWR FrameStrobe_O[2] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput143 net149 VGND VGND VPWR VPWR N2BEGb[2] sky130_fd_sc_hd__buf_2
Xoutput132 net138 VGND VGND VPWR VPWR N1BEG[3] sky130_fd_sc_hd__buf_2
XANTENNA_14 S4END[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput176 net182 VGND VGND VPWR VPWR NN4BEG[5] sky130_fd_sc_hd__buf_2
Xoutput165 net171 VGND VGND VPWR VPWR NN4BEG[0] sky130_fd_sc_hd__buf_2
Xoutput154 net160 VGND VGND VPWR VPWR N4BEG[14] sky130_fd_sc_hd__buf_2
X_120_ FrameStrobe[15] VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__clkbuf_1
XFILLER_7_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput187 net193 VGND VGND VPWR VPWR VALUE_top5 sky130_fd_sc_hd__buf_2
X_051_ net3 net17 VGND VGND VPWR VPWR Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput45 S2MID[0] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__buf_1
Xinput67 SS4END[15] VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__buf_1
Xinput56 S4END[3] VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__buf_1
Xinput34 S1END[1] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_7_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput12 FrameData[1] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__buf_1
Xinput23 FrameData[2] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_4_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_103_ net30 VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__buf_1
XFILLER_7_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_034_ net25 net14 VGND VGND VPWR VPWR Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_8_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_180 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_017_ net52 net60 net74 net82 Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit28.Q Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit29.Q
+ VGND VGND VPWR VPWR Inst_S_EF_DAC8_switch_matrix.N2BEG6 sky130_fd_sc_hd__mux4_1
XFILLER_8_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_15 net194 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput100 net106 VGND VGND VPWR VPWR FrameData_O[30] sky130_fd_sc_hd__buf_2
Xoutput122 net128 VGND VGND VPWR VPWR FrameStrobe_O[3] sky130_fd_sc_hd__buf_2
Xoutput155 net161 VGND VGND VPWR VPWR N4BEG[15] sky130_fd_sc_hd__buf_2
Xoutput144 net150 VGND VGND VPWR VPWR N2BEGb[3] sky130_fd_sc_hd__buf_2
Xoutput133 net139 VGND VGND VPWR VPWR N2BEG[0] sky130_fd_sc_hd__buf_2
Xoutput111 net117 VGND VGND VPWR VPWR FrameStrobe_O[11] sky130_fd_sc_hd__buf_2
Xoutput166 net172 VGND VGND VPWR VPWR NN4BEG[10] sky130_fd_sc_hd__buf_2
Xoutput177 net183 VGND VGND VPWR VPWR NN4BEG[6] sky130_fd_sc_hd__buf_2
XFILLER_7_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_050_ net2 net17 VGND VGND VPWR VPWR Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput188 net194 VGND VGND VPWR VPWR VALUE_top6 sky130_fd_sc_hd__buf_2
Xinput68 SS4END[1] VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput46 S2MID[1] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__buf_1
Xinput35 S1END[2] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__buf_1
XFILLER_11_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput24 FrameData[30] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_10_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput57 S4END[4] VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__buf_1
Xinput13 FrameData[20] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_7_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_033_ net24 net13 VGND VGND VPWR VPWR Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
X_102_ net28 VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__buf_1
XFILLER_6_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_016_ net51 net59 net67 net81 Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit30.Q Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit31.Q
+ VGND VGND VPWR VPWR Inst_S_EF_DAC8_switch_matrix.N2BEG7 sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_4_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput112 net118 VGND VGND VPWR VPWR FrameStrobe_O[12] sky130_fd_sc_hd__buf_2
Xoutput123 net129 VGND VGND VPWR VPWR FrameStrobe_O[4] sky130_fd_sc_hd__buf_2
Xoutput167 net173 VGND VGND VPWR VPWR NN4BEG[11] sky130_fd_sc_hd__buf_2
Xoutput178 net184 VGND VGND VPWR VPWR NN4BEG[7] sky130_fd_sc_hd__buf_2
Xoutput156 net162 VGND VGND VPWR VPWR N4BEG[1] sky130_fd_sc_hd__buf_2
Xoutput145 net151 VGND VGND VPWR VPWR N2BEGb[4] sky130_fd_sc_hd__buf_2
XANTENNA_16 net144 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput134 net140 VGND VGND VPWR VPWR N2BEG[1] sky130_fd_sc_hd__buf_2
Xoutput101 net107 VGND VGND VPWR VPWR FrameData_O[31] sky130_fd_sc_hd__buf_2
XFILLER_9_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_6_Left_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput189 net195 VGND VGND VPWR VPWR VALUE_top7 sky130_fd_sc_hd__buf_2
Xinput36 S1END[3] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__clkbuf_1
Xinput25 FrameData[31] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput14 FrameData[21] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__buf_1
Xinput58 S4END[5] VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput47 S2MID[2] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__buf_1
Xinput69 SS4END[2] VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__buf_1
XFILLER_6_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_032_ net23 net13 VGND VGND VPWR VPWR Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
X_101_ net27 VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__buf_1
XFILLER_3_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_9_Left_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_015_ net50 net80 net66 net73 Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit1.Q Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit0.Q
+ VGND VGND VPWR VPWR Inst_S_EF_DAC8_switch_matrix.N2BEGb0 sky130_fd_sc_hd__mux4_1
XFILLER_8_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_250 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_12 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput124 net130 VGND VGND VPWR VPWR FrameStrobe_O[5] sky130_fd_sc_hd__buf_2
Xoutput168 net174 VGND VGND VPWR VPWR NN4BEG[12] sky130_fd_sc_hd__buf_2
Xoutput179 net185 VGND VGND VPWR VPWR NN4BEG[8] sky130_fd_sc_hd__buf_2
Xoutput146 net152 VGND VGND VPWR VPWR N2BEGb[5] sky130_fd_sc_hd__buf_2
Xoutput113 net119 VGND VGND VPWR VPWR FrameStrobe_O[13] sky130_fd_sc_hd__buf_2
Xoutput157 net163 VGND VGND VPWR VPWR N4BEG[2] sky130_fd_sc_hd__buf_2
Xoutput135 net141 VGND VGND VPWR VPWR N2BEG[2] sky130_fd_sc_hd__buf_2
Xoutput102 net108 VGND VGND VPWR VPWR FrameData_O[3] sky130_fd_sc_hd__buf_2
XANTENNA_17 net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput37 S2END[0] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__buf_1
Xinput48 S2MID[3] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__buf_1
Xinput59 S4END[6] VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__buf_1
Xinput15 FrameData[22] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__buf_1
XFILLER_6_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput26 FrameData[3] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__dlymetal6s2s_1
X_177_ UserCLK VGND VGND VPWR VPWR net187 sky130_fd_sc_hd__buf_2
XFILLER_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_031_ net22 net13 VGND VGND VPWR VPWR Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
X_100_ net26 VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__clkbuf_2
XFILLER_8_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_014_ net49 net79 net65 net72 Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit3.Q Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit2.Q
+ VGND VGND VPWR VPWR Inst_S_EF_DAC8_switch_matrix.N2BEGb1 sky130_fd_sc_hd__mux4_1
XFILLER_5_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput114 net120 VGND VGND VPWR VPWR FrameStrobe_O[14] sky130_fd_sc_hd__buf_2
Xoutput125 net131 VGND VGND VPWR VPWR FrameStrobe_O[6] sky130_fd_sc_hd__buf_2
Xoutput169 net175 VGND VGND VPWR VPWR NN4BEG[13] sky130_fd_sc_hd__buf_2
Xoutput158 net164 VGND VGND VPWR VPWR N4BEG[3] sky130_fd_sc_hd__buf_2
Xoutput136 net142 VGND VGND VPWR VPWR N2BEG[3] sky130_fd_sc_hd__buf_2
Xoutput147 net153 VGND VGND VPWR VPWR N2BEGb[6] sky130_fd_sc_hd__buf_2
XFILLER_9_362 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_262 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput103 net109 VGND VGND VPWR VPWR FrameData_O[4] sky130_fd_sc_hd__buf_2
XFILLER_2_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_18 net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput38 S2END[1] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__buf_1
Xinput49 S2MID[4] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__clkbuf_1
X_176_ net67 VGND VGND VPWR VPWR net177 sky130_fd_sc_hd__clkbuf_1
Xinput16 FrameData[23] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__buf_1
XFILLER_6_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput27 FrameData[4] VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__clkbuf_1
XFILLER_9_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_030_ net21 net13 VGND VGND VPWR VPWR Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
X_159_ net60 VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_013_ net48 net78 net64 net71 Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit5.Q Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit4.Q
+ VGND VGND VPWR VPWR Inst_S_EF_DAC8_switch_matrix.N2BEGb2 sky130_fd_sc_hd__mux4_1
XFILLER_3_198 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput159 net165 VGND VGND VPWR VPWR N4BEG[4] sky130_fd_sc_hd__buf_2
Xoutput148 net154 VGND VGND VPWR VPWR N2BEGb[7] sky130_fd_sc_hd__buf_2
Xoutput137 net143 VGND VGND VPWR VPWR N2BEG[4] sky130_fd_sc_hd__buf_2
Xoutput115 net121 VGND VGND VPWR VPWR FrameStrobe_O[15] sky130_fd_sc_hd__buf_2
Xoutput126 net132 VGND VGND VPWR VPWR FrameStrobe_O[7] sky130_fd_sc_hd__buf_2
XFILLER_9_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput104 net110 VGND VGND VPWR VPWR FrameData_O[5] sky130_fd_sc_hd__buf_2
XANTENNA_19 net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput39 S2END[2] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__buf_1
XFILLER_10_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput17 FrameData[24] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__buf_1
XFILLER_6_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput28 FrameData[5] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__clkbuf_1
X_175_ net74 VGND VGND VPWR VPWR net176 sky130_fd_sc_hd__clkbuf_1
XFILLER_3_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_089_ net8 VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__buf_1
X_158_ net61 VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__buf_1
X_012_ net47 net77 net63 net70 Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit7.Q Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit6.Q
+ VGND VGND VPWR VPWR Inst_S_EF_DAC8_switch_matrix.N2BEGb3 sky130_fd_sc_hd__mux4_1
XFILLER_3_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput116 net122 VGND VGND VPWR VPWR FrameStrobe_O[16] sky130_fd_sc_hd__buf_2
Xoutput127 net133 VGND VGND VPWR VPWR FrameStrobe_O[8] sky130_fd_sc_hd__buf_2
Xoutput138 net144 VGND VGND VPWR VPWR N2BEG[5] sky130_fd_sc_hd__buf_2
XFILLER_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput149 net155 VGND VGND VPWR VPWR N4BEG[0] sky130_fd_sc_hd__buf_2
Xoutput105 net111 VGND VGND VPWR VPWR FrameData_O[6] sky130_fd_sc_hd__buf_2
XFILLER_10_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput18 FrameData[25] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__buf_1
XFILLER_6_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput29 FrameData[6] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__buf_1
X_174_ net75 VGND VGND VPWR VPWR net175 sky130_fd_sc_hd__clkbuf_1
XFILLER_3_80 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_157_ net62 VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__clkbuf_1
X_088_ net7 VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_8_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_011_ net46 net62 net76 net69 Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit8.Q Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit9.Q
+ VGND VGND VPWR VPWR Inst_S_EF_DAC8_switch_matrix.N2BEGb4 sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_4_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput117 net123 VGND VGND VPWR VPWR FrameStrobe_O[17] sky130_fd_sc_hd__buf_2
Xoutput128 net134 VGND VGND VPWR VPWR FrameStrobe_O[9] sky130_fd_sc_hd__buf_2
Xoutput139 net145 VGND VGND VPWR VPWR N2BEG[6] sky130_fd_sc_hd__buf_2
Xoutput106 net112 VGND VGND VPWR VPWR FrameData_O[7] sky130_fd_sc_hd__buf_2
Xinput19 FrameData[26] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__buf_1
X_173_ net76 VGND VGND VPWR VPWR net174 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_1_Left_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_156_ net63 VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__clkbuf_1
X_087_ net6 VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__buf_1
XFILLER_8_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XS_EF_DAC8_190 VGND VGND VPWR VPWR S_EF_DAC8_190/HI Co sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_8_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_010_ net45 net61 net75 net68 Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit10.Q Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit11.Q
+ VGND VGND VPWR VPWR Inst_S_EF_DAC8_switch_matrix.N2BEGb5 sky130_fd_sc_hd__mux4_1
X_139_ Inst_S_EF_DAC8_switch_matrix.N2BEGb2 VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_5_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput118 net124 VGND VGND VPWR VPWR FrameStrobe_O[18] sky130_fd_sc_hd__buf_2
Xoutput129 net135 VGND VGND VPWR VPWR N1BEG[0] sky130_fd_sc_hd__buf_2
Xoutput107 net113 VGND VGND VPWR VPWR FrameData_O[8] sky130_fd_sc_hd__buf_2
XFILLER_10_343 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_172_ net77 VGND VGND VPWR VPWR net173 sky130_fd_sc_hd__clkbuf_1
XFILLER_5_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_144 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_086_ net5 VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__clkbuf_2
X_155_ net64 VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_8_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_069_ net28 net17 VGND VGND VPWR VPWR Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
X_138_ Inst_S_EF_DAC8_switch_matrix.N2BEGb1 VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__buf_1
XFILLER_0_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput119 net125 VGND VGND VPWR VPWR FrameStrobe_O[19] sky130_fd_sc_hd__buf_2
Xoutput90 net96 VGND VGND VPWR VPWR FrameData_O[21] sky130_fd_sc_hd__buf_2
XFILLER_9_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_2_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput108 net114 VGND VGND VPWR VPWR FrameData_O[9] sky130_fd_sc_hd__buf_2
XFILLER_10_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_171_ net78 VGND VGND VPWR VPWR net172 sky130_fd_sc_hd__buf_1
XFILLER_10_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_8_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_085_ net4 VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__clkbuf_2
X_154_ net65 VGND VGND VPWR VPWR net170 sky130_fd_sc_hd__buf_1
XFILLER_2_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_137_ Inst_S_EF_DAC8_switch_matrix.N2BEGb0 VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__buf_1
X_068_ net27 net17 VGND VGND VPWR VPWR Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_2_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput109 net115 VGND VGND VPWR VPWR FrameStrobe_O[0] sky130_fd_sc_hd__buf_2
XFILLER_9_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput91 net97 VGND VGND VPWR VPWR FrameData_O[22] sky130_fd_sc_hd__buf_2
Xoutput80 net86 VGND VGND VPWR VPWR FrameData_O[12] sky130_fd_sc_hd__buf_2
X_170_ net79 VGND VGND VPWR VPWR net186 sky130_fd_sc_hd__buf_1
XFILLER_5_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_5_Left_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_153_ net66 VGND VGND VPWR VPWR net169 sky130_fd_sc_hd__clkbuf_1
XFILLER_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_168 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_084_ net3 VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__buf_1
XFILLER_2_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_136_ Inst_S_EF_DAC8_switch_matrix.N2BEG7 VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__clkbuf_1
XFILLER_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_067_ net26 net16 VGND VGND VPWR VPWR Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_8_Left_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_119_ FrameStrobe[14] VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__clkbuf_1
XFILLER_7_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput92 net98 VGND VGND VPWR VPWR FrameData_O[23] sky130_fd_sc_hd__buf_2
Xoutput81 net87 VGND VGND VPWR VPWR FrameData_O[13] sky130_fd_sc_hd__buf_2
XFILLER_10_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_9_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_152_ S4END[8] VGND VGND VPWR VPWR net168 sky130_fd_sc_hd__buf_1
X_083_ net2 VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__buf_1
X_135_ Inst_S_EF_DAC8_switch_matrix.N2BEG6 VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__clkbuf_1
X_066_ net25 net16 VGND VGND VPWR VPWR Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
X_118_ FrameStrobe[13] VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__clkbuf_1
X_049_ net38 net16 VGND VGND VPWR VPWR Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_4_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_1 net110 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput93 net99 VGND VGND VPWR VPWR FrameData_O[24] sky130_fd_sc_hd__buf_2
XFILLER_9_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput82 net88 VGND VGND VPWR VPWR FrameData_O[14] sky130_fd_sc_hd__buf_2
XFILLER_10_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_166 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_151_ S4END[9] VGND VGND VPWR VPWR net167 sky130_fd_sc_hd__buf_1
X_082_ net38 VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__clkbuf_2
XFILLER_2_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_065_ net24 net18 VGND VGND VPWR VPWR Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_134_ Inst_S_EF_DAC8_switch_matrix.N2BEG5 VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__buf_1
X_117_ FrameStrobe[12] VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__clkbuf_1
X_048_ net37 net16 VGND VGND VPWR VPWR Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_6_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_2 FrameStrobe[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput94 net100 VGND VGND VPWR VPWR FrameData_O[25] sky130_fd_sc_hd__buf_2
XFILLER_9_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput83 net89 VGND VGND VPWR VPWR FrameData_O[15] sky130_fd_sc_hd__buf_2
XFILLER_0_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_150_ S4END[10] VGND VGND VPWR VPWR net166 sky130_fd_sc_hd__clkbuf_2
X_081_ net37 VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__clkbuf_2
XFILLER_5_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_064_ net23 net15 VGND VGND VPWR VPWR Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
X_133_ Inst_S_EF_DAC8_switch_matrix.N2BEG4 VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__clkbuf_1
X_116_ FrameStrobe[11] VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__clkbuf_1
X_047_ net36 net15 VGND VGND VPWR VPWR Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_3 FrameStrobe[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput95 net101 VGND VGND VPWR VPWR FrameData_O[26] sky130_fd_sc_hd__buf_2
Xoutput84 net90 VGND VGND VPWR VPWR FrameData_O[16] sky130_fd_sc_hd__buf_2
XFILLER_6_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_080_ net36 VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_8_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_323 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_132_ Inst_S_EF_DAC8_switch_matrix.N2BEG3 VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__clkbuf_1
X_063_ net22 net15 VGND VGND VPWR VPWR Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_2_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_046_ net35 net15 VGND VGND VPWR VPWR Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
X_115_ FrameStrobe[10] VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_5_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_4 FrameStrobe[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_029_ net20 net13 VGND VGND VPWR VPWR Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_3_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_2_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput96 net102 VGND VGND VPWR VPWR FrameData_O[27] sky130_fd_sc_hd__buf_2
Xoutput85 net91 VGND VGND VPWR VPWR FrameData_O[17] sky130_fd_sc_hd__buf_2
XFILLER_0_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
.ends

