* NGSPICE file created from S_CPU_IRQ.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlxtp_1 abstract view
.subckt sky130_fd_sc_hd__dlxtp_1 D GATE VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

.subckt S_CPU_IRQ Co FrameData[0] FrameData[10] FrameData[11] FrameData[12] FrameData[13]
+ FrameData[14] FrameData[15] FrameData[16] FrameData[17] FrameData[18] FrameData[19]
+ FrameData[1] FrameData[20] FrameData[21] FrameData[22] FrameData[23] FrameData[24]
+ FrameData[25] FrameData[26] FrameData[27] FrameData[28] FrameData[29] FrameData[2]
+ FrameData[30] FrameData[31] FrameData[3] FrameData[4] FrameData[5] FrameData[6]
+ FrameData[7] FrameData[8] FrameData[9] FrameData_O[0] FrameData_O[10] FrameData_O[11]
+ FrameData_O[12] FrameData_O[13] FrameData_O[14] FrameData_O[15] FrameData_O[16]
+ FrameData_O[17] FrameData_O[18] FrameData_O[19] FrameData_O[1] FrameData_O[20] FrameData_O[21]
+ FrameData_O[22] FrameData_O[23] FrameData_O[24] FrameData_O[25] FrameData_O[26]
+ FrameData_O[27] FrameData_O[28] FrameData_O[29] FrameData_O[2] FrameData_O[30] FrameData_O[31]
+ FrameData_O[3] FrameData_O[4] FrameData_O[5] FrameData_O[6] FrameData_O[7] FrameData_O[8]
+ FrameData_O[9] FrameStrobe[0] FrameStrobe[10] FrameStrobe[11] FrameStrobe[12] FrameStrobe[13]
+ FrameStrobe[14] FrameStrobe[15] FrameStrobe[16] FrameStrobe[17] FrameStrobe[18]
+ FrameStrobe[19] FrameStrobe[1] FrameStrobe[2] FrameStrobe[3] FrameStrobe[4] FrameStrobe[5]
+ FrameStrobe[6] FrameStrobe[7] FrameStrobe[8] FrameStrobe[9] FrameStrobe_O[0] FrameStrobe_O[10]
+ FrameStrobe_O[11] FrameStrobe_O[12] FrameStrobe_O[13] FrameStrobe_O[14] FrameStrobe_O[15]
+ FrameStrobe_O[16] FrameStrobe_O[17] FrameStrobe_O[18] FrameStrobe_O[19] FrameStrobe_O[1]
+ FrameStrobe_O[2] FrameStrobe_O[3] FrameStrobe_O[4] FrameStrobe_O[5] FrameStrobe_O[6]
+ FrameStrobe_O[7] FrameStrobe_O[8] FrameStrobe_O[9] IRQ_top0 IRQ_top1 IRQ_top2 IRQ_top3
+ N1BEG[0] N1BEG[1] N1BEG[2] N1BEG[3] N2BEG[0] N2BEG[1] N2BEG[2] N2BEG[3] N2BEG[4]
+ N2BEG[5] N2BEG[6] N2BEG[7] N2BEGb[0] N2BEGb[1] N2BEGb[2] N2BEGb[3] N2BEGb[4] N2BEGb[5]
+ N2BEGb[6] N2BEGb[7] N4BEG[0] N4BEG[10] N4BEG[11] N4BEG[12] N4BEG[13] N4BEG[14] N4BEG[15]
+ N4BEG[1] N4BEG[2] N4BEG[3] N4BEG[4] N4BEG[5] N4BEG[6] N4BEG[7] N4BEG[8] N4BEG[9]
+ NN4BEG[0] NN4BEG[10] NN4BEG[11] NN4BEG[12] NN4BEG[13] NN4BEG[14] NN4BEG[15] NN4BEG[1]
+ NN4BEG[2] NN4BEG[3] NN4BEG[4] NN4BEG[5] NN4BEG[6] NN4BEG[7] NN4BEG[8] NN4BEG[9]
+ S1END[0] S1END[1] S1END[2] S1END[3] S2END[0] S2END[1] S2END[2] S2END[3] S2END[4]
+ S2END[5] S2END[6] S2END[7] S2MID[0] S2MID[1] S2MID[2] S2MID[3] S2MID[4] S2MID[5]
+ S2MID[6] S2MID[7] S4END[0] S4END[10] S4END[11] S4END[12] S4END[13] S4END[14] S4END[15]
+ S4END[1] S4END[2] S4END[3] S4END[4] S4END[5] S4END[6] S4END[7] S4END[8] S4END[9]
+ SS4END[0] SS4END[10] SS4END[11] SS4END[12] SS4END[13] SS4END[14] SS4END[15] SS4END[1]
+ SS4END[2] SS4END[3] SS4END[4] SS4END[5] SS4END[6] SS4END[7] SS4END[8] SS4END[9]
+ UserCLK UserCLKo VGND VPWR
XFILLER_10_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_376 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_0_Left_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_131_ net24 VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__clkbuf_1
X_062_ net12 net14 VGND VGND VPWR VPWR Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_045_ _002_ _014_ _018_ VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__o21a_1
X_114_ FrameStrobe[17] VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_5_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_227 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_5 FrameData[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_028_ net34 net38 net42 net46 Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit29.Q Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit30.Q
+ VGND VGND VPWR VPWR _004_ sky130_fd_sc_hd__mux4_1
XFILLER_3_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput86 net87 VGND VGND VPWR VPWR FrameStrobe_O[17] sky130_fd_sc_hd__buf_2
Xoutput97 net98 VGND VGND VPWR VPWR FrameStrobe_O[9] sky130_fd_sc_hd__buf_2
Xoutput64 net65 VGND VGND VPWR VPWR FrameData_O[26] sky130_fd_sc_hd__buf_2
Xoutput53 net54 VGND VGND VPWR VPWR FrameData_O[16] sky130_fd_sc_hd__buf_2
Xoutput75 net76 VGND VGND VPWR VPWR FrameData_O[7] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_2_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_130_ net25 VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__buf_1
XFILLER_9_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_061_ net11 net3 VGND VGND VPWR VPWR Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_2_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_044_ _015_ _016_ _017_ Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit24.Q Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit25.Q
+ VGND VGND VPWR VPWR _018_ sky130_fd_sc_hd__a221o_1
X_113_ FrameStrobe[16] VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_5_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_239 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_027_ Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit22.Q VGND VGND VPWR VPWR _003_ sky130_fd_sc_hd__inv_2
XANTENNA_6 FrameData[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput87 net88 VGND VGND VPWR VPWR FrameStrobe_O[18] sky130_fd_sc_hd__buf_2
Xoutput65 net66 VGND VGND VPWR VPWR FrameData_O[27] sky130_fd_sc_hd__buf_2
Xoutput54 net55 VGND VGND VPWR VPWR FrameData_O[17] sky130_fd_sc_hd__buf_2
XFILLER_0_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput98 net99 VGND VGND VPWR VPWR IRQ_top0 sky130_fd_sc_hd__buf_2
Xoutput76 net77 VGND VGND VPWR VPWR FrameData_O[8] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_2_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_060_ net10 net3 VGND VGND VPWR VPWR Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_112_ FrameStrobe[15] VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__clkbuf_1
X_043_ net20 net24 Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit23.Q VGND VGND VPWR VPWR
+ _017_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_5_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_026_ Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit25.Q VGND VGND VPWR VPWR _002_ sky130_fd_sc_hd__inv_2
XANTENNA_7 FrameData[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput88 net89 VGND VGND VPWR VPWR FrameStrobe_O[19] sky130_fd_sc_hd__buf_2
Xoutput55 net56 VGND VGND VPWR VPWR FrameData_O[18] sky130_fd_sc_hd__buf_2
Xoutput66 net67 VGND VGND VPWR VPWR FrameData_O[28] sky130_fd_sc_hd__buf_2
XFILLER_0_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput99 net100 VGND VGND VPWR VPWR IRQ_top1 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_2_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput77 net78 VGND VGND VPWR VPWR FrameData_O[9] sky130_fd_sc_hd__buf_2
XFILLER_8_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_11_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_4_Left_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_111_ FrameStrobe[14] VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__clkbuf_1
X_042_ net16 Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit23.Q Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit24.Q
+ VGND VGND VPWR VPWR _016_ sky130_fd_sc_hd__o21ba_1
XFILLER_6_271 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_8 net63 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_025_ Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit28.Q VGND VGND VPWR VPWR _001_ sky130_fd_sc_hd__inv_2
Xoutput89 net90 VGND VGND VPWR VPWR FrameStrobe_O[1] sky130_fd_sc_hd__buf_2
Xoutput78 net79 VGND VGND VPWR VPWR FrameStrobe_O[0] sky130_fd_sc_hd__buf_2
Xoutput67 net68 VGND VGND VPWR VPWR FrameData_O[29] sky130_fd_sc_hd__buf_2
Xoutput56 net57 VGND VGND VPWR VPWR FrameData_O[19] sky130_fd_sc_hd__buf_2
XFILLER_0_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_110_ FrameStrobe[13] VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__clkbuf_1
X_041_ net28 Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit23.Q VGND VGND VPWR VPWR _015_
+ sky130_fd_sc_hd__nand2b_1
XFILLER_6_283 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_024_ Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit31.Q VGND VGND VPWR VPWR _000_ sky130_fd_sc_hd__inv_2
XANTENNA_9 FrameStrobe[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput57 net58 VGND VGND VPWR VPWR FrameData_O[1] sky130_fd_sc_hd__buf_2
Xoutput46 net47 VGND VGND VPWR VPWR FrameData_O[0] sky130_fd_sc_hd__buf_2
Xoutput79 net80 VGND VGND VPWR VPWR FrameStrobe_O[10] sky130_fd_sc_hd__buf_2
XFILLER_8_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput68 net69 VGND VGND VPWR VPWR FrameData_O[2] sky130_fd_sc_hd__buf_2
XFILLER_8_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_11_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_040_ net32 net36 net40 net44 Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit23.Q Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit24.Q
+ VGND VGND VPWR VPWR _014_ sky130_fd_sc_hd__mux4_1
XFILLER_6_295 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_169_ UserCLK VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__buf_2
XFILLER_10_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput58 net59 VGND VGND VPWR VPWR FrameData_O[20] sky130_fd_sc_hd__buf_2
Xoutput69 net70 VGND VGND VPWR VPWR FrameData_O[30] sky130_fd_sc_hd__buf_2
XFILLER_8_346 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput47 net48 VGND VGND VPWR VPWR FrameData_O[10] sky130_fd_sc_hd__buf_2
XFILLER_7_71 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_11_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_168_ net39 VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__clkbuf_1
X_099_ FrameStrobe[2] VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__clkbuf_1
XFILLER_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_255 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput59 net60 VGND VGND VPWR VPWR FrameData_O[21] sky130_fd_sc_hd__buf_2
XFILLER_0_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput48 net49 VGND VGND VPWR VPWR FrameData_O[11] sky130_fd_sc_hd__buf_2
XFILLER_8_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_11_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_9_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_167_ net40 VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__buf_1
X_098_ FrameStrobe[1] VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__clkbuf_1
XFILLER_10_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_11_Left_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput49 net50 VGND VGND VPWR VPWR FrameData_O[12] sky130_fd_sc_hd__buf_2
XFILLER_8_315 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_9_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_251 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_097_ net14 VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__buf_1
X_166_ net41 VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__clkbuf_1
XFILLER_3_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_149_ net34 VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_6_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_371 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_263 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_207 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_165_ net42 VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__clkbuf_1
XFILLER_6_222 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_096_ net13 VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__buf_1
XFILLER_10_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_148_ net35 VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_6_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_079_ FrameData[14] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__clkbuf_1
XFILLER_8_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_172 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_9_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_095_ net12 VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__buf_1
XFILLER_6_234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_164_ net43 VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__clkbuf_1
XFILLER_10_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_6_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_078_ FrameData[13] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__clkbuf_2
X_147_ net36 VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__clkbuf_1
XFILLER_8_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XS_CPU_IRQ_155 VGND VGND VPWR VPWR S_CPU_IRQ_155/HI Co sky130_fd_sc_hd__conb_1
XPHY_EDGE_ROW_3_Left_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_163_ net44 VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__buf_1
X_094_ net11 VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__clkbuf_2
X_146_ net37 VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__clkbuf_1
X_077_ FrameData[12] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_6_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_129_ net26 VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_3_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_093_ net10 VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__buf_1
X_162_ net45 VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__clkbuf_1
XFILLER_1_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput1 FrameData[20] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_6_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_076_ FrameData[11] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__clkbuf_2
X_145_ net38 VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__buf_1
XFILLER_0_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_059_ net9 net3 VGND VGND VPWR VPWR Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
X_128_ net27 VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_3_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_161_ net46 VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__clkbuf_1
XFILLER_6_259 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_092_ net9 VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__buf_1
XFILLER_10_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput2 FrameData[21] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__buf_1
XFILLER_5_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_144_ S4END[8] VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_6_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_075_ FrameData[10] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__clkbuf_2
XFILLER_2_90 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_058_ net8 net3 VGND VGND VPWR VPWR Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
X_127_ net28 VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__clkbuf_1
XFILLER_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_3_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_160_ SS4END[8] VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__buf_1
XFILLER_6_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_091_ net8 VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__buf_1
Xinput3 FrameData[22] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_7_Left_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_143_ S4END[9] VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__buf_1
X_074_ FrameData[9] VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__clkbuf_2
XFILLER_11_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_057_ net7 net3 VGND VGND VPWR VPWR Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
X_126_ net29 VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__buf_1
XFILLER_8_119 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_109_ FrameStrobe[12] VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__clkbuf_1
XFILLER_7_130 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_144 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_090_ net7 VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput4 FrameData[23] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__buf_1
XFILLER_5_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_142_ S4END[10] VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__buf_1
XFILLER_2_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_073_ FrameData[8] VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__clkbuf_2
X_125_ net30 VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__buf_1
X_056_ net6 net3 VGND VGND VPWR VPWR Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_7_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput40 SS4END[2] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_10_Left_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_7_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_108_ FrameStrobe[11] VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__clkbuf_1
XFILLER_7_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_039_ _001_ _009_ _013_ VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__o21a_1
XFILLER_7_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput5 FrameData[24] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__buf_1
XFILLER_1_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_141_ S4END[11] VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__buf_1
XFILLER_2_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_276 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_072_ FrameData[7] VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__clkbuf_2
XANTENNA_10 FrameStrobe[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput150 net151 VGND VGND VPWR VPWR NN4BEG[6] sky130_fd_sc_hd__buf_2
X_055_ net5 net3 VGND VGND VPWR VPWR Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
X_124_ S2MID[4] VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__clkbuf_1
XFILLER_7_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput30 S4END[0] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__buf_1
Xinput41 SS4END[3] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__buf_1
XFILLER_6_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_7_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_038_ _010_ _011_ _012_ Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit27.Q Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit28.Q
+ VGND VGND VPWR VPWR _013_ sky130_fd_sc_hd__a221o_1
X_107_ FrameStrobe[10] VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__clkbuf_1
XFILLER_3_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_190 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput6 FrameData[25] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_1
X_140_ S4END[12] VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__buf_1
XFILLER_2_288 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_071_ FrameData[6] VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__clkbuf_2
XFILLER_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput140 net141 VGND VGND VPWR VPWR NN4BEG[11] sky130_fd_sc_hd__buf_2
Xoutput151 net152 VGND VGND VPWR VPWR NN4BEG[7] sky130_fd_sc_hd__buf_2
XANTENNA_11 FrameStrobe[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput31 S4END[1] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__buf_1
Xinput20 S2END[2] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__buf_1
X_123_ S2MID[5] VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__clkbuf_1
X_054_ net4 net3 VGND VGND VPWR VPWR Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_7_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput42 SS4END[4] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__buf_1
XFILLER_4_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_106_ FrameStrobe[9] VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__clkbuf_1
X_037_ net21 net25 Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit26.Q VGND VGND VPWR VPWR
+ _012_ sky130_fd_sc_hd__mux2_1
XFILLER_3_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_239 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput7 FrameData[26] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_1_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_070_ FrameData[5] VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__clkbuf_2
XFILLER_4_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput141 net142 VGND VGND VPWR VPWR NN4BEG[12] sky130_fd_sc_hd__buf_2
Xoutput152 net153 VGND VGND VPWR VPWR NN4BEG[8] sky130_fd_sc_hd__buf_2
Xoutput130 net131 VGND VGND VPWR VPWR N4BEG[2] sky130_fd_sc_hd__buf_2
XANTENNA_12 FrameStrobe[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_322 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_053_ net2 net3 VGND VGND VPWR VPWR Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
X_122_ S2MID[6] VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__clkbuf_1
XFILLER_7_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput43 SS4END[5] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput32 S4END[2] VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__buf_1
Xinput21 S2END[3] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__clkbuf_1
Xinput10 FrameData[29] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__buf_1
XFILLER_6_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_105_ FrameStrobe[8] VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__clkbuf_1
XFILLER_4_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_036_ net17 Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit26.Q Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit27.Q
+ VGND VGND VPWR VPWR _011_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_10_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput8 FrameData[27] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_1_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_2_Left_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput153 net154 VGND VGND VPWR VPWR NN4BEG[9] sky130_fd_sc_hd__buf_2
Xoutput142 net143 VGND VGND VPWR VPWR NN4BEG[13] sky130_fd_sc_hd__buf_2
Xoutput131 net132 VGND VGND VPWR VPWR N4BEG[3] sky130_fd_sc_hd__buf_2
Xoutput120 net121 VGND VGND VPWR VPWR N2BEGb[6] sky130_fd_sc_hd__buf_2
XANTENNA_13 net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_052_ net1 net3 VGND VGND VPWR VPWR Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
X_121_ S2MID[7] VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__clkbuf_1
XFILLER_7_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput33 S4END[3] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__clkbuf_1
Xinput22 S2END[4] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__buf_1
Xinput11 FrameData[30] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__buf_1
Xinput44 SS4END[6] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_7_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_035_ net29 Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit26.Q VGND VGND VPWR VPWR _010_
+ sky130_fd_sc_hd__nand2b_1
X_104_ FrameStrobe[7] VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__clkbuf_1
XFILLER_3_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_4_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput9 FrameData[28] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_1_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput143 net144 VGND VGND VPWR VPWR NN4BEG[14] sky130_fd_sc_hd__buf_2
Xoutput132 net133 VGND VGND VPWR VPWR N4BEG[4] sky130_fd_sc_hd__buf_2
Xoutput121 net122 VGND VGND VPWR VPWR N2BEGb[7] sky130_fd_sc_hd__buf_2
Xoutput110 net111 VGND VGND VPWR VPWR N2BEG[4] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_14 S2MID[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput154 net155 VGND VGND VPWR VPWR UserCLKo sky130_fd_sc_hd__buf_1
X_051_ _003_ _019_ _023_ VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__o21a_1
XFILLER_7_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_120_ net15 VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__buf_1
Xinput45 SS4END[7] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__buf_1
Xinput34 S4END[4] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__buf_1
Xinput23 S2END[5] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__buf_1
Xinput12 FrameData[31] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_7_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_103_ FrameStrobe[6] VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__clkbuf_1
X_034_ net33 net37 net41 net45 Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit26.Q Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit27.Q
+ VGND VGND VPWR VPWR _009_ sky130_fd_sc_hd__mux4_1
XFILLER_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_264 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_15 FrameStrobe[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput144 net145 VGND VGND VPWR VPWR NN4BEG[15] sky130_fd_sc_hd__buf_2
Xoutput133 net134 VGND VGND VPWR VPWR N4BEG[5] sky130_fd_sc_hd__buf_2
Xoutput111 net112 VGND VGND VPWR VPWR N2BEG[5] sky130_fd_sc_hd__buf_2
Xoutput122 net123 VGND VGND VPWR VPWR N4BEG[0] sky130_fd_sc_hd__buf_2
XFILLER_7_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput100 net101 VGND VGND VPWR VPWR IRQ_top2 sky130_fd_sc_hd__buf_2
X_050_ _020_ _021_ _022_ Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit21.Q Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit22.Q
+ VGND VGND VPWR VPWR _023_ sky130_fd_sc_hd__a221o_1
Xinput35 S4END[5] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__buf_1
Xinput24 S2END[6] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__buf_1
XFILLER_11_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_7_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_351 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput13 FrameStrobe[0] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_2_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_102_ FrameStrobe[5] VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__clkbuf_1
X_033_ _000_ _004_ _008_ VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__o21a_1
XFILLER_6_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_16 net148 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput123 net124 VGND VGND VPWR VPWR N4BEG[10] sky130_fd_sc_hd__buf_2
Xoutput145 net146 VGND VGND VPWR VPWR NN4BEG[1] sky130_fd_sc_hd__buf_2
Xoutput134 net135 VGND VGND VPWR VPWR N4BEG[6] sky130_fd_sc_hd__buf_2
Xoutput112 net113 VGND VGND VPWR VPWR N2BEG[6] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_6_Left_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput101 net102 VGND VGND VPWR VPWR IRQ_top3 sky130_fd_sc_hd__buf_2
Xinput36 S4END[6] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__buf_1
Xinput25 S2END[7] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__buf_1
Xinput14 S1END[0] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__buf_1
XFILLER_6_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_101_ FrameStrobe[4] VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__clkbuf_1
X_032_ _005_ _006_ _007_ Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit30.Q Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit31.Q
+ VGND VGND VPWR VPWR _008_ sky130_fd_sc_hd__a221o_1
XFILLER_3_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_98 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_32 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_9_Left_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput146 net147 VGND VGND VPWR VPWR NN4BEG[2] sky130_fd_sc_hd__buf_2
Xoutput135 net136 VGND VGND VPWR VPWR N4BEG[7] sky130_fd_sc_hd__buf_2
Xoutput113 net114 VGND VGND VPWR VPWR N2BEG[7] sky130_fd_sc_hd__buf_2
Xoutput124 net125 VGND VGND VPWR VPWR N4BEG[11] sky130_fd_sc_hd__buf_2
Xoutput102 net103 VGND VGND VPWR VPWR N1BEG[0] sky130_fd_sc_hd__buf_2
Xinput37 S4END[7] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__buf_1
Xinput26 S2MID[0] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__clkbuf_1
XFILLER_10_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput15 S1END[1] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__buf_1
XFILLER_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_031_ net22 net26 Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit29.Q VGND VGND VPWR VPWR
+ _007_ sky130_fd_sc_hd__mux2_1
X_100_ FrameStrobe[3] VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__clkbuf_1
XFILLER_8_44 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput147 net148 VGND VGND VPWR VPWR NN4BEG[3] sky130_fd_sc_hd__buf_2
Xoutput125 net126 VGND VGND VPWR VPWR N4BEG[12] sky130_fd_sc_hd__buf_2
Xoutput136 net137 VGND VGND VPWR VPWR N4BEG[8] sky130_fd_sc_hd__buf_2
Xoutput103 net104 VGND VGND VPWR VPWR N1BEG[1] sky130_fd_sc_hd__buf_2
Xoutput114 net115 VGND VGND VPWR VPWR N2BEGb[0] sky130_fd_sc_hd__buf_2
XFILLER_1_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput38 SS4END[0] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__buf_1
Xinput27 S2MID[1] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__buf_1
Xinput16 S1END[2] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__buf_1
XFILLER_6_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_56 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_030_ net18 Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit29.Q Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit30.Q
+ VGND VGND VPWR VPWR _006_ sky130_fd_sc_hd__o21ba_1
X_159_ SS4END[9] VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__buf_1
XFILLER_0_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput126 net127 VGND VGND VPWR VPWR N4BEG[13] sky130_fd_sc_hd__buf_2
Xoutput115 net116 VGND VGND VPWR VPWR N2BEGb[1] sky130_fd_sc_hd__buf_2
Xoutput104 net105 VGND VGND VPWR VPWR N1BEG[2] sky130_fd_sc_hd__buf_2
Xoutput148 net149 VGND VGND VPWR VPWR NN4BEG[4] sky130_fd_sc_hd__buf_2
Xoutput137 net138 VGND VGND VPWR VPWR N4BEG[9] sky130_fd_sc_hd__buf_2
XFILLER_9_363 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput39 SS4END[1] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput28 S2MID[2] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__buf_1
Xinput17 S1END[3] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__buf_1
XFILLER_6_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_158_ SS4END[10] VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__buf_1
XFILLER_8_68 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_089_ net6 VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__clkbuf_2
XFILLER_3_100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_375 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput149 net150 VGND VGND VPWR VPWR NN4BEG[5] sky130_fd_sc_hd__buf_2
Xoutput138 net139 VGND VGND VPWR VPWR NN4BEG[0] sky130_fd_sc_hd__buf_2
XFILLER_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput127 net128 VGND VGND VPWR VPWR N4BEG[14] sky130_fd_sc_hd__buf_2
Xoutput116 net117 VGND VGND VPWR VPWR N2BEGb[2] sky130_fd_sc_hd__buf_2
Xoutput105 net106 VGND VGND VPWR VPWR N1BEG[3] sky130_fd_sc_hd__buf_2
Xinput18 S2END[0] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__buf_1
Xinput29 S2MID[3] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__buf_1
XFILLER_10_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_157_ SS4END[11] VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__buf_1
XFILLER_6_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_088_ net5 VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_8_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput128 net129 VGND VGND VPWR VPWR N4BEG[15] sky130_fd_sc_hd__buf_2
Xoutput117 net118 VGND VGND VPWR VPWR N2BEGb[3] sky130_fd_sc_hd__buf_2
Xoutput106 net107 VGND VGND VPWR VPWR N2BEG[0] sky130_fd_sc_hd__buf_2
Xoutput139 net140 VGND VGND VPWR VPWR NN4BEG[10] sky130_fd_sc_hd__buf_2
XFILLER_9_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput19 S2END[1] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_1_Left_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_156_ SS4END[12] VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__buf_1
XFILLER_8_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_087_ net4 VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_8_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_139_ S4END[13] VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__buf_1
XFILLER_0_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput129 net130 VGND VGND VPWR VPWR N4BEG[1] sky130_fd_sc_hd__buf_2
Xoutput118 net119 VGND VGND VPWR VPWR N2BEGb[4] sky130_fd_sc_hd__buf_2
Xoutput107 net108 VGND VGND VPWR VPWR N2BEG[1] sky130_fd_sc_hd__buf_2
XFILLER_9_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_155_ SS4END[13] VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__buf_1
XFILLER_6_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_086_ net2 VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_8_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_138_ S4END[14] VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__buf_1
X_069_ FrameData[4] VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__clkbuf_1
XFILLER_9_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput90 net91 VGND VGND VPWR VPWR FrameStrobe_O[2] sky130_fd_sc_hd__buf_2
Xoutput119 net120 VGND VGND VPWR VPWR N2BEGb[5] sky130_fd_sc_hd__buf_2
Xoutput108 net109 VGND VGND VPWR VPWR N2BEG[2] sky130_fd_sc_hd__buf_2
XFILLER_9_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_154_ SS4END[14] VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_8_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_085_ net1 VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__buf_1
XFILLER_6_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_137_ S4END[15] VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__buf_1
X_068_ FrameData[3] VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__clkbuf_1
XFILLER_9_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_72 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput109 net110 VGND VGND VPWR VPWR N2BEG[3] sky130_fd_sc_hd__buf_2
XFILLER_9_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput91 net92 VGND VGND VPWR VPWR FrameStrobe_O[3] sky130_fd_sc_hd__buf_2
Xoutput80 net81 VGND VGND VPWR VPWR FrameStrobe_O[11] sky130_fd_sc_hd__buf_2
XFILLER_10_312 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_5_Left_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_084_ FrameData[19] VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__clkbuf_1
X_153_ SS4END[15] VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__buf_1
XFILLER_6_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_330 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_136_ net19 VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__buf_1
XFILLER_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_182 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_067_ FrameData[2] VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_8_Left_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_119_ net16 VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__clkbuf_1
XFILLER_7_252 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput81 net82 VGND VGND VPWR VPWR FrameStrobe_O[12] sky130_fd_sc_hd__buf_2
Xoutput92 net93 VGND VGND VPWR VPWR FrameStrobe_O[4] sky130_fd_sc_hd__buf_2
XFILLER_11_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput70 net71 VGND VGND VPWR VPWR FrameData_O[31] sky130_fd_sc_hd__buf_2
XFILLER_10_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_339 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_199 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_30 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_083_ FrameData[18] VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__clkbuf_2
X_152_ net31 VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__clkbuf_1
XFILLER_6_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_342 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_40 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_135_ net20 VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_066_ FrameData[1] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__clkbuf_2
XFILLER_11_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_264 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_118_ net17 VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__buf_1
X_049_ net19 net23 Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit20.Q VGND VGND VPWR VPWR
+ _022_ sky130_fd_sc_hd__mux2_1
Xfanout3 net14 VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_2
XFILLER_4_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_1 FrameData[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput93 net94 VGND VGND VPWR VPWR FrameStrobe_O[5] sky130_fd_sc_hd__buf_2
Xoutput60 net61 VGND VGND VPWR VPWR FrameData_O[22] sky130_fd_sc_hd__buf_2
Xoutput82 net83 VGND VGND VPWR VPWR FrameStrobe_O[13] sky130_fd_sc_hd__buf_2
XFILLER_9_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput71 net72 VGND VGND VPWR VPWR FrameData_O[3] sky130_fd_sc_hd__buf_2
XFILLER_10_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_336 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_340 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_166 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_082_ FrameData[17] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__clkbuf_2
X_151_ net32 VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__clkbuf_1
XFILLER_2_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_134_ net21 VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__clkbuf_1
X_065_ FrameData[0] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__clkbuf_1
XFILLER_9_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_117_ net18 VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__buf_1
X_048_ net15 Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit20.Q Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit21.Q
+ VGND VGND VPWR VPWR _021_ sky130_fd_sc_hd__o21ba_1
XFILLER_7_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_2 FrameData[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput83 net84 VGND VGND VPWR VPWR FrameStrobe_O[14] sky130_fd_sc_hd__buf_2
Xoutput94 net95 VGND VGND VPWR VPWR FrameStrobe_O[6] sky130_fd_sc_hd__buf_2
Xoutput61 net62 VGND VGND VPWR VPWR FrameData_O[23] sky130_fd_sc_hd__buf_2
XFILLER_9_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput50 net51 VGND VGND VPWR VPWR FrameData_O[13] sky130_fd_sc_hd__buf_2
XFILLER_0_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput72 net73 VGND VGND VPWR VPWR FrameData_O[4] sky130_fd_sc_hd__buf_2
XFILLER_10_348 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_352 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_081_ FrameData[16] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__clkbuf_2
XFILLER_2_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_150_ net33 VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__clkbuf_1
XFILLER_2_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_133_ net22 VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__buf_1
XFILLER_7_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_047_ net27 Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit20.Q VGND VGND VPWR VPWR _020_
+ sky130_fd_sc_hd__nand2b_1
X_116_ FrameStrobe[19] VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_3 FrameData[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_32 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput62 net63 VGND VGND VPWR VPWR FrameData_O[24] sky130_fd_sc_hd__buf_2
Xoutput84 net85 VGND VGND VPWR VPWR FrameStrobe_O[15] sky130_fd_sc_hd__buf_2
Xoutput95 net96 VGND VGND VPWR VPWR FrameStrobe_O[7] sky130_fd_sc_hd__buf_2
XFILLER_9_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput73 net74 VGND VGND VPWR VPWR FrameData_O[5] sky130_fd_sc_hd__buf_2
Xoutput51 net52 VGND VGND VPWR VPWR FrameData_O[14] sky130_fd_sc_hd__buf_2
XFILLER_6_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_364 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_080_ FrameData[15] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__clkbuf_1
XFILLER_8_180 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_063_ net13 net14 VGND VGND VPWR VPWR Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
X_132_ net23 VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__clkbuf_1
XFILLER_2_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_115_ FrameStrobe[18] VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__clkbuf_1
X_046_ net31 net35 net39 net43 Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit20.Q Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit21.Q
+ VGND VGND VPWR VPWR _019_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_5_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_4 FrameData[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_44 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_029_ net30 Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit29.Q VGND VGND VPWR VPWR _005_
+ sky130_fd_sc_hd__nand2b_1
XFILLER_3_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput52 net53 VGND VGND VPWR VPWR FrameData_O[15] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_2_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput85 net86 VGND VGND VPWR VPWR FrameStrobe_O[16] sky130_fd_sc_hd__buf_2
Xoutput96 net97 VGND VGND VPWR VPWR FrameStrobe_O[8] sky130_fd_sc_hd__buf_2
Xoutput63 net64 VGND VGND VPWR VPWR FrameData_O[25] sky130_fd_sc_hd__buf_2
Xoutput74 net75 VGND VGND VPWR VPWR FrameData_O[6] sky130_fd_sc_hd__buf_2
.ends

