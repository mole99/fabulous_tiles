* NGSPICE file created from N_term_single2.ext - technology: ihp-sg13g2

* Black-box entry subcircuit for sg13g2_decap_8 abstract view
.subckt sg13g2_decap_8 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_2 abstract view
.subckt sg13g2_fill_2 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_1 abstract view
.subckt sg13g2_buf_1 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_1 abstract view
.subckt sg13g2_fill_1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_antennanp abstract view
.subckt sg13g2_antennanp VDD VSS A
.ends

* Black-box entry subcircuit for sg13g2_decap_4 abstract view
.subckt sg13g2_decap_4 VDD VSS
.ends

.subckt N_term_single2 FrameData[0] FrameData[10] FrameData[11] FrameData[12] FrameData[13]
+ FrameData[14] FrameData[15] FrameData[16] FrameData[17] FrameData[18] FrameData[19]
+ FrameData[1] FrameData[20] FrameData[21] FrameData[22] FrameData[23] FrameData[24]
+ FrameData[25] FrameData[26] FrameData[27] FrameData[28] FrameData[29] FrameData[2]
+ FrameData[30] FrameData[31] FrameData[3] FrameData[4] FrameData[5] FrameData[6]
+ FrameData[7] FrameData[8] FrameData[9] FrameData_O[0] FrameData_O[10] FrameData_O[11]
+ FrameData_O[12] FrameData_O[13] FrameData_O[14] FrameData_O[15] FrameData_O[16]
+ FrameData_O[17] FrameData_O[18] FrameData_O[19] FrameData_O[1] FrameData_O[20] FrameData_O[21]
+ FrameData_O[22] FrameData_O[23] FrameData_O[24] FrameData_O[25] FrameData_O[26]
+ FrameData_O[27] FrameData_O[28] FrameData_O[29] FrameData_O[2] FrameData_O[30] FrameData_O[31]
+ FrameData_O[3] FrameData_O[4] FrameData_O[5] FrameData_O[6] FrameData_O[7] FrameData_O[8]
+ FrameData_O[9] FrameStrobe[0] FrameStrobe[10] FrameStrobe[11] FrameStrobe[12] FrameStrobe[13]
+ FrameStrobe[14] FrameStrobe[15] FrameStrobe[16] FrameStrobe[17] FrameStrobe[18]
+ FrameStrobe[19] FrameStrobe[1] FrameStrobe[2] FrameStrobe[3] FrameStrobe[4] FrameStrobe[5]
+ FrameStrobe[6] FrameStrobe[7] FrameStrobe[8] FrameStrobe[9] FrameStrobe_O[0] FrameStrobe_O[10]
+ FrameStrobe_O[11] FrameStrobe_O[12] FrameStrobe_O[13] FrameStrobe_O[14] FrameStrobe_O[15]
+ FrameStrobe_O[16] FrameStrobe_O[17] FrameStrobe_O[18] FrameStrobe_O[19] FrameStrobe_O[1]
+ FrameStrobe_O[2] FrameStrobe_O[3] FrameStrobe_O[4] FrameStrobe_O[5] FrameStrobe_O[6]
+ FrameStrobe_O[7] FrameStrobe_O[8] FrameStrobe_O[9] N1END[0] N1END[1] N1END[2] N1END[3]
+ N2END[0] N2END[1] N2END[2] N2END[3] N2END[4] N2END[5] N2END[6] N2END[7] N2MID[0]
+ N2MID[1] N2MID[2] N2MID[3] N2MID[4] N2MID[5] N2MID[6] N2MID[7] N4END[0] N4END[10]
+ N4END[11] N4END[12] N4END[13] N4END[14] N4END[15] N4END[1] N4END[2] N4END[3] N4END[4]
+ N4END[5] N4END[6] N4END[7] N4END[8] N4END[9] NN4END[0] NN4END[10] NN4END[11] NN4END[12]
+ NN4END[13] NN4END[14] NN4END[15] NN4END[1] NN4END[2] NN4END[3] NN4END[4] NN4END[5]
+ NN4END[6] NN4END[7] NN4END[8] NN4END[9] S1BEG[0] S1BEG[1] S1BEG[2] S1BEG[3] S2BEG[0]
+ S2BEG[1] S2BEG[2] S2BEG[3] S2BEG[4] S2BEG[5] S2BEG[6] S2BEG[7] S2BEGb[0] S2BEGb[1]
+ S2BEGb[2] S2BEGb[3] S2BEGb[4] S2BEGb[5] S2BEGb[6] S2BEGb[7] S4BEG[0] S4BEG[10] S4BEG[11]
+ S4BEG[12] S4BEG[13] S4BEG[14] S4BEG[15] S4BEG[1] S4BEG[2] S4BEG[3] S4BEG[4] S4BEG[5]
+ S4BEG[6] S4BEG[7] S4BEG[8] S4BEG[9] SS4BEG[0] SS4BEG[10] SS4BEG[11] SS4BEG[12] SS4BEG[13]
+ SS4BEG[14] SS4BEG[15] SS4BEG[1] SS4BEG[2] SS4BEG[3] SS4BEG[4] SS4BEG[5] SS4BEG[6]
+ SS4BEG[7] SS4BEG[8] SS4BEG[9] UserCLK UserCLKo VGND VPWR
XFILLER_10_306 VPWR VGND sg13g2_decap_8
XFILLER_7_7 VPWR VGND sg13g2_decap_8
XFILLER_2_505 VPWR VGND sg13g2_fill_2
XFILLER_9_126 VPWR VGND sg13g2_decap_8
XFILLER_5_387 VPWR VGND sg13g2_decap_8
XFILLER_3_56 VPWR VGND sg13g2_decap_8
XFILLER_10_147 VPWR VGND sg13g2_fill_2
XFILLER_5_140 VPWR VGND sg13g2_decap_8
XFILLER_9_490 VPWR VGND sg13g2_decap_8
XFILLER_7_416 VPWR VGND sg13g2_decap_8
X_062_ N2MID[1] net63 VPWR VGND sg13g2_buf_1
XFILLER_9_77 VPWR VGND sg13g2_decap_8
XFILLER_6_460 VPWR VGND sg13g2_decap_8
XFILLER_0_35 VPWR VGND sg13g2_decap_8
XFILLER_2_165 VPWR VGND sg13g2_fill_1
XFILLER_11_264 VPWR VGND sg13g2_fill_1
XFILLER_11_231 VPWR VGND sg13g2_decap_8
X_045_ FrameStrobe[13] net37 VPWR VGND sg13g2_buf_1
XFILLER_7_279 VPWR VGND sg13g2_decap_8
XFILLER_7_202 VPWR VGND sg13g2_decap_8
XFILLER_3_485 VPWR VGND sg13g2_decap_8
XFILLER_4_238 VPWR VGND sg13g2_fill_1
XFILLER_4_227 VPWR VGND sg13g2_decap_8
XFILLER_0_433 VPWR VGND sg13g2_decap_8
X_028_ FrameData[28] net21 VPWR VGND sg13g2_buf_1
XFILLER_6_56 VPWR VGND sg13g2_decap_8
XANTENNA_5 VPWR VGND net1 sg13g2_antennanp
XFILLER_9_319 VPWR VGND sg13g2_decap_8
Xoutput20 net20 FrameData_O[27] VPWR VGND sg13g2_buf_1
Xoutput42 net42 FrameStrobe_O[18] VPWR VGND sg13g2_buf_1
Xoutput7 net7 FrameData_O[15] VPWR VGND sg13g2_buf_1
Xoutput31 net31 FrameData_O[8] VPWR VGND sg13g2_buf_1
Xoutput53 net53 S1BEG[0] VPWR VGND sg13g2_buf_1
Xoutput64 net64 S2BEG[7] VPWR VGND sg13g2_buf_1
Xoutput86 net86 S4BEG[7] VPWR VGND sg13g2_buf_1
Xoutput75 net75 S4BEG[11] VPWR VGND sg13g2_buf_1
Xoutput97 net97 SS4BEG[2] VPWR VGND sg13g2_buf_1
XFILLER_11_0 VPWR VGND sg13g2_decap_4
XFILLER_9_105 VPWR VGND sg13g2_decap_8
XFILLER_5_366 VPWR VGND sg13g2_decap_8
XFILLER_5_344 VPWR VGND sg13g2_decap_8
XFILLER_3_35 VPWR VGND sg13g2_decap_8
XFILLER_8_182 VPWR VGND sg13g2_decap_8
XFILLER_10_126 VPWR VGND sg13g2_fill_2
XFILLER_6_119 VPWR VGND sg13g2_decap_8
XFILLER_2_369 VPWR VGND sg13g2_fill_1
XFILLER_5_196 VPWR VGND sg13g2_decap_8
XFILLER_1_380 VPWR VGND sg13g2_decap_8
XFILLER_11_446 VPWR VGND sg13g2_fill_1
XFILLER_11_413 VPWR VGND sg13g2_decap_8
XFILLER_9_56 VPWR VGND sg13g2_decap_8
X_061_ N2MID[2] net62 VPWR VGND sg13g2_buf_1
XFILLER_0_14 VPWR VGND sg13g2_decap_8
XFILLER_2_133 VPWR VGND sg13g2_fill_2
XFILLER_2_144 VPWR VGND sg13g2_decap_8
XFILLER_2_177 VPWR VGND sg13g2_decap_8
XFILLER_4_409 VPWR VGND sg13g2_decap_8
XFILLER_11_276 VPWR VGND sg13g2_decap_8
XFILLER_11_243 VPWR VGND sg13g2_decap_8
X_044_ FrameStrobe[12] net36 VPWR VGND sg13g2_buf_1
XFILLER_7_258 VPWR VGND sg13g2_decap_8
XFILLER_3_464 VPWR VGND sg13g2_decap_8
XFILLER_4_206 VPWR VGND sg13g2_decap_8
XFILLER_0_489 VPWR VGND sg13g2_decap_4
X_027_ FrameData[27] net20 VPWR VGND sg13g2_buf_1
XFILLER_8_512 VPWR VGND sg13g2_decap_8
XFILLER_6_35 VPWR VGND sg13g2_decap_8
XANTENNA_6 VPWR VGND net27 sg13g2_antennanp
XFILLER_3_283 VPWR VGND sg13g2_decap_8
XFILLER_1_209 VPWR VGND sg13g2_decap_8
Xoutput43 net43 FrameStrobe_O[19] VPWR VGND sg13g2_buf_1
Xoutput21 net21 FrameData_O[28] VPWR VGND sg13g2_buf_1
Xoutput10 net10 FrameData_O[18] VPWR VGND sg13g2_buf_1
Xoutput8 net8 FrameData_O[16] VPWR VGND sg13g2_buf_1
Xoutput54 net54 S1BEG[1] VPWR VGND sg13g2_buf_1
Xoutput65 net65 S2BEGb[0] VPWR VGND sg13g2_buf_1
Xoutput87 net87 S4BEG[8] VPWR VGND sg13g2_buf_1
Xoutput76 net76 S4BEG[12] VPWR VGND sg13g2_buf_1
Xoutput98 net98 SS4BEG[3] VPWR VGND sg13g2_buf_1
Xoutput32 net32 FrameData_O[9] VPWR VGND sg13g2_buf_1
XFILLER_8_386 VPWR VGND sg13g2_decap_8
XFILLER_8_353 VPWR VGND sg13g2_fill_1
XFILLER_5_323 VPWR VGND sg13g2_decap_8
XFILLER_8_161 VPWR VGND sg13g2_decap_8
XFILLER_3_14 VPWR VGND sg13g2_decap_8
XFILLER_10_105 VPWR VGND sg13g2_decap_8
XFILLER_5_175 VPWR VGND sg13g2_decap_8
XFILLER_11_458 VPWR VGND sg13g2_decap_8
XFILLER_11_425 VPWR VGND sg13g2_decap_8
XFILLER_9_35 VPWR VGND sg13g2_decap_8
X_060_ N2MID[3] net61 VPWR VGND sg13g2_buf_1
XFILLER_2_112 VPWR VGND sg13g2_decap_8
XFILLER_6_495 VPWR VGND sg13g2_decap_8
X_043_ FrameStrobe[11] net35 VPWR VGND sg13g2_buf_1
XFILLER_7_237 VPWR VGND sg13g2_decap_8
XFILLER_6_281 VPWR VGND sg13g2_decap_8
XFILLER_3_443 VPWR VGND sg13g2_decap_8
XFILLER_1_0 VPWR VGND sg13g2_decap_8
X_026_ FrameData[26] net19 VPWR VGND sg13g2_buf_1
XANTENNA_7 VPWR VGND FrameStrobe[3] sg13g2_antennanp
XFILLER_6_14 VPWR VGND sg13g2_decap_8
XFILLER_0_468 VPWR VGND sg13g2_decap_8
XFILLER_3_273 VPWR VGND sg13g2_decap_4
Xoutput22 net22 FrameData_O[29] VPWR VGND sg13g2_buf_1
Xoutput44 net44 FrameStrobe_O[1] VPWR VGND sg13g2_buf_1
Xoutput33 net33 FrameStrobe_O[0] VPWR VGND sg13g2_buf_1
Xoutput11 net11 FrameData_O[19] VPWR VGND sg13g2_buf_1
Xoutput9 net9 FrameData_O[17] VPWR VGND sg13g2_buf_1
Xoutput55 net55 S1BEG[2] VPWR VGND sg13g2_buf_1
XFILLER_0_210 VPWR VGND sg13g2_decap_8
Xoutput66 net66 S2BEGb[1] VPWR VGND sg13g2_buf_1
Xoutput88 net88 S4BEG[9] VPWR VGND sg13g2_buf_1
Xoutput77 net77 S4BEG[13] VPWR VGND sg13g2_buf_1
Xoutput99 net99 SS4BEG[4] VPWR VGND sg13g2_buf_1
X_009_ FrameData[9] net32 VPWR VGND sg13g2_buf_1
XFILLER_8_365 VPWR VGND sg13g2_decap_8
XFILLER_2_519 VPWR VGND sg13g2_fill_1
XFILLER_8_140 VPWR VGND sg13g2_decap_8
XFILLER_5_302 VPWR VGND sg13g2_decap_8
XFILLER_10_128 VPWR VGND sg13g2_fill_1
XFILLER_5_7 VPWR VGND sg13g2_decap_8
XFILLER_2_316 VPWR VGND sg13g2_fill_1
XFILLER_2_338 VPWR VGND sg13g2_fill_1
XFILLER_5_154 VPWR VGND sg13g2_decap_8
XFILLER_4_91 VPWR VGND sg13g2_decap_8
XFILLER_0_49 VPWR VGND sg13g2_decap_8
XFILLER_9_14 VPWR VGND sg13g2_decap_8
XFILLER_6_474 VPWR VGND sg13g2_decap_8
XFILLER_11_212 VPWR VGND sg13g2_fill_1
X_042_ FrameStrobe[10] net34 VPWR VGND sg13g2_buf_1
XFILLER_7_216 VPWR VGND sg13g2_decap_8
XFILLER_3_499 VPWR VGND sg13g2_decap_8
XFILLER_3_422 VPWR VGND sg13g2_decap_8
XFILLER_6_260 VPWR VGND sg13g2_decap_8
XFILLER_1_81 VPWR VGND sg13g2_decap_8
X_025_ FrameData[25] net18 VPWR VGND sg13g2_buf_1
XANTENNA_8 VPWR VGND FrameStrobe[4] sg13g2_antennanp
XFILLER_0_447 VPWR VGND sg13g2_decap_8
XFILLER_3_252 VPWR VGND sg13g2_decap_8
Xoutput34 net34 FrameStrobe_O[10] VPWR VGND sg13g2_buf_1
Xoutput45 net45 FrameStrobe_O[2] VPWR VGND sg13g2_buf_1
XFILLER_5_506 VPWR VGND sg13g2_decap_8
Xoutput56 net56 S1BEG[3] VPWR VGND sg13g2_buf_1
Xoutput67 net67 S2BEGb[2] VPWR VGND sg13g2_buf_1
Xoutput78 net78 S4BEG[14] VPWR VGND sg13g2_buf_1
Xoutput89 net89 SS4BEG[0] VPWR VGND sg13g2_buf_1
Xoutput12 net12 FrameData_O[1] VPWR VGND sg13g2_buf_1
Xoutput23 net23 FrameData_O[2] VPWR VGND sg13g2_buf_1
XFILLER_8_333 VPWR VGND sg13g2_fill_2
XFILLER_8_311 VPWR VGND sg13g2_decap_4
X_008_ FrameData[8] net31 VPWR VGND sg13g2_buf_1
XFILLER_7_91 VPWR VGND sg13g2_decap_8
XFILLER_9_119 VPWR VGND sg13g2_decap_8
XFILLER_5_358 VPWR VGND sg13g2_fill_2
XFILLER_3_49 VPWR VGND sg13g2_decap_8
XFILLER_8_196 VPWR VGND sg13g2_decap_8
XFILLER_5_133 VPWR VGND sg13g2_decap_8
XFILLER_9_483 VPWR VGND sg13g2_decap_8
XFILLER_1_394 VPWR VGND sg13g2_fill_2
XFILLER_7_409 VPWR VGND sg13g2_decap_8
XFILLER_4_70 VPWR VGND sg13g2_decap_8
XFILLER_2_158 VPWR VGND sg13g2_decap_8
XFILLER_10_482 VPWR VGND sg13g2_decap_8
XFILLER_10_460 VPWR VGND sg13g2_decap_8
XFILLER_6_453 VPWR VGND sg13g2_decap_8
XFILLER_0_28 VPWR VGND sg13g2_decap_8
XFILLER_9_291 VPWR VGND sg13g2_decap_8
XFILLER_11_257 VPWR VGND sg13g2_decap_8
XFILLER_11_224 VPWR VGND sg13g2_decap_8
X_041_ FrameStrobe[9] net52 VPWR VGND sg13g2_buf_1
XFILLER_3_478 VPWR VGND sg13g2_decap_8
XFILLER_3_401 VPWR VGND sg13g2_decap_8
XFILLER_10_91 VPWR VGND sg13g2_decap_8
X_024_ FrameData[24] net17 VPWR VGND sg13g2_buf_1
XANTENNA_9 VPWR VGND FrameData[10] sg13g2_antennanp
XFILLER_6_49 VPWR VGND sg13g2_decap_8
XFILLER_3_231 VPWR VGND sg13g2_decap_8
XFILLER_3_297 VPWR VGND sg13g2_decap_8
Xoutput24 net24 FrameData_O[30] VPWR VGND sg13g2_buf_1
Xoutput35 net35 FrameStrobe_O[11] VPWR VGND sg13g2_buf_1
Xoutput46 net46 FrameStrobe_O[3] VPWR VGND sg13g2_buf_1
Xoutput13 net13 FrameData_O[20] VPWR VGND sg13g2_buf_1
Xoutput57 net57 S2BEG[0] VPWR VGND sg13g2_buf_1
X_007_ FrameData[7] net30 VPWR VGND sg13g2_buf_1
Xoutput68 net68 S2BEGb[3] VPWR VGND sg13g2_buf_1
Xoutput79 net79 S4BEG[15] VPWR VGND sg13g2_buf_1
XFILLER_11_4 VPWR VGND sg13g2_fill_1
XFILLER_7_70 VPWR VGND sg13g2_decap_8
XFILLER_5_337 VPWR VGND sg13g2_decap_8
XFILLER_3_28 VPWR VGND sg13g2_decap_8
XFILLER_8_175 VPWR VGND sg13g2_decap_8
XFILLER_4_381 VPWR VGND sg13g2_decap_8
XFILLER_10_119 VPWR VGND sg13g2_decap_8
XFILLER_2_329 VPWR VGND sg13g2_fill_1
XFILLER_9_462 VPWR VGND sg13g2_decap_8
XFILLER_5_189 VPWR VGND sg13g2_decap_8
XFILLER_5_112 VPWR VGND sg13g2_decap_8
XFILLER_1_373 VPWR VGND sg13g2_decap_8
XFILLER_11_439 VPWR VGND sg13g2_decap_8
XFILLER_11_406 VPWR VGND sg13g2_decap_8
XFILLER_10_450 VPWR VGND sg13g2_decap_4
XFILLER_9_49 VPWR VGND sg13g2_decap_8
XFILLER_6_432 VPWR VGND sg13g2_decap_8
XFILLER_2_126 VPWR VGND sg13g2_decap_8
XFILLER_1_192 VPWR VGND sg13g2_decap_8
XFILLER_11_269 VPWR VGND sg13g2_decap_8
X_040_ FrameStrobe[8] net51 VPWR VGND sg13g2_buf_1
XFILLER_3_457 VPWR VGND sg13g2_decap_8
XFILLER_6_295 VPWR VGND sg13g2_decap_8
XFILLER_6_251 VPWR VGND sg13g2_fill_1
XFILLER_10_70 VPWR VGND sg13g2_decap_8
XFILLER_8_505 VPWR VGND sg13g2_decap_8
X_023_ FrameData[23] net16 VPWR VGND sg13g2_buf_1
XFILLER_6_28 VPWR VGND sg13g2_decap_8
Xoutput36 net36 FrameStrobe_O[12] VPWR VGND sg13g2_buf_1
Xoutput47 net47 FrameStrobe_O[4] VPWR VGND sg13g2_buf_1
Xoutput25 net25 FrameData_O[31] VPWR VGND sg13g2_buf_1
Xoutput14 net14 FrameData_O[21] VPWR VGND sg13g2_buf_1
XFILLER_8_379 VPWR VGND sg13g2_decap_8
XFILLER_8_346 VPWR VGND sg13g2_decap_8
XFILLER_8_335 VPWR VGND sg13g2_fill_1
X_006_ FrameData[6] net29 VPWR VGND sg13g2_buf_1
Xoutput58 net58 S2BEG[1] VPWR VGND sg13g2_buf_1
XFILLER_0_224 VPWR VGND sg13g2_fill_1
Xoutput69 net69 S2BEGb[4] VPWR VGND sg13g2_buf_1
XFILLER_5_316 VPWR VGND sg13g2_decap_8
XFILLER_8_154 VPWR VGND sg13g2_decap_8
XFILLER_4_360 VPWR VGND sg13g2_decap_8
XFILLER_5_168 VPWR VGND sg13g2_decap_8
XFILLER_1_352 VPWR VGND sg13g2_decap_8
XFILLER_1_396 VPWR VGND sg13g2_fill_1
XFILLER_9_441 VPWR VGND sg13g2_decap_8
XFILLER_10_473 VPWR VGND sg13g2_fill_1
XFILLER_9_28 VPWR VGND sg13g2_decap_8
XFILLER_6_411 VPWR VGND sg13g2_decap_8
XFILLER_2_105 VPWR VGND sg13g2_decap_8
XFILLER_3_7 VPWR VGND sg13g2_decap_8
XFILLER_6_488 VPWR VGND sg13g2_decap_8
XFILLER_3_436 VPWR VGND sg13g2_decap_8
XFILLER_10_292 VPWR VGND sg13g2_decap_4
XFILLER_6_274 VPWR VGND sg13g2_decap_8
X_099_ NN4END[4] net91 VPWR VGND sg13g2_buf_1
XFILLER_2_491 VPWR VGND sg13g2_decap_8
XFILLER_1_95 VPWR VGND sg13g2_decap_8
X_022_ FrameData[22] net15 VPWR VGND sg13g2_buf_1
XFILLER_3_266 VPWR VGND sg13g2_decap_8
XFILLER_3_277 VPWR VGND sg13g2_fill_2
Xoutput37 net37 FrameStrobe_O[13] VPWR VGND sg13g2_buf_1
Xoutput48 net48 FrameStrobe_O[5] VPWR VGND sg13g2_buf_1
Xoutput15 net15 FrameData_O[22] VPWR VGND sg13g2_buf_1
Xoutput59 net59 S2BEG[2] VPWR VGND sg13g2_buf_1
XFILLER_0_203 VPWR VGND sg13g2_decap_8
Xoutput26 net26 FrameData_O[3] VPWR VGND sg13g2_buf_1
XFILLER_8_358 VPWR VGND sg13g2_decap_8
X_005_ FrameData[5] net28 VPWR VGND sg13g2_buf_1
XFILLER_8_133 VPWR VGND sg13g2_decap_8
XFILLER_5_147 VPWR VGND sg13g2_decap_8
XFILLER_9_497 VPWR VGND sg13g2_decap_8
XFILLER_9_420 VPWR VGND sg13g2_decap_8
XFILLER_4_84 VPWR VGND sg13g2_decap_8
XFILLER_2_139 VPWR VGND sg13g2_fill_1
XFILLER_6_467 VPWR VGND sg13g2_decap_8
XFILLER_1_172 VPWR VGND sg13g2_decap_4
XFILLER_11_238 VPWR VGND sg13g2_fill_1
XFILLER_11_205 VPWR VGND sg13g2_decap_8
XFILLER_9_272 VPWR VGND sg13g2_decap_4
XFILLER_7_209 VPWR VGND sg13g2_decap_8
XFILLER_10_282 VPWR VGND sg13g2_decap_4
XFILLER_6_242 VPWR VGND sg13g2_decap_8
XFILLER_3_415 VPWR VGND sg13g2_decap_8
X_098_ NN4END[5] net90 VPWR VGND sg13g2_buf_1
XFILLER_1_74 VPWR VGND sg13g2_decap_8
XFILLER_2_470 VPWR VGND sg13g2_decap_8
X_021_ FrameData[21] net14 VPWR VGND sg13g2_buf_1
XFILLER_3_212 VPWR VGND sg13g2_decap_8
XFILLER_3_245 VPWR VGND sg13g2_decap_8
Xoutput38 net38 FrameStrobe_O[14] VPWR VGND sg13g2_buf_1
Xoutput49 net49 FrameStrobe_O[6] VPWR VGND sg13g2_buf_1
Xoutput16 net16 FrameData_O[23] VPWR VGND sg13g2_buf_1
Xoutput27 net27 FrameData_O[4] VPWR VGND sg13g2_buf_1
XFILLER_8_326 VPWR VGND sg13g2_decap_8
XFILLER_8_304 VPWR VGND sg13g2_decap_8
XFILLER_4_521 VPWR VGND sg13g2_fill_2
X_004_ FrameData[4] net27 VPWR VGND sg13g2_buf_1
XFILLER_7_381 VPWR VGND sg13g2_decap_8
XFILLER_7_84 VPWR VGND sg13g2_decap_8
XFILLER_8_189 VPWR VGND sg13g2_decap_8
XFILLER_8_112 VPWR VGND sg13g2_decap_8
XFILLER_4_395 VPWR VGND sg13g2_decap_8
XFILLER_5_126 VPWR VGND sg13g2_decap_8
XFILLER_1_343 VPWR VGND sg13g2_fill_1
XFILLER_9_476 VPWR VGND sg13g2_decap_8
XFILLER_4_192 VPWR VGND sg13g2_decap_8
XFILLER_4_63 VPWR VGND sg13g2_decap_8
XFILLER_1_387 VPWR VGND sg13g2_decap_8
XFILLER_6_446 VPWR VGND sg13g2_decap_8
XFILLER_1_151 VPWR VGND sg13g2_decap_8
XFILLER_11_217 VPWR VGND sg13g2_decap_8
XFILLER_9_284 VPWR VGND sg13g2_decap_8
XFILLER_10_250 VPWR VGND sg13g2_fill_2
XFILLER_6_210 VPWR VGND sg13g2_decap_8
XFILLER_1_42 VPWR VGND sg13g2_decap_8
X_097_ NN4END[6] net104 VPWR VGND sg13g2_buf_1
XFILLER_8_519 VPWR VGND sg13g2_decap_4
X_020_ FrameData[20] net13 VPWR VGND sg13g2_buf_1
XFILLER_10_84 VPWR VGND sg13g2_decap_8
Xoutput39 net39 FrameStrobe_O[15] VPWR VGND sg13g2_buf_1
Xoutput17 net17 FrameData_O[24] VPWR VGND sg13g2_buf_1
Xoutput28 net28 FrameData_O[5] VPWR VGND sg13g2_buf_1
XFILLER_4_500 VPWR VGND sg13g2_decap_8
X_003_ FrameData[3] net26 VPWR VGND sg13g2_buf_1
XFILLER_7_360 VPWR VGND sg13g2_decap_8
XFILLER_7_63 VPWR VGND sg13g2_decap_8
XFILLER_8_168 VPWR VGND sg13g2_decap_8
XFILLER_4_374 VPWR VGND sg13g2_decap_8
XFILLER_5_105 VPWR VGND sg13g2_decap_8
XFILLER_9_455 VPWR VGND sg13g2_decap_8
XFILLER_4_171 VPWR VGND sg13g2_decap_8
XFILLER_4_42 VPWR VGND sg13g2_decap_8
XFILLER_1_333 VPWR VGND sg13g2_fill_2
XFILLER_1_366 VPWR VGND sg13g2_decap_8
XFILLER_2_119 VPWR VGND sg13g2_decap_8
XFILLER_10_498 VPWR VGND sg13g2_decap_8
XFILLER_10_454 VPWR VGND sg13g2_fill_2
XFILLER_8_0 VPWR VGND sg13g2_decap_8
XFILLER_6_425 VPWR VGND sg13g2_decap_8
XFILLER_1_185 VPWR VGND sg13g2_decap_8
XFILLER_9_252 VPWR VGND sg13g2_fill_2
XFILLER_1_7 VPWR VGND sg13g2_fill_2
XFILLER_6_288 VPWR VGND sg13g2_decap_8
X_096_ NN4END[7] net103 VPWR VGND sg13g2_buf_1
XFILLER_1_21 VPWR VGND sg13g2_decap_8
XFILLER_10_63 VPWR VGND sg13g2_decap_8
Xoutput18 net18 FrameData_O[25] VPWR VGND sg13g2_buf_1
XFILLER_0_217 VPWR VGND sg13g2_decap_8
Xoutput29 net29 FrameData_O[6] VPWR VGND sg13g2_buf_1
X_079_ N4END[8] net86 VPWR VGND sg13g2_buf_1
XFILLER_8_339 VPWR VGND sg13g2_decap_8
X_002_ FrameData[2] net23 VPWR VGND sg13g2_buf_1
XFILLER_11_9 VPWR VGND sg13g2_decap_8
XFILLER_7_42 VPWR VGND sg13g2_decap_8
XFILLER_5_309 VPWR VGND sg13g2_decap_8
XFILLER_8_147 VPWR VGND sg13g2_decap_8
XFILLER_4_353 VPWR VGND sg13g2_decap_8
XFILLER_9_434 VPWR VGND sg13g2_decap_8
XFILLER_1_312 VPWR VGND sg13g2_decap_8
XFILLER_4_150 VPWR VGND sg13g2_decap_8
XFILLER_4_98 VPWR VGND sg13g2_decap_8
XFILLER_4_21 VPWR VGND sg13g2_decap_8
XFILLER_10_444 VPWR VGND sg13g2_fill_2
XFILLER_6_404 VPWR VGND sg13g2_decap_8
XFILLER_9_231 VPWR VGND sg13g2_decap_8
XFILLER_5_492 VPWR VGND sg13g2_decap_8
XFILLER_3_429 VPWR VGND sg13g2_decap_8
XFILLER_10_296 VPWR VGND sg13g2_fill_1
XFILLER_6_267 VPWR VGND sg13g2_decap_8
XFILLER_1_88 VPWR VGND sg13g2_decap_8
XFILLER_2_484 VPWR VGND sg13g2_decap_8
X_095_ NN4END[8] net102 VPWR VGND sg13g2_buf_1
XFILLER_10_42 VPWR VGND sg13g2_decap_8
XFILLER_3_226 VPWR VGND sg13g2_fill_1
XFILLER_3_259 VPWR VGND sg13g2_decap_8
XFILLER_7_521 VPWR VGND sg13g2_fill_2
XFILLER_2_292 VPWR VGND sg13g2_decap_4
X_078_ N4END[9] net85 VPWR VGND sg13g2_buf_1
Xoutput19 net19 FrameData_O[26] VPWR VGND sg13g2_buf_1
X_001_ FrameData[1] net12 VPWR VGND sg13g2_buf_1
XFILLER_11_380 VPWR VGND sg13g2_decap_8
XFILLER_7_395 VPWR VGND sg13g2_decap_8
XFILLER_7_98 VPWR VGND sg13g2_decap_8
XFILLER_7_21 VPWR VGND sg13g2_decap_8
XFILLER_8_126 VPWR VGND sg13g2_decap_8
XFILLER_4_332 VPWR VGND sg13g2_decap_8
XFILLER_9_413 VPWR VGND sg13g2_decap_8
XFILLER_4_77 VPWR VGND sg13g2_decap_8
XFILLER_10_489 VPWR VGND sg13g2_fill_1
XFILLER_10_467 VPWR VGND sg13g2_fill_2
XFILLER_9_298 VPWR VGND sg13g2_decap_8
XFILLER_9_265 VPWR VGND sg13g2_decap_8
XFILLER_9_210 VPWR VGND sg13g2_decap_8
XFILLER_5_471 VPWR VGND sg13g2_decap_8
XFILLER_1_176 VPWR VGND sg13g2_fill_1
XFILLER_1_165 VPWR VGND sg13g2_decap_8
XFILLER_1_132 VPWR VGND sg13g2_fill_2
XFILLER_1_121 VPWR VGND sg13g2_fill_2
XFILLER_3_408 VPWR VGND sg13g2_decap_8
XFILLER_1_9 VPWR VGND sg13g2_fill_1
XFILLER_10_286 VPWR VGND sg13g2_fill_2
XFILLER_10_264 VPWR VGND sg13g2_fill_1
XFILLER_6_235 VPWR VGND sg13g2_decap_8
X_094_ NN4END[9] net101 VPWR VGND sg13g2_buf_1
XFILLER_2_463 VPWR VGND sg13g2_decap_8
XFILLER_1_67 VPWR VGND sg13g2_decap_8
XFILLER_1_56 VPWR VGND sg13g2_decap_8
XFILLER_10_98 VPWR VGND sg13g2_decap_8
XFILLER_10_21 VPWR VGND sg13g2_decap_8
XFILLER_3_205 VPWR VGND sg13g2_decap_8
XFILLER_3_238 VPWR VGND sg13g2_decap_8
XFILLER_7_500 VPWR VGND sg13g2_decap_8
X_077_ N4END[10] net84 VPWR VGND sg13g2_buf_1
XFILLER_8_319 VPWR VGND sg13g2_decap_8
XFILLER_7_374 VPWR VGND sg13g2_decap_8
XFILLER_7_352 VPWR VGND sg13g2_fill_2
XFILLER_7_341 VPWR VGND sg13g2_decap_8
XFILLER_7_77 VPWR VGND sg13g2_decap_8
XFILLER_4_514 VPWR VGND sg13g2_decap_8
X_000_ FrameData[0] net1 VPWR VGND sg13g2_buf_1
XFILLER_8_105 VPWR VGND sg13g2_decap_8
XFILLER_4_388 VPWR VGND sg13g2_decap_8
XFILLER_4_311 VPWR VGND sg13g2_decap_8
XFILLER_7_182 VPWR VGND sg13g2_fill_2
XFILLER_5_119 VPWR VGND sg13g2_decap_8
XFILLER_9_469 VPWR VGND sg13g2_decap_8
XFILLER_4_185 VPWR VGND sg13g2_decap_8
XFILLER_4_56 VPWR VGND sg13g2_decap_8
XFILLER_8_491 VPWR VGND sg13g2_decap_8
XFILLER_10_435 VPWR VGND sg13g2_decap_4
XFILLER_6_439 VPWR VGND sg13g2_decap_8
XFILLER_1_199 VPWR VGND sg13g2_fill_2
XFILLER_1_144 VPWR VGND sg13g2_decap_8
XFILLER_5_450 VPWR VGND sg13g2_decap_8
XFILLER_10_276 VPWR VGND sg13g2_fill_2
XFILLER_6_203 VPWR VGND sg13g2_decap_8
XFILLER_6_0 VPWR VGND sg13g2_decap_8
X_093_ NN4END[10] net100 VPWR VGND sg13g2_buf_1
XFILLER_1_35 VPWR VGND sg13g2_decap_8
XFILLER_10_77 VPWR VGND sg13g2_decap_8
XFILLER_2_261 VPWR VGND sg13g2_decap_8
X_076_ N4END[11] net83 VPWR VGND sg13g2_buf_1
XANTENNA_50 VPWR VGND net1 sg13g2_antennanp
XFILLER_7_320 VPWR VGND sg13g2_decap_8
XFILLER_7_56 VPWR VGND sg13g2_decap_8
X_059_ N2MID[4] net60 VPWR VGND sg13g2_buf_1
XFILLER_7_161 VPWR VGND sg13g2_decap_8
XFILLER_4_367 VPWR VGND sg13g2_decap_8
XFILLER_1_326 VPWR VGND sg13g2_decap_8
XFILLER_1_359 VPWR VGND sg13g2_decap_8
XFILLER_9_448 VPWR VGND sg13g2_decap_8
XFILLER_4_164 VPWR VGND sg13g2_decap_8
XFILLER_4_35 VPWR VGND sg13g2_decap_8
XFILLER_8_470 VPWR VGND sg13g2_decap_8
XFILLER_10_425 VPWR VGND sg13g2_decap_4
XFILLER_6_418 VPWR VGND sg13g2_decap_8
XFILLER_1_123 VPWR VGND sg13g2_fill_1
XFILLER_9_245 VPWR VGND sg13g2_decap_8
XFILLER_10_233 VPWR VGND sg13g2_fill_2
XFILLER_1_14 VPWR VGND sg13g2_decap_8
X_092_ NN4END[11] net99 VPWR VGND sg13g2_buf_1
XFILLER_2_410 VPWR VGND sg13g2_decap_8
XFILLER_2_421 VPWR VGND sg13g2_fill_1
XFILLER_2_498 VPWR VGND sg13g2_decap_8
XFILLER_10_56 VPWR VGND sg13g2_decap_8
XFILLER_5_281 VPWR VGND sg13g2_decap_8
X_075_ N4END[12] net82 VPWR VGND sg13g2_buf_1
XFILLER_2_240 VPWR VGND sg13g2_decap_8
XANTENNA_51 VPWR VGND net27 sg13g2_antennanp
XANTENNA_40 VPWR VGND net1 sg13g2_antennanp
XFILLER_11_394 VPWR VGND sg13g2_fill_1
XFILLER_11_361 VPWR VGND sg13g2_decap_8
XFILLER_7_35 VPWR VGND sg13g2_decap_8
X_058_ N2MID[5] net59 VPWR VGND sg13g2_buf_1
XFILLER_11_191 VPWR VGND sg13g2_decap_8
XFILLER_7_140 VPWR VGND sg13g2_decap_8
XFILLER_4_346 VPWR VGND sg13g2_decap_8
XFILLER_7_195 VPWR VGND sg13g2_decap_8
XFILLER_9_427 VPWR VGND sg13g2_decap_8
XFILLER_4_14 VPWR VGND sg13g2_decap_8
XFILLER_1_305 VPWR VGND sg13g2_decap_8
XFILLER_10_415 VPWR VGND sg13g2_decap_4
XFILLER_10_404 VPWR VGND sg13g2_fill_1
XFILLER_1_102 VPWR VGND sg13g2_decap_8
XFILLER_9_224 VPWR VGND sg13g2_decap_8
XFILLER_5_485 VPWR VGND sg13g2_decap_8
XFILLER_8_290 VPWR VGND sg13g2_decap_8
XFILLER_10_256 VPWR VGND sg13g2_decap_4
XFILLER_10_223 VPWR VGND sg13g2_decap_4
XFILLER_6_249 VPWR VGND sg13g2_fill_2
X_091_ NN4END[12] net98 VPWR VGND sg13g2_buf_1
XFILLER_2_477 VPWR VGND sg13g2_decap_8
XFILLER_10_35 VPWR VGND sg13g2_decap_8
XFILLER_7_514 VPWR VGND sg13g2_decap_8
X_074_ N4END[13] net81 VPWR VGND sg13g2_buf_1
XFILLER_3_219 VPWR VGND sg13g2_decap_8
XFILLER_2_285 VPWR VGND sg13g2_decap_8
XANTENNA_30 VPWR VGND net1 sg13g2_antennanp
XANTENNA_41 VPWR VGND net27 sg13g2_antennanp
XFILLER_2_91 VPWR VGND sg13g2_decap_8
XANTENNA_52 VPWR VGND FrameData[5] sg13g2_antennanp
XFILLER_11_373 VPWR VGND sg13g2_decap_8
XFILLER_7_388 VPWR VGND sg13g2_decap_8
XFILLER_7_14 VPWR VGND sg13g2_decap_8
X_057_ N2MID[6] net58 VPWR VGND sg13g2_buf_1
XFILLER_8_119 VPWR VGND sg13g2_decap_8
XFILLER_4_325 VPWR VGND sg13g2_decap_8
XFILLER_9_406 VPWR VGND sg13g2_decap_8
XFILLER_1_339 VPWR VGND sg13g2_decap_4
XFILLER_4_199 VPWR VGND sg13g2_decap_8
XFILLER_4_144 VPWR VGND sg13g2_fill_2
XFILLER_4_133 VPWR VGND sg13g2_decap_8
XFILLER_1_158 VPWR VGND sg13g2_decap_8
XFILLER_1_114 VPWR VGND sg13g2_decap_8
XFILLER_9_258 VPWR VGND sg13g2_decap_8
XFILLER_9_203 VPWR VGND sg13g2_decap_8
XFILLER_5_464 VPWR VGND sg13g2_decap_8
XFILLER_5_91 VPWR VGND sg13g2_decap_8
XFILLER_10_246 VPWR VGND sg13g2_decap_4
XFILLER_6_228 VPWR VGND sg13g2_decap_8
XFILLER_6_217 VPWR VGND sg13g2_decap_8
XFILLER_1_49 VPWR VGND sg13g2_decap_8
X_090_ NN4END[13] net97 VPWR VGND sg13g2_buf_1
XFILLER_2_456 VPWR VGND sg13g2_decap_8
XFILLER_5_261 VPWR VGND sg13g2_decap_8
XFILLER_10_14 VPWR VGND sg13g2_decap_8
XFILLER_4_0 VPWR VGND sg13g2_decap_8
X_073_ N4END[14] net80 VPWR VGND sg13g2_buf_1
XFILLER_2_275 VPWR VGND sg13g2_decap_4
XANTENNA_20 VPWR VGND net22 sg13g2_antennanp
XANTENNA_53 VPWR VGND FrameData[6] sg13g2_antennanp
XFILLER_4_507 VPWR VGND sg13g2_decap_8
XANTENNA_31 VPWR VGND net27 sg13g2_antennanp
XFILLER_2_70 VPWR VGND sg13g2_decap_8
XANTENNA_42 VPWR VGND FrameData[5] sg13g2_antennanp
XFILLER_7_367 VPWR VGND sg13g2_decap_8
XFILLER_7_334 VPWR VGND sg13g2_decap_8
XFILLER_7_301 VPWR VGND sg13g2_fill_1
X_056_ N2MID[7] net57 VPWR VGND sg13g2_buf_1
XFILLER_4_304 VPWR VGND sg13g2_decap_8
XFILLER_11_160 VPWR VGND sg13g2_fill_1
X_039_ FrameStrobe[7] net50 VPWR VGND sg13g2_buf_1
XFILLER_7_175 VPWR VGND sg13g2_decap_8
XFILLER_3_381 VPWR VGND sg13g2_decap_8
XFILLER_8_91 VPWR VGND sg13g2_decap_8
XFILLER_4_178 VPWR VGND sg13g2_decap_8
XFILLER_4_112 VPWR VGND sg13g2_decap_8
XFILLER_4_49 VPWR VGND sg13g2_decap_8
XFILLER_10_439 VPWR VGND sg13g2_fill_1
XFILLER_8_484 VPWR VGND sg13g2_decap_8
XFILLER_8_7 VPWR VGND sg13g2_decap_8
XFILLER_5_443 VPWR VGND sg13g2_decap_8
XFILLER_5_70 VPWR VGND sg13g2_decap_8
XFILLER_10_269 VPWR VGND sg13g2_decap_8
XFILLER_1_28 VPWR VGND sg13g2_decap_8
XFILLER_5_295 VPWR VGND sg13g2_decap_8
XFILLER_5_240 VPWR VGND sg13g2_decap_8
XFILLER_1_490 VPWR VGND sg13g2_decap_8
X_072_ N4END[15] net73 VPWR VGND sg13g2_buf_1
XFILLER_2_221 VPWR VGND sg13g2_fill_1
XFILLER_2_254 VPWR VGND sg13g2_decap_8
XANTENNA_54 VPWR VGND FrameData[7] sg13g2_antennanp
XANTENNA_43 VPWR VGND FrameData[6] sg13g2_antennanp
XANTENNA_21 VPWR VGND net27 sg13g2_antennanp
XANTENNA_32 VPWR VGND FrameData[5] sg13g2_antennanp
XANTENNA_10 VPWR VGND FrameData[5] sg13g2_antennanp
XFILLER_11_342 VPWR VGND sg13g2_fill_1
XFILLER_7_313 VPWR VGND sg13g2_decap_8
XFILLER_7_49 VPWR VGND sg13g2_decap_8
X_055_ N1END[0] net56 VPWR VGND sg13g2_buf_1
XFILLER_6_390 VPWR VGND sg13g2_decap_8
XFILLER_11_172 VPWR VGND sg13g2_decap_8
X_038_ FrameStrobe[6] net49 VPWR VGND sg13g2_buf_1
XFILLER_7_154 VPWR VGND sg13g2_decap_8
XFILLER_3_360 VPWR VGND sg13g2_decap_8
XFILLER_8_70 VPWR VGND sg13g2_decap_8
XFILLER_1_319 VPWR VGND sg13g2_decap_8
XFILLER_4_157 VPWR VGND sg13g2_decap_8
XFILLER_4_28 VPWR VGND sg13g2_decap_8
XFILLER_8_463 VPWR VGND sg13g2_decap_8
XFILLER_10_429 VPWR VGND sg13g2_fill_2
XFILLER_9_238 VPWR VGND sg13g2_decap_8
XFILLER_1_138 VPWR VGND sg13g2_fill_2
XFILLER_5_499 VPWR VGND sg13g2_decap_8
XFILLER_5_422 VPWR VGND sg13g2_decap_8
XFILLER_0_182 VPWR VGND sg13g2_decap_8
XFILLER_2_403 VPWR VGND sg13g2_decap_8
XFILLER_10_49 VPWR VGND sg13g2_decap_8
X_071_ N2END[0] net72 VPWR VGND sg13g2_buf_1
XFILLER_2_233 VPWR VGND sg13g2_decap_8
XFILLER_11_321 VPWR VGND sg13g2_decap_8
XANTENNA_44 VPWR VGND FrameData[7] sg13g2_antennanp
XANTENNA_33 VPWR VGND FrameData[6] sg13g2_antennanp
XANTENNA_11 VPWR VGND FrameData[6] sg13g2_antennanp
XANTENNA_55 VPWR VGND net1 sg13g2_antennanp
XANTENNA_22 VPWR VGND FrameData[5] sg13g2_antennanp
XFILLER_11_387 VPWR VGND sg13g2_decap_8
XFILLER_11_354 VPWR VGND sg13g2_decap_8
XFILLER_7_28 VPWR VGND sg13g2_decap_8
X_054_ N1END[1] net55 VPWR VGND sg13g2_buf_1
XFILLER_4_339 VPWR VGND sg13g2_decap_8
X_037_ FrameStrobe[5] net48 VPWR VGND sg13g2_buf_1
XFILLER_7_188 VPWR VGND sg13g2_decap_8
XFILLER_7_133 VPWR VGND sg13g2_decap_8
XFILLER_0_523 VPWR VGND sg13g2_fill_1
XFILLER_3_394 VPWR VGND sg13g2_decap_8
XFILLER_8_442 VPWR VGND sg13g2_decap_8
XFILLER_3_191 VPWR VGND sg13g2_decap_8
XFILLER_10_419 VPWR VGND sg13g2_fill_2
XFILLER_1_128 VPWR VGND sg13g2_decap_4
XFILLER_9_217 VPWR VGND sg13g2_decap_8
XFILLER_5_478 VPWR VGND sg13g2_decap_8
XFILLER_5_401 VPWR VGND sg13g2_decap_8
XFILLER_0_161 VPWR VGND sg13g2_decap_8
XFILLER_10_227 VPWR VGND sg13g2_fill_2
XFILLER_10_216 VPWR VGND sg13g2_decap_8
XFILLER_8_283 VPWR VGND sg13g2_decap_8
XFILLER_5_231 VPWR VGND sg13g2_decap_4
XFILLER_10_28 VPWR VGND sg13g2_decap_8
XFILLER_5_275 VPWR VGND sg13g2_fill_2
XFILLER_11_503 VPWR VGND sg13g2_fill_1
XFILLER_7_507 VPWR VGND sg13g2_decap_8
X_070_ N2END[1] net71 VPWR VGND sg13g2_buf_1
XFILLER_2_84 VPWR VGND sg13g2_decap_8
XANTENNA_12 VPWR VGND FrameData[7] sg13g2_antennanp
XANTENNA_34 VPWR VGND FrameData[7] sg13g2_antennanp
XANTENNA_23 VPWR VGND FrameData[6] sg13g2_antennanp
XANTENNA_45 VPWR VGND net1 sg13g2_antennanp
XANTENNA_56 VPWR VGND net27 sg13g2_antennanp
XFILLER_11_399 VPWR VGND sg13g2_decap_8
XFILLER_11_82 VPWR VGND sg13g2_fill_1
XFILLER_7_348 VPWR VGND sg13g2_decap_4
X_053_ N1END[2] net54 VPWR VGND sg13g2_buf_1
XFILLER_2_0 VPWR VGND sg13g2_decap_8
XFILLER_7_112 VPWR VGND sg13g2_decap_8
XFILLER_4_318 VPWR VGND sg13g2_decap_8
X_036_ FrameStrobe[4] net47 VPWR VGND sg13g2_buf_1
XFILLER_4_126 VPWR VGND sg13g2_decap_8
XFILLER_8_498 VPWR VGND sg13g2_decap_8
XFILLER_8_421 VPWR VGND sg13g2_decap_8
X_019_ FrameData[19] net11 VPWR VGND sg13g2_buf_1
XFILLER_3_181 VPWR VGND sg13g2_decap_4
XFILLER_10_409 VPWR VGND sg13g2_fill_2
XFILLER_5_457 VPWR VGND sg13g2_decap_8
XFILLER_0_140 VPWR VGND sg13g2_decap_8
XFILLER_8_262 VPWR VGND sg13g2_decap_8
XFILLER_5_84 VPWR VGND sg13g2_decap_8
XFILLER_10_239 VPWR VGND sg13g2_decap_8
XFILLER_6_7 VPWR VGND sg13g2_decap_8
XFILLER_5_254 VPWR VGND sg13g2_decap_8
XFILLER_5_210 VPWR VGND sg13g2_decap_8
XFILLER_2_202 VPWR VGND sg13g2_decap_8
XFILLER_2_268 VPWR VGND sg13g2_decap_8
XFILLER_2_279 VPWR VGND sg13g2_fill_2
XANTENNA_24 VPWR VGND FrameData[7] sg13g2_antennanp
XANTENNA_46 VPWR VGND net27 sg13g2_antennanp
XANTENNA_35 VPWR VGND net1 sg13g2_antennanp
XANTENNA_13 VPWR VGND net1 sg13g2_antennanp
XFILLER_2_63 VPWR VGND sg13g2_decap_8
XFILLER_11_94 VPWR VGND sg13g2_decap_8
XFILLER_11_61 VPWR VGND sg13g2_decap_8
XFILLER_7_327 VPWR VGND sg13g2_decap_8
X_052_ N1END[3] net53 VPWR VGND sg13g2_buf_1
XFILLER_11_186 VPWR VGND sg13g2_fill_1
XFILLER_11_153 VPWR VGND sg13g2_decap_8
XFILLER_11_120 VPWR VGND sg13g2_decap_8
X_104_ UserCLK net105 VPWR VGND sg13g2_buf_1
X_035_ FrameStrobe[3] net46 VPWR VGND sg13g2_buf_1
XFILLER_7_168 VPWR VGND sg13g2_decap_8
XFILLER_3_374 VPWR VGND sg13g2_decap_8
XFILLER_8_84 VPWR VGND sg13g2_decap_8
XFILLER_4_105 VPWR VGND sg13g2_decap_8
XFILLER_8_477 VPWR VGND sg13g2_decap_8
XFILLER_8_400 VPWR VGND sg13g2_decap_8
X_018_ FrameData[18] net10 VPWR VGND sg13g2_buf_1
XFILLER_5_436 VPWR VGND sg13g2_decap_8
XFILLER_0_196 VPWR VGND sg13g2_decap_8
XFILLER_10_0 VPWR VGND sg13g2_decap_8
XFILLER_8_241 VPWR VGND sg13g2_decap_8
XFILLER_5_63 VPWR VGND sg13g2_decap_8
XFILLER_2_417 VPWR VGND sg13g2_decap_4
XFILLER_5_288 VPWR VGND sg13g2_decap_8
XFILLER_1_483 VPWR VGND sg13g2_decap_8
XFILLER_2_247 VPWR VGND sg13g2_decap_8
XANTENNA_14 VPWR VGND net22 sg13g2_antennanp
XFILLER_1_280 VPWR VGND sg13g2_fill_2
XFILLER_1_291 VPWR VGND sg13g2_decap_8
XFILLER_2_42 VPWR VGND sg13g2_decap_8
XANTENNA_47 VPWR VGND FrameData[5] sg13g2_antennanp
XANTENNA_25 VPWR VGND net1 sg13g2_antennanp
XANTENNA_36 VPWR VGND net27 sg13g2_antennanp
XFILLER_11_368 VPWR VGND sg13g2_fill_1
XFILLER_11_335 VPWR VGND sg13g2_decap_8
XFILLER_11_302 VPWR VGND sg13g2_decap_8
X_051_ FrameStrobe[19] net43 VPWR VGND sg13g2_buf_1
XFILLER_7_306 VPWR VGND sg13g2_decap_8
XFILLER_10_390 VPWR VGND sg13g2_decap_8
XFILLER_11_198 VPWR VGND sg13g2_decap_8
XFILLER_11_165 VPWR VGND sg13g2_decap_8
X_034_ FrameStrobe[2] net45 VPWR VGND sg13g2_buf_1
XFILLER_7_147 VPWR VGND sg13g2_decap_8
XFILLER_3_353 VPWR VGND sg13g2_decap_8
X_103_ NN4END[0] net95 VPWR VGND sg13g2_buf_1
XFILLER_8_63 VPWR VGND sg13g2_decap_8
XFILLER_8_456 VPWR VGND sg13g2_decap_8
X_017_ FrameData[17] net9 VPWR VGND sg13g2_buf_1
XFILLER_5_415 VPWR VGND sg13g2_decap_8
XFILLER_1_109 VPWR VGND sg13g2_fill_1
XFILLER_8_297 VPWR VGND sg13g2_decap_8
XFILLER_5_42 VPWR VGND sg13g2_decap_8
XFILLER_0_175 VPWR VGND sg13g2_decap_8
XFILLER_1_462 VPWR VGND sg13g2_decap_8
XFILLER_2_226 VPWR VGND sg13g2_decap_8
XANTENNA_48 VPWR VGND FrameData[6] sg13g2_antennanp
XANTENNA_26 VPWR VGND net27 sg13g2_antennanp
XFILLER_2_21 VPWR VGND sg13g2_decap_8
XFILLER_2_98 VPWR VGND sg13g2_decap_8
XANTENNA_37 VPWR VGND FrameData[5] sg13g2_antennanp
XANTENNA_15 VPWR VGND net27 sg13g2_antennanp
XFILLER_11_347 VPWR VGND sg13g2_decap_8
XFILLER_11_30 VPWR VGND sg13g2_fill_1
X_050_ FrameStrobe[18] net42 VPWR VGND sg13g2_buf_1
XFILLER_9_392 VPWR VGND sg13g2_decap_8
Xoutput100 net100 SS4BEG[5] VPWR VGND sg13g2_buf_1
XFILLER_6_351 VPWR VGND sg13g2_decap_4
XFILLER_3_513 VPWR VGND sg13g2_fill_2
X_033_ FrameStrobe[1] net44 VPWR VGND sg13g2_buf_1
XFILLER_7_126 VPWR VGND sg13g2_decap_8
XFILLER_3_332 VPWR VGND sg13g2_decap_8
XFILLER_0_0 VPWR VGND sg13g2_decap_8
X_102_ NN4END[1] net94 VPWR VGND sg13g2_buf_1
XFILLER_8_42 VPWR VGND sg13g2_decap_8
XFILLER_8_435 VPWR VGND sg13g2_decap_8
X_016_ FrameData[16] net8 VPWR VGND sg13g2_buf_1
XFILLER_3_162 VPWR VGND sg13g2_fill_1
XFILLER_8_276 VPWR VGND sg13g2_fill_2
XFILLER_8_210 VPWR VGND sg13g2_decap_8
XFILLER_5_21 VPWR VGND sg13g2_decap_8
XFILLER_0_154 VPWR VGND sg13g2_decap_8
XFILLER_10_209 VPWR VGND sg13g2_decap_8
XFILLER_5_98 VPWR VGND sg13g2_decap_8
XFILLER_4_493 VPWR VGND sg13g2_decap_8
XFILLER_5_268 VPWR VGND sg13g2_decap_8
XFILLER_5_235 VPWR VGND sg13g2_fill_1
XFILLER_5_224 VPWR VGND sg13g2_decap_8
XFILLER_1_441 VPWR VGND sg13g2_decap_8
XFILLER_4_7 VPWR VGND sg13g2_decap_8
XFILLER_1_282 VPWR VGND sg13g2_fill_1
XFILLER_2_77 VPWR VGND sg13g2_decap_8
XFILLER_9_371 VPWR VGND sg13g2_decap_8
XANTENNA_49 VPWR VGND FrameData[7] sg13g2_antennanp
XANTENNA_38 VPWR VGND FrameData[6] sg13g2_antennanp
Xoutput101 net101 SS4BEG[6] VPWR VGND sg13g2_buf_1
XANTENNA_27 VPWR VGND FrameData[5] sg13g2_antennanp
XANTENNA_16 VPWR VGND FrameData[5] sg13g2_antennanp
XFILLER_11_75 VPWR VGND sg13g2_decap_8
XFILLER_11_42 VPWR VGND sg13g2_decap_8
XFILLER_6_385 VPWR VGND sg13g2_fill_1
XFILLER_6_330 VPWR VGND sg13g2_decap_8
XFILLER_11_134 VPWR VGND sg13g2_fill_1
XFILLER_11_101 VPWR VGND sg13g2_decap_8
X_032_ FrameStrobe[0] net33 VPWR VGND sg13g2_buf_1
XFILLER_7_105 VPWR VGND sg13g2_decap_8
XFILLER_3_388 VPWR VGND sg13g2_fill_2
X_101_ NN4END[2] net93 VPWR VGND sg13g2_buf_1
XFILLER_3_311 VPWR VGND sg13g2_decap_8
XFILLER_8_98 VPWR VGND sg13g2_decap_8
XFILLER_8_21 VPWR VGND sg13g2_decap_8
XFILLER_6_182 VPWR VGND sg13g2_decap_8
XFILLER_4_119 VPWR VGND sg13g2_decap_8
XFILLER_8_414 VPWR VGND sg13g2_decap_8
X_015_ FrameData[15] net7 VPWR VGND sg13g2_buf_1
XFILLER_3_152 VPWR VGND sg13g2_decap_4
XFILLER_3_174 VPWR VGND sg13g2_decap_8
XFILLER_3_185 VPWR VGND sg13g2_fill_2
XFILLER_0_133 VPWR VGND sg13g2_decap_8
XFILLER_8_255 VPWR VGND sg13g2_decap_8
XFILLER_5_77 VPWR VGND sg13g2_decap_8
XFILLER_4_472 VPWR VGND sg13g2_decap_8
XFILLER_5_247 VPWR VGND sg13g2_decap_8
XFILLER_5_203 VPWR VGND sg13g2_decap_8
XFILLER_1_420 VPWR VGND sg13g2_decap_8
XFILLER_1_497 VPWR VGND sg13g2_fill_1
XFILLER_2_217 VPWR VGND sg13g2_decap_4
XFILLER_2_56 VPWR VGND sg13g2_decap_8
XANTENNA_39 VPWR VGND FrameData[7] sg13g2_antennanp
XANTENNA_17 VPWR VGND FrameData[6] sg13g2_antennanp
XANTENNA_28 VPWR VGND FrameData[6] sg13g2_antennanp
Xoutput102 net102 SS4BEG[7] VPWR VGND sg13g2_buf_1
XFILLER_11_316 VPWR VGND sg13g2_fill_1
XFILLER_11_87 VPWR VGND sg13g2_decap_8
XFILLER_3_515 VPWR VGND sg13g2_fill_1
XFILLER_6_397 VPWR VGND sg13g2_decap_8
XFILLER_11_179 VPWR VGND sg13g2_decap_8
XFILLER_11_146 VPWR VGND sg13g2_decap_8
XFILLER_11_113 VPWR VGND sg13g2_decap_8
X_031_ FrameData[31] net25 VPWR VGND sg13g2_buf_1
X_100_ NN4END[3] net92 VPWR VGND sg13g2_buf_1
XFILLER_8_77 VPWR VGND sg13g2_decap_8
XFILLER_6_161 VPWR VGND sg13g2_decap_8
XFILLER_3_367 VPWR VGND sg13g2_decap_8
X_014_ FrameData[14] net6 VPWR VGND sg13g2_buf_1
XFILLER_3_131 VPWR VGND sg13g2_decap_8
XFILLER_5_429 VPWR VGND sg13g2_decap_8
XFILLER_0_189 VPWR VGND sg13g2_decap_8
XFILLER_0_112 VPWR VGND sg13g2_decap_8
XFILLER_8_278 VPWR VGND sg13g2_fill_1
XFILLER_8_234 VPWR VGND sg13g2_decap_8
XFILLER_5_56 VPWR VGND sg13g2_decap_8
XFILLER_4_451 VPWR VGND sg13g2_decap_8
XFILLER_1_476 VPWR VGND sg13g2_decap_8
XFILLER_6_502 VPWR VGND sg13g2_decap_8
XFILLER_1_251 VPWR VGND sg13g2_fill_2
XANTENNA_18 VPWR VGND FrameData[7] sg13g2_antennanp
XANTENNA_29 VPWR VGND FrameData[7] sg13g2_antennanp
XFILLER_1_273 VPWR VGND sg13g2_decap_8
Xoutput103 net103 SS4BEG[8] VPWR VGND sg13g2_buf_1
XFILLER_2_35 VPWR VGND sg13g2_decap_8
XFILLER_11_328 VPWR VGND sg13g2_decap_8
XFILLER_10_383 VPWR VGND sg13g2_decap_8
X_030_ FrameData[30] net24 VPWR VGND sg13g2_buf_1
XFILLER_8_56 VPWR VGND sg13g2_decap_8
XFILLER_3_346 VPWR VGND sg13g2_decap_8
XFILLER_10_191 VPWR VGND sg13g2_decap_8
XFILLER_6_140 VPWR VGND sg13g2_decap_8
X_013_ FrameData[13] net5 VPWR VGND sg13g2_buf_1
XFILLER_8_449 VPWR VGND sg13g2_decap_8
XFILLER_7_493 VPWR VGND sg13g2_decap_8
XFILLER_3_198 VPWR VGND sg13g2_decap_8
XFILLER_5_408 VPWR VGND sg13g2_decap_8
XFILLER_0_168 VPWR VGND sg13g2_decap_8
XFILLER_8_224 VPWR VGND sg13g2_decap_4
XFILLER_5_35 VPWR VGND sg13g2_decap_8
XFILLER_4_430 VPWR VGND sg13g2_decap_8
XFILLER_1_455 VPWR VGND sg13g2_decap_8
XFILLER_9_522 VPWR VGND sg13g2_fill_1
XFILLER_9_511 VPWR VGND sg13g2_decap_8
XFILLER_4_282 VPWR VGND sg13g2_decap_8
XFILLER_9_385 VPWR VGND sg13g2_decap_8
XFILLER_9_0 VPWR VGND sg13g2_decap_8
Xoutput104 net104 SS4BEG[9] VPWR VGND sg13g2_buf_1
XANTENNA_19 VPWR VGND net1 sg13g2_antennanp
XFILLER_2_14 VPWR VGND sg13g2_decap_8
XFILLER_11_56 VPWR VGND sg13g2_fill_1
XFILLER_11_23 VPWR VGND sg13g2_decap_8
XFILLER_3_506 VPWR VGND sg13g2_decap_8
XFILLER_2_7 VPWR VGND sg13g2_decap_8
XFILLER_10_362 VPWR VGND sg13g2_decap_8
XFILLER_6_355 VPWR VGND sg13g2_fill_2
XFILLER_6_344 VPWR VGND sg13g2_decap_8
XFILLER_9_182 VPWR VGND sg13g2_decap_8
XFILLER_7_119 VPWR VGND sg13g2_decap_8
XFILLER_3_325 VPWR VGND sg13g2_decap_8
XFILLER_10_170 VPWR VGND sg13g2_decap_8
XFILLER_8_35 VPWR VGND sg13g2_decap_8
XFILLER_6_196 VPWR VGND sg13g2_decap_8
X_089_ NN4END[14] net96 VPWR VGND sg13g2_buf_1
XFILLER_8_428 VPWR VGND sg13g2_decap_8
XFILLER_7_472 VPWR VGND sg13g2_decap_8
X_012_ FrameData[12] net4 VPWR VGND sg13g2_buf_1
XFILLER_0_91 VPWR VGND sg13g2_decap_8
XFILLER_8_269 VPWR VGND sg13g2_decap_8
XFILLER_8_203 VPWR VGND sg13g2_decap_8
XFILLER_5_14 VPWR VGND sg13g2_decap_8
XFILLER_4_486 VPWR VGND sg13g2_decap_8
XFILLER_0_147 VPWR VGND sg13g2_decap_8
XFILLER_5_217 VPWR VGND sg13g2_decap_8
XFILLER_1_401 VPWR VGND sg13g2_fill_1
XFILLER_1_434 VPWR VGND sg13g2_decap_8
XFILLER_4_261 VPWR VGND sg13g2_decap_8
XFILLER_10_522 VPWR VGND sg13g2_fill_1
XFILLER_9_364 VPWR VGND sg13g2_decap_8
XFILLER_1_253 VPWR VGND sg13g2_fill_1
XFILLER_1_242 VPWR VGND sg13g2_fill_1
XFILLER_1_231 VPWR VGND sg13g2_fill_1
XFILLER_11_35 VPWR VGND sg13g2_decap_8
Xoutput105 net105 UserCLKo VPWR VGND sg13g2_buf_1
XFILLER_11_68 VPWR VGND sg13g2_decap_8
XFILLER_10_341 VPWR VGND sg13g2_decap_8
XFILLER_6_323 VPWR VGND sg13g2_decap_8
XFILLER_9_161 VPWR VGND sg13g2_decap_8
XFILLER_11_127 VPWR VGND sg13g2_decap_8
XFILLER_3_91 VPWR VGND sg13g2_decap_8
XFILLER_3_304 VPWR VGND sg13g2_decap_8
XFILLER_8_14 VPWR VGND sg13g2_decap_8
XFILLER_6_175 VPWR VGND sg13g2_decap_8
X_088_ NN4END[15] net89 VPWR VGND sg13g2_buf_1
XFILLER_8_407 VPWR VGND sg13g2_decap_8
X_011_ FrameData[11] net3 VPWR VGND sg13g2_buf_1
XFILLER_3_112 VPWR VGND sg13g2_decap_8
XFILLER_3_145 VPWR VGND sg13g2_decap_8
XFILLER_3_156 VPWR VGND sg13g2_fill_2
XFILLER_3_167 VPWR VGND sg13g2_decap_8
XFILLER_11_491 VPWR VGND sg13g2_decap_8
XFILLER_7_451 VPWR VGND sg13g2_decap_8
XFILLER_0_70 VPWR VGND sg13g2_decap_8
XFILLER_8_248 VPWR VGND sg13g2_decap_8
XFILLER_0_126 VPWR VGND sg13g2_decap_8
XFILLER_10_7 VPWR VGND sg13g2_decap_8
XFILLER_4_465 VPWR VGND sg13g2_decap_8
XFILLER_1_413 VPWR VGND sg13g2_decap_8
XFILLER_6_91 VPWR VGND sg13g2_decap_8
XFILLER_6_516 VPWR VGND sg13g2_decap_8
XFILLER_1_265 VPWR VGND sg13g2_decap_4
XFILLER_1_298 VPWR VGND sg13g2_decap_8
XFILLER_2_49 VPWR VGND sg13g2_decap_8
XFILLER_11_309 VPWR VGND sg13g2_decap_8
XFILLER_10_320 VPWR VGND sg13g2_decap_8
XFILLER_6_302 VPWR VGND sg13g2_decap_8
XFILLER_10_397 VPWR VGND sg13g2_decap_8
XFILLER_9_140 VPWR VGND sg13g2_decap_8
XFILLER_11_139 VPWR VGND sg13g2_decap_8
XFILLER_3_70 VPWR VGND sg13g2_decap_8
XFILLER_6_154 VPWR VGND sg13g2_decap_8
X_087_ N4END[0] net79 VPWR VGND sg13g2_buf_1
XFILLER_2_382 VPWR VGND sg13g2_decap_8
X_010_ FrameData[10] net2 VPWR VGND sg13g2_buf_1
XFILLER_7_430 VPWR VGND sg13g2_decap_8
XFILLER_9_91 VPWR VGND sg13g2_decap_8
XFILLER_0_105 VPWR VGND sg13g2_decap_8
XFILLER_5_49 VPWR VGND sg13g2_decap_8
XFILLER_4_444 VPWR VGND sg13g2_decap_8
XFILLER_7_293 VPWR VGND sg13g2_decap_4
XFILLER_4_296 VPWR VGND sg13g2_decap_4
XFILLER_1_469 VPWR VGND sg13g2_decap_8
XFILLER_6_70 VPWR VGND sg13g2_decap_8
XFILLER_2_28 VPWR VGND sg13g2_decap_8
XFILLER_9_399 VPWR VGND sg13g2_decap_8
XFILLER_10_376 VPWR VGND sg13g2_decap_8
XFILLER_7_0 VPWR VGND sg13g2_decap_8
XFILLER_9_196 VPWR VGND sg13g2_decap_8
XFILLER_5_380 VPWR VGND sg13g2_decap_8
XFILLER_10_184 VPWR VGND sg13g2_decap_8
XFILLER_10_140 VPWR VGND sg13g2_decap_8
XFILLER_8_49 VPWR VGND sg13g2_decap_8
XFILLER_6_133 VPWR VGND sg13g2_decap_8
XFILLER_3_339 VPWR VGND sg13g2_decap_8
XFILLER_0_7 VPWR VGND sg13g2_decap_8
X_086_ N4END[1] net78 VPWR VGND sg13g2_buf_1
XFILLER_2_350 VPWR VGND sg13g2_fill_2
XFILLER_7_486 VPWR VGND sg13g2_decap_8
X_069_ N2END[2] net70 VPWR VGND sg13g2_buf_1
XFILLER_9_70 VPWR VGND sg13g2_decap_8
XFILLER_8_228 VPWR VGND sg13g2_fill_2
XFILLER_8_217 VPWR VGND sg13g2_decap_8
XFILLER_5_28 VPWR VGND sg13g2_decap_8
XFILLER_4_423 VPWR VGND sg13g2_decap_8
XFILLER_11_290 VPWR VGND sg13g2_fill_1
XFILLER_7_272 VPWR VGND sg13g2_decap_8
XFILLER_9_504 VPWR VGND sg13g2_decap_8
XFILLER_1_448 VPWR VGND sg13g2_decap_8
XFILLER_4_275 VPWR VGND sg13g2_decap_8
XFILLER_4_220 VPWR VGND sg13g2_decap_8
XFILLER_1_223 VPWR VGND sg13g2_decap_4
XFILLER_9_378 VPWR VGND sg13g2_decap_8
XFILLER_9_312 VPWR VGND sg13g2_decap_8
Xoutput90 net90 SS4BEG[10] VPWR VGND sg13g2_buf_1
XFILLER_11_49 VPWR VGND sg13g2_decap_8
XFILLER_11_16 VPWR VGND sg13g2_decap_8
XFILLER_10_355 VPWR VGND sg13g2_decap_8
XFILLER_6_337 VPWR VGND sg13g2_decap_8
XFILLER_11_108 VPWR VGND sg13g2_fill_1
XFILLER_9_175 VPWR VGND sg13g2_decap_8
XFILLER_8_28 VPWR VGND sg13g2_decap_8
XFILLER_3_318 VPWR VGND sg13g2_decap_8
XFILLER_10_163 VPWR VGND sg13g2_decap_8
XFILLER_6_189 VPWR VGND sg13g2_decap_8
XFILLER_6_112 VPWR VGND sg13g2_decap_8
XFILLER_2_362 VPWR VGND sg13g2_fill_1
X_085_ N4END[2] net77 VPWR VGND sg13g2_buf_1
XFILLER_3_126 VPWR VGND sg13g2_fill_1
XFILLER_11_472 VPWR VGND sg13g2_fill_1
XFILLER_7_465 VPWR VGND sg13g2_decap_8
XFILLER_2_170 VPWR VGND sg13g2_decap_8
X_068_ N2END[3] net69 VPWR VGND sg13g2_buf_1
XFILLER_0_84 VPWR VGND sg13g2_decap_8
XFILLER_4_479 VPWR VGND sg13g2_decap_8
XFILLER_4_402 VPWR VGND sg13g2_decap_8
XFILLER_7_251 VPWR VGND sg13g2_decap_8
XFILLER_1_427 VPWR VGND sg13g2_decap_8
XFILLER_4_254 VPWR VGND sg13g2_decap_8
XFILLER_4_243 VPWR VGND sg13g2_fill_2
XFILLER_0_482 VPWR VGND sg13g2_decap_8
Xoutput1 net1 FrameData_O[0] VPWR VGND sg13g2_buf_1
Xoutput80 net80 S4BEG[1] VPWR VGND sg13g2_buf_1
Xoutput91 net91 SS4BEG[11] VPWR VGND sg13g2_buf_1
XFILLER_10_334 VPWR VGND sg13g2_decap_8
XFILLER_10_301 VPWR VGND sg13g2_fill_1
XFILLER_6_316 VPWR VGND sg13g2_decap_8
XFILLER_9_154 VPWR VGND sg13g2_decap_8
XFILLER_3_84 VPWR VGND sg13g2_decap_8
XFILLER_6_168 VPWR VGND sg13g2_decap_8
X_084_ N4END[3] net76 VPWR VGND sg13g2_buf_1
XFILLER_2_374 VPWR VGND sg13g2_decap_4
XFILLER_2_396 VPWR VGND sg13g2_decap_8
XFILLER_11_484 VPWR VGND sg13g2_decap_8
XFILLER_11_451 VPWR VGND sg13g2_decap_8
XFILLER_7_444 VPWR VGND sg13g2_decap_8
XFILLER_3_105 VPWR VGND sg13g2_decap_8
XFILLER_3_138 VPWR VGND sg13g2_decap_8
XFILLER_0_63 VPWR VGND sg13g2_decap_8
X_067_ N2END[4] net68 VPWR VGND sg13g2_buf_1
XFILLER_4_458 VPWR VGND sg13g2_decap_8
XFILLER_0_119 VPWR VGND sg13g2_decap_8
XFILLER_7_230 VPWR VGND sg13g2_fill_2
XFILLER_1_406 VPWR VGND sg13g2_decap_8
XFILLER_0_461 VPWR VGND sg13g2_decap_8
XFILLER_10_505 VPWR VGND sg13g2_decap_4
XFILLER_6_84 VPWR VGND sg13g2_decap_8
XFILLER_6_509 VPWR VGND sg13g2_decap_8
XFILLER_1_258 VPWR VGND sg13g2_decap_8
XFILLER_1_236 VPWR VGND sg13g2_fill_2
XFILLER_5_520 VPWR VGND sg13g2_fill_2
Xoutput2 net2 FrameData_O[10] VPWR VGND sg13g2_buf_1
Xoutput70 net70 S2BEGb[5] VPWR VGND sg13g2_buf_1
Xoutput81 net81 S4BEG[2] VPWR VGND sg13g2_buf_1
Xoutput92 net92 SS4BEG[12] VPWR VGND sg13g2_buf_1
XFILLER_10_313 VPWR VGND sg13g2_decap_8
XFILLER_9_133 VPWR VGND sg13g2_decap_8
XFILLER_5_394 VPWR VGND sg13g2_decap_8
XFILLER_3_63 VPWR VGND sg13g2_decap_8
XFILLER_10_198 VPWR VGND sg13g2_decap_8
XFILLER_6_147 VPWR VGND sg13g2_decap_8
XFILLER_5_0 VPWR VGND sg13g2_decap_8
X_083_ N4END[4] net75 VPWR VGND sg13g2_buf_1
XFILLER_9_84 VPWR VGND sg13g2_decap_8
XFILLER_7_423 VPWR VGND sg13g2_decap_8
XFILLER_0_42 VPWR VGND sg13g2_decap_8
X_066_ N2END[5] net67 VPWR VGND sg13g2_buf_1
XFILLER_4_437 VPWR VGND sg13g2_decap_8
X_049_ FrameStrobe[17] net41 VPWR VGND sg13g2_buf_1
XFILLER_7_286 VPWR VGND sg13g2_decap_8
XFILLER_3_492 VPWR VGND sg13g2_decap_8
XFILLER_9_518 VPWR VGND sg13g2_decap_4
XFILLER_4_289 VPWR VGND sg13g2_decap_8
XFILLER_4_245 VPWR VGND sg13g2_fill_1
XFILLER_4_234 VPWR VGND sg13g2_decap_4
XFILLER_0_440 VPWR VGND sg13g2_decap_8
XANTENNA_1 VPWR VGND FrameData[10] sg13g2_antennanp
XFILLER_6_63 VPWR VGND sg13g2_decap_8
XFILLER_9_7 VPWR VGND sg13g2_decap_8
XFILLER_9_326 VPWR VGND sg13g2_decap_8
Xoutput3 net3 FrameData_O[11] VPWR VGND sg13g2_buf_1
Xoutput60 net60 S2BEG[3] VPWR VGND sg13g2_buf_1
Xoutput71 net71 S2BEGb[6] VPWR VGND sg13g2_buf_1
Xoutput82 net82 S4BEG[3] VPWR VGND sg13g2_buf_1
Xoutput93 net93 SS4BEG[13] VPWR VGND sg13g2_buf_1
XFILLER_10_369 VPWR VGND sg13g2_decap_8
XFILLER_9_189 VPWR VGND sg13g2_decap_8
XFILLER_9_112 VPWR VGND sg13g2_decap_8
XFILLER_5_373 VPWR VGND sg13g2_decap_8
XFILLER_5_351 VPWR VGND sg13g2_decap_8
XFILLER_3_42 VPWR VGND sg13g2_decap_8
XFILLER_10_177 VPWR VGND sg13g2_fill_2
XFILLER_6_126 VPWR VGND sg13g2_decap_8
X_082_ N4END[5] net74 VPWR VGND sg13g2_buf_1
XFILLER_2_321 VPWR VGND sg13g2_decap_4
XFILLER_2_343 VPWR VGND sg13g2_decap_8
XFILLER_11_420 VPWR VGND sg13g2_fill_1
XFILLER_7_479 VPWR VGND sg13g2_decap_8
XFILLER_7_402 VPWR VGND sg13g2_decap_8
X_065_ N2END[6] net66 VPWR VGND sg13g2_buf_1
XFILLER_0_98 VPWR VGND sg13g2_decap_8
XFILLER_0_21 VPWR VGND sg13g2_decap_8
XFILLER_2_151 VPWR VGND sg13g2_decap_8
XFILLER_2_184 VPWR VGND sg13g2_decap_8
XFILLER_2_195 VPWR VGND sg13g2_decap_8
XFILLER_9_63 VPWR VGND sg13g2_decap_8
XFILLER_11_283 VPWR VGND sg13g2_decap_8
XFILLER_11_250 VPWR VGND sg13g2_decap_8
XFILLER_7_265 VPWR VGND sg13g2_decap_8
XFILLER_7_232 VPWR VGND sg13g2_fill_1
XFILLER_4_416 VPWR VGND sg13g2_decap_8
X_048_ FrameStrobe[16] net40 VPWR VGND sg13g2_buf_1
XFILLER_3_471 VPWR VGND sg13g2_decap_8
XFILLER_4_268 VPWR VGND sg13g2_decap_8
XFILLER_4_213 VPWR VGND sg13g2_decap_8
XFILLER_6_42 VPWR VGND sg13g2_decap_8
XANTENNA_2 VPWR VGND FrameData[5] sg13g2_antennanp
XFILLER_3_290 VPWR VGND sg13g2_decap_8
XFILLER_1_216 VPWR VGND sg13g2_decap_8
Xoutput50 net50 FrameStrobe_O[7] VPWR VGND sg13g2_buf_1
XFILLER_9_305 VPWR VGND sg13g2_decap_8
XFILLER_5_522 VPWR VGND sg13g2_fill_1
Xoutput4 net4 FrameData_O[12] VPWR VGND sg13g2_buf_1
Xoutput61 net61 S2BEG[4] VPWR VGND sg13g2_buf_1
Xoutput72 net72 S2BEGb[7] VPWR VGND sg13g2_buf_1
Xoutput83 net83 S4BEG[4] VPWR VGND sg13g2_buf_1
Xoutput94 net94 SS4BEG[14] VPWR VGND sg13g2_buf_1
XFILLER_8_393 VPWR VGND sg13g2_decap_8
XFILLER_10_348 VPWR VGND sg13g2_decap_8
XFILLER_9_168 VPWR VGND sg13g2_decap_8
XFILLER_5_330 VPWR VGND sg13g2_decap_8
XFILLER_3_21 VPWR VGND sg13g2_decap_8
XFILLER_3_98 VPWR VGND sg13g2_decap_8
XFILLER_10_156 VPWR VGND sg13g2_decap_8
XFILLER_10_112 VPWR VGND sg13g2_decap_8
XFILLER_6_105 VPWR VGND sg13g2_decap_8
XFILLER_2_300 VPWR VGND sg13g2_decap_4
X_081_ N4END[6] net88 VPWR VGND sg13g2_buf_1
XFILLER_5_182 VPWR VGND sg13g2_decap_8
XFILLER_3_119 VPWR VGND sg13g2_decap_8
XFILLER_11_498 VPWR VGND sg13g2_fill_1
XFILLER_11_465 VPWR VGND sg13g2_decap_8
XFILLER_11_432 VPWR VGND sg13g2_decap_8
XFILLER_7_458 VPWR VGND sg13g2_decap_8
X_064_ N2END[7] net65 VPWR VGND sg13g2_buf_1
XFILLER_9_42 VPWR VGND sg13g2_decap_8
XFILLER_0_77 VPWR VGND sg13g2_decap_8
XFILLER_11_295 VPWR VGND sg13g2_decap_8
X_047_ FrameStrobe[15] net39 VPWR VGND sg13g2_buf_1
XFILLER_7_244 VPWR VGND sg13g2_decap_8
XFILLER_3_450 VPWR VGND sg13g2_decap_8
XFILLER_6_98 VPWR VGND sg13g2_decap_8
XFILLER_6_21 VPWR VGND sg13g2_decap_8
XANTENNA_3 VPWR VGND FrameData[6] sg13g2_antennanp
XFILLER_0_475 VPWR VGND sg13g2_decap_8
Xoutput40 net40 FrameStrobe_O[16] VPWR VGND sg13g2_buf_1
Xoutput51 net51 FrameStrobe_O[8] VPWR VGND sg13g2_buf_1
Xoutput5 net5 FrameData_O[13] VPWR VGND sg13g2_buf_1
Xoutput62 net62 S2BEG[5] VPWR VGND sg13g2_buf_1
Xoutput73 net73 S4BEG[0] VPWR VGND sg13g2_buf_1
Xoutput84 net84 S4BEG[5] VPWR VGND sg13g2_buf_1
Xoutput95 net95 SS4BEG[15] VPWR VGND sg13g2_buf_1
XFILLER_8_372 VPWR VGND sg13g2_decap_8
XFILLER_10_327 VPWR VGND sg13g2_decap_8
XFILLER_6_309 VPWR VGND sg13g2_decap_8
XFILLER_9_147 VPWR VGND sg13g2_decap_8
XFILLER_3_77 VPWR VGND sg13g2_decap_8
X_080_ N4END[7] net87 VPWR VGND sg13g2_buf_1
XFILLER_10_179 VPWR VGND sg13g2_fill_1
XFILLER_2_334 VPWR VGND sg13g2_decap_4
XFILLER_2_356 VPWR VGND sg13g2_fill_2
XFILLER_2_367 VPWR VGND sg13g2_fill_2
XFILLER_2_389 VPWR VGND sg13g2_decap_8
XFILLER_5_161 VPWR VGND sg13g2_decap_8
XFILLER_11_477 VPWR VGND sg13g2_decap_8
XFILLER_7_437 VPWR VGND sg13g2_decap_8
X_063_ N2MID[0] net64 VPWR VGND sg13g2_buf_1
XFILLER_3_0 VPWR VGND sg13g2_decap_8
XFILLER_9_98 VPWR VGND sg13g2_decap_8
XFILLER_9_21 VPWR VGND sg13g2_decap_8
XFILLER_6_481 VPWR VGND sg13g2_decap_8
XFILLER_0_56 VPWR VGND sg13g2_decap_8
X_046_ FrameStrobe[14] net38 VPWR VGND sg13g2_buf_1
XFILLER_7_223 VPWR VGND sg13g2_decap_8
XFILLER_0_454 VPWR VGND sg13g2_decap_8
XFILLER_10_509 VPWR VGND sg13g2_fill_2
X_029_ FrameData[29] net22 VPWR VGND sg13g2_buf_1
XANTENNA_4 VPWR VGND FrameData[7] sg13g2_antennanp
XFILLER_6_77 VPWR VGND sg13g2_decap_8
Xoutput41 net41 FrameStrobe_O[17] VPWR VGND sg13g2_buf_1
Xoutput52 net52 FrameStrobe_O[9] VPWR VGND sg13g2_buf_1
Xoutput6 net6 FrameData_O[14] VPWR VGND sg13g2_buf_1
XFILLER_5_513 VPWR VGND sg13g2_decap_8
Xoutput30 net30 FrameData_O[7] VPWR VGND sg13g2_buf_1
Xoutput63 net63 S2BEG[6] VPWR VGND sg13g2_buf_1
Xoutput85 net85 S4BEG[6] VPWR VGND sg13g2_buf_1
Xoutput74 net74 S4BEG[10] VPWR VGND sg13g2_buf_1
Xoutput96 net96 SS4BEG[1] VPWR VGND sg13g2_buf_1
.ends

