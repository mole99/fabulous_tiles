module S_WARMBOOT (BOOT_top,
    CONFIGURED_top,
    Co,
    RESET_top,
    SLOT_top0,
    SLOT_top1,
    SLOT_top2,
    SLOT_top3,
    UserCLK,
    UserCLKo,
    VPWR,
    VGND,
    FrameData,
    FrameData_O,
    FrameStrobe,
    FrameStrobe_O,
    N1BEG,
    N2BEG,
    N2BEGb,
    N4BEG,
    NN4BEG,
    S1END,
    S2END,
    S2MID,
    S4END,
    SS4END);
 output BOOT_top;
 input CONFIGURED_top;
 output Co;
 input RESET_top;
 output SLOT_top0;
 output SLOT_top1;
 output SLOT_top2;
 output SLOT_top3;
 input UserCLK;
 output UserCLKo;
 inout VPWR;
 inout VGND;
 input [31:0] FrameData;
 output [31:0] FrameData_O;
 input [19:0] FrameStrobe;
 output [19:0] FrameStrobe_O;
 output [3:0] N1BEG;
 output [7:0] N2BEG;
 output [7:0] N2BEGb;
 output [15:0] N4BEG;
 output [15:0] NN4BEG;
 input [3:0] S1END;
 input [7:0] S2END;
 input [7:0] S2MID;
 input [15:0] S4END;
 input [15:0] SS4END;

 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire \Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit13.Q ;
 wire \Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit14.Q ;
 wire \Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit15.Q ;
 wire \Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit16.Q ;
 wire \Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit17.Q ;
 wire \Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit18.Q ;
 wire \Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit19.Q ;
 wire \Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit20.Q ;
 wire \Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit21.Q ;
 wire \Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit22.Q ;
 wire \Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit23.Q ;
 wire \Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit24.Q ;
 wire \Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit25.Q ;
 wire \Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit26.Q ;
 wire \Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit27.Q ;
 wire \Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit28.Q ;
 wire \Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit29.Q ;
 wire \Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit30.Q ;
 wire \Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit31.Q ;
 wire \Inst_S_WARMBOOT_switch_matrix.N1BEG0 ;
 wire \Inst_S_WARMBOOT_switch_matrix.N1BEG1 ;
 wire \Inst_S_WARMBOOT_switch_matrix.N1BEG2 ;
 wire \Inst_S_WARMBOOT_switch_matrix.N1BEG3 ;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire net7;
 wire net8;
 wire net9;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net167;

 sg13g2_inv_1 _016_ (.VDD(VPWR),
    .Y(_000_),
    .A(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit19.Q ),
    .VSS(VGND));
 sg13g2_inv_1 _017_ (.VDD(VPWR),
    .Y(_001_),
    .A(net1),
    .VSS(VGND));
 sg13g2_mux4_1 _018_ (.S0(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit17.Q ),
    .A0(net28),
    .A1(net40),
    .A2(net32),
    .A3(net36),
    .S1(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit18.Q ),
    .X(_002_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _019_ (.VDD(VPWR),
    .Y(_003_),
    .A(_002_),
    .VSS(VGND));
 sg13g2_mux2_1 _020_ (.A0(net44),
    .A1(net48),
    .S(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit17.Q ),
    .X(_004_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _021_ (.Y(_005_),
    .B(_004_),
    .A_N(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit18.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _022_ (.A0(net52),
    .A1(net56),
    .S(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit17.Q ),
    .X(_006_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _023_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit18.Q ),
    .A2(_006_),
    .Y(_007_),
    .B1(_000_));
 sg13g2_a221oi_1 _024_ (.VSS(VGND),
    .VDD(VPWR),
    .B2(_007_),
    .C1(_001_),
    .B1(_005_),
    .A1(_000_),
    .Y(net57),
    .A2(_003_));
 sg13g2_mux4_1 _025_ (.S0(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit29.Q ),
    .A0(net44),
    .A1(net48),
    .A2(net52),
    .A3(net56),
    .S1(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit30.Q ),
    .X(_008_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _026_ (.S0(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit29.Q ),
    .A0(net28),
    .A1(net40),
    .A2(net32),
    .A3(net36),
    .S1(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit30.Q ),
    .X(_009_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _027_ (.A0(_009_),
    .A1(_008_),
    .S(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit31.Q ),
    .X(net165),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _028_ (.S0(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit26.Q ),
    .A0(net43),
    .A1(net47),
    .A2(net51),
    .A3(net55),
    .S1(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit27.Q ),
    .X(_010_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _029_ (.S0(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit26.Q ),
    .A0(net27),
    .A1(net39),
    .A2(net31),
    .A3(net35),
    .S1(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit27.Q ),
    .X(_011_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _030_ (.A0(_011_),
    .A1(_010_),
    .S(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit28.Q ),
    .X(net164),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _031_ (.S0(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit23.Q ),
    .A0(net42),
    .A1(net46),
    .A2(net50),
    .A3(net54),
    .S1(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit24.Q ),
    .X(_012_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _032_ (.S0(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit23.Q ),
    .A0(net26),
    .A1(net38),
    .A2(net30),
    .A3(net34),
    .S1(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit24.Q ),
    .X(_013_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _033_ (.A0(_013_),
    .A1(_012_),
    .S(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit25.Q ),
    .X(net163),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _034_ (.S0(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit20.Q ),
    .A0(net41),
    .A1(net45),
    .A2(net49),
    .A3(net53),
    .S1(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit21.Q ),
    .X(_014_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _035_ (.S0(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit20.Q ),
    .A0(net25),
    .A1(net37),
    .A2(net29),
    .A3(net33),
    .S1(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit21.Q ),
    .X(_015_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _036_ (.A0(_015_),
    .A1(_014_),
    .S(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit22.Q ),
    .X(net162),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _037_ (.A0(net25),
    .A1(net24),
    .S(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit16.Q ),
    .X(\Inst_S_WARMBOOT_switch_matrix.N1BEG3 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _038_ (.A0(net26),
    .A1(net24),
    .S(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit15.Q ),
    .X(\Inst_S_WARMBOOT_switch_matrix.N1BEG2 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _039_ (.A0(net27),
    .A1(net24),
    .S(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit14.Q ),
    .X(\Inst_S_WARMBOOT_switch_matrix.N1BEG1 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _040_ (.A0(net28),
    .A1(net24),
    .S(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit13.Q ),
    .X(\Inst_S_WARMBOOT_switch_matrix.N1BEG0 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _041_ (.D(net2),
    .GATE(net7),
    .Q(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit13.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _042_ (.D(net3),
    .GATE(net7),
    .Q(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit14.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _043_ (.D(net4),
    .GATE(net7),
    .Q(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit15.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _044_ (.D(net5),
    .GATE(net7),
    .Q(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit16.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _045_ (.D(net6),
    .GATE(net9),
    .Q(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit17.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _046_ (.D(net10),
    .GATE(net9),
    .Q(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit18.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _047_ (.D(net11),
    .GATE(net7),
    .Q(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit19.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _048_ (.D(net12),
    .GATE(net8),
    .Q(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit20.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _049_ (.D(net13),
    .GATE(net8),
    .Q(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit21.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _050_ (.D(net14),
    .GATE(net8),
    .Q(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit22.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _051_ (.D(net15),
    .GATE(net8),
    .Q(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit23.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _052_ (.D(net16),
    .GATE(net8),
    .Q(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit24.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _053_ (.D(net17),
    .GATE(net8),
    .Q(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit25.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _054_ (.D(net18),
    .GATE(net9),
    .Q(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit26.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _055_ (.D(net19),
    .GATE(net8),
    .Q(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit27.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _056_ (.D(net20),
    .GATE(net9),
    .Q(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit28.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _057_ (.D(net21),
    .GATE(net7),
    .Q(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit29.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _058_ (.D(net22),
    .GATE(net7),
    .Q(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit30.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _059_ (.D(net23),
    .GATE(net7),
    .Q(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit31.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_antennanp ANTENNA_1 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[10]));
 sg13g2_buf_1 _061_ (.A(FrameData[0]),
    .X(net58),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _062_ (.A(FrameData[1]),
    .X(net69),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _063_ (.A(FrameData[2]),
    .X(net80),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _064_ (.A(FrameData[3]),
    .X(net83),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _065_ (.A(FrameData[4]),
    .X(net84),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _066_ (.A(FrameData[5]),
    .X(net85),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _067_ (.A(FrameData[6]),
    .X(net86),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _068_ (.A(FrameData[7]),
    .X(net87),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _069_ (.A(FrameData[8]),
    .X(net88),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _070_ (.A(FrameData[9]),
    .X(net89),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _071_ (.A(FrameData[10]),
    .X(net59),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _072_ (.A(FrameData[11]),
    .X(net60),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _073_ (.A(FrameData[12]),
    .X(net61),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _074_ (.A(net2),
    .X(net62),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _075_ (.A(net3),
    .X(net63),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _076_ (.A(net4),
    .X(net64),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _077_ (.A(net5),
    .X(net65),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _078_ (.A(net6),
    .X(net66),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _079_ (.A(net10),
    .X(net67),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _080_ (.A(net11),
    .X(net68),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _081_ (.A(net12),
    .X(net70),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _082_ (.A(net13),
    .X(net71),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _083_ (.A(net14),
    .X(net72),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _084_ (.A(net15),
    .X(net73),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _085_ (.A(net16),
    .X(net74),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _086_ (.A(net17),
    .X(net75),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _087_ (.A(net18),
    .X(net76),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _088_ (.A(net19),
    .X(net77),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _089_ (.A(net20),
    .X(net78),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _090_ (.A(net21),
    .X(net79),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _091_ (.A(net22),
    .X(net81),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _092_ (.A(net23),
    .X(net82),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _093_ (.A(net8),
    .X(net90),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _094_ (.A(FrameStrobe[1]),
    .X(net101),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _095_ (.A(FrameStrobe[2]),
    .X(net102),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _096_ (.A(FrameStrobe[3]),
    .X(net103),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _097_ (.A(FrameStrobe[4]),
    .X(net104),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _098_ (.A(FrameStrobe[5]),
    .X(net105),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _099_ (.A(FrameStrobe[6]),
    .X(net106),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _100_ (.A(FrameStrobe[7]),
    .X(net107),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _101_ (.A(FrameStrobe[8]),
    .X(net108),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _102_ (.A(FrameStrobe[9]),
    .X(net109),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _103_ (.A(FrameStrobe[10]),
    .X(net91),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _104_ (.A(FrameStrobe[11]),
    .X(net92),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _105_ (.A(FrameStrobe[12]),
    .X(net93),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _106_ (.A(FrameStrobe[13]),
    .X(net94),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _107_ (.A(FrameStrobe[14]),
    .X(net95),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _108_ (.A(FrameStrobe[15]),
    .X(net96),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _109_ (.A(FrameStrobe[16]),
    .X(net97),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _110_ (.A(FrameStrobe[17]),
    .X(net98),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _111_ (.A(FrameStrobe[18]),
    .X(net99),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _112_ (.A(FrameStrobe[19]),
    .X(net100),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _113_ (.A(\Inst_S_WARMBOOT_switch_matrix.N1BEG0 ),
    .X(net110),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _114_ (.A(\Inst_S_WARMBOOT_switch_matrix.N1BEG1 ),
    .X(net111),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _115_ (.A(\Inst_S_WARMBOOT_switch_matrix.N1BEG2 ),
    .X(net112),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _116_ (.A(\Inst_S_WARMBOOT_switch_matrix.N1BEG3 ),
    .X(net113),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _117_ (.A(S2MID[7]),
    .X(net114),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _118_ (.A(S2MID[6]),
    .X(net115),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _119_ (.A(S2MID[5]),
    .X(net116),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _120_ (.A(S2MID[4]),
    .X(net117),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _121_ (.A(net40),
    .X(net118),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _122_ (.A(net39),
    .X(net119),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _123_ (.A(net38),
    .X(net120),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _124_ (.A(net37),
    .X(net121),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _125_ (.A(net36),
    .X(net122),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _126_ (.A(net35),
    .X(net123),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _127_ (.A(net34),
    .X(net124),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _128_ (.A(net33),
    .X(net125),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _129_ (.A(net32),
    .X(net126),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _130_ (.A(net31),
    .X(net127),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _131_ (.A(net30),
    .X(net128),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _132_ (.A(net29),
    .X(net129),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _133_ (.A(S4END[15]),
    .X(net130),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _134_ (.A(S4END[14]),
    .X(net137),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _135_ (.A(S4END[13]),
    .X(net138),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _136_ (.A(S4END[12]),
    .X(net139),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _137_ (.A(S4END[11]),
    .X(net140),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _138_ (.A(S4END[10]),
    .X(net141),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _139_ (.A(S4END[9]),
    .X(net142),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _140_ (.A(S4END[8]),
    .X(net143),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _141_ (.A(net48),
    .X(net144),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _142_ (.A(net47),
    .X(net145),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _143_ (.A(net46),
    .X(net131),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _144_ (.A(net45),
    .X(net132),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _145_ (.A(net44),
    .X(net133),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _146_ (.A(net43),
    .X(net134),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _147_ (.A(net42),
    .X(net135),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _148_ (.A(net41),
    .X(net136),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _149_ (.A(SS4END[15]),
    .X(net146),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _150_ (.A(SS4END[14]),
    .X(net153),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _151_ (.A(SS4END[13]),
    .X(net154),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _152_ (.A(SS4END[12]),
    .X(net155),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _153_ (.A(SS4END[11]),
    .X(net156),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _154_ (.A(SS4END[10]),
    .X(net157),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _155_ (.A(SS4END[9]),
    .X(net158),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _156_ (.A(SS4END[8]),
    .X(net159),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _157_ (.A(net56),
    .X(net160),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _158_ (.A(net55),
    .X(net161),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _159_ (.A(net54),
    .X(net147),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _160_ (.A(net53),
    .X(net148),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _161_ (.A(net52),
    .X(net149),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _162_ (.A(net51),
    .X(net150),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _163_ (.A(net50),
    .X(net151),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _164_ (.A(net49),
    .X(net152),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _165_ (.A(UserCLK),
    .X(net166),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout7 (.A(net9),
    .X(net7),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout8 (.A(net9),
    .X(net8),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout9 (.A(FrameStrobe[0]),
    .X(net9),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input1 (.A(CONFIGURED_top),
    .X(net1),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input2 (.A(FrameData[13]),
    .X(net2),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input3 (.A(FrameData[14]),
    .X(net3),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input4 (.A(FrameData[15]),
    .X(net4),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input5 (.A(FrameData[16]),
    .X(net5),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input6 (.A(FrameData[17]),
    .X(net6),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input7 (.A(FrameData[18]),
    .X(net10),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input8 (.A(FrameData[19]),
    .X(net11),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input9 (.A(FrameData[20]),
    .X(net12),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input10 (.A(FrameData[21]),
    .X(net13),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input11 (.A(FrameData[22]),
    .X(net14),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input12 (.A(FrameData[23]),
    .X(net15),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input13 (.A(FrameData[24]),
    .X(net16),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input14 (.A(FrameData[25]),
    .X(net17),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input15 (.A(FrameData[26]),
    .X(net18),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input16 (.A(FrameData[27]),
    .X(net19),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input17 (.A(FrameData[28]),
    .X(net20),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input18 (.A(FrameData[29]),
    .X(net21),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input19 (.A(FrameData[30]),
    .X(net22),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input20 (.A(FrameData[31]),
    .X(net23),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input21 (.A(RESET_top),
    .X(net24),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input22 (.A(S1END[0]),
    .X(net25),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input23 (.A(S1END[1]),
    .X(net26),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input24 (.A(S1END[2]),
    .X(net27),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input25 (.A(S1END[3]),
    .X(net28),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input26 (.A(S2END[0]),
    .X(net29),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input27 (.A(S2END[1]),
    .X(net30),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input28 (.A(S2END[2]),
    .X(net31),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input29 (.A(S2END[3]),
    .X(net32),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input30 (.A(S2END[4]),
    .X(net33),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input31 (.A(S2END[5]),
    .X(net34),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input32 (.A(S2END[6]),
    .X(net35),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input33 (.A(S2END[7]),
    .X(net36),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input34 (.A(S2MID[0]),
    .X(net37),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input35 (.A(S2MID[1]),
    .X(net38),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input36 (.A(S2MID[2]),
    .X(net39),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input37 (.A(S2MID[3]),
    .X(net40),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input38 (.A(S4END[0]),
    .X(net41),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input39 (.A(S4END[1]),
    .X(net42),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input40 (.A(S4END[2]),
    .X(net43),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input41 (.A(S4END[3]),
    .X(net44),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input42 (.A(S4END[4]),
    .X(net45),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input43 (.A(S4END[5]),
    .X(net46),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input44 (.A(S4END[6]),
    .X(net47),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input45 (.A(S4END[7]),
    .X(net48),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input46 (.A(SS4END[0]),
    .X(net49),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input47 (.A(SS4END[1]),
    .X(net50),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input48 (.A(SS4END[2]),
    .X(net51),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input49 (.A(SS4END[3]),
    .X(net52),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input50 (.A(SS4END[4]),
    .X(net53),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input51 (.A(SS4END[5]),
    .X(net54),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input52 (.A(SS4END[6]),
    .X(net55),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input53 (.A(SS4END[7]),
    .X(net56),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output54 (.A(net57),
    .X(BOOT_top),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output55 (.A(net58),
    .X(FrameData_O[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output56 (.A(net59),
    .X(FrameData_O[10]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output57 (.A(net60),
    .X(FrameData_O[11]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output58 (.A(net61),
    .X(FrameData_O[12]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output59 (.A(net62),
    .X(FrameData_O[13]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output60 (.A(net63),
    .X(FrameData_O[14]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output61 (.A(net64),
    .X(FrameData_O[15]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output62 (.A(net65),
    .X(FrameData_O[16]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output63 (.A(net66),
    .X(FrameData_O[17]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output64 (.A(net67),
    .X(FrameData_O[18]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output65 (.A(net68),
    .X(FrameData_O[19]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output66 (.A(net69),
    .X(FrameData_O[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output67 (.A(net70),
    .X(FrameData_O[20]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output68 (.A(net71),
    .X(FrameData_O[21]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output69 (.A(net72),
    .X(FrameData_O[22]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output70 (.A(net73),
    .X(FrameData_O[23]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output71 (.A(net74),
    .X(FrameData_O[24]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output72 (.A(net75),
    .X(FrameData_O[25]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output73 (.A(net76),
    .X(FrameData_O[26]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output74 (.A(net77),
    .X(FrameData_O[27]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output75 (.A(net78),
    .X(FrameData_O[28]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output76 (.A(net79),
    .X(FrameData_O[29]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output77 (.A(net80),
    .X(FrameData_O[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output78 (.A(net81),
    .X(FrameData_O[30]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output79 (.A(net82),
    .X(FrameData_O[31]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output80 (.A(net83),
    .X(FrameData_O[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output81 (.A(net84),
    .X(FrameData_O[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output82 (.A(net85),
    .X(FrameData_O[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output83 (.A(net86),
    .X(FrameData_O[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output84 (.A(net87),
    .X(FrameData_O[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output85 (.A(net88),
    .X(FrameData_O[8]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output86 (.A(net89),
    .X(FrameData_O[9]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output87 (.A(net90),
    .X(FrameStrobe_O[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output88 (.A(net91),
    .X(FrameStrobe_O[10]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output89 (.A(net92),
    .X(FrameStrobe_O[11]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output90 (.A(net93),
    .X(FrameStrobe_O[12]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output91 (.A(net94),
    .X(FrameStrobe_O[13]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output92 (.A(net95),
    .X(FrameStrobe_O[14]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output93 (.A(net96),
    .X(FrameStrobe_O[15]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output94 (.A(net97),
    .X(FrameStrobe_O[16]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output95 (.A(net98),
    .X(FrameStrobe_O[17]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output96 (.A(net99),
    .X(FrameStrobe_O[18]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output97 (.A(net100),
    .X(FrameStrobe_O[19]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output98 (.A(net101),
    .X(FrameStrobe_O[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output99 (.A(net102),
    .X(FrameStrobe_O[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output100 (.A(net103),
    .X(FrameStrobe_O[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output101 (.A(net104),
    .X(FrameStrobe_O[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output102 (.A(net105),
    .X(FrameStrobe_O[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output103 (.A(net106),
    .X(FrameStrobe_O[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output104 (.A(net107),
    .X(FrameStrobe_O[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output105 (.A(net108),
    .X(FrameStrobe_O[8]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output106 (.A(net109),
    .X(FrameStrobe_O[9]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output107 (.A(net110),
    .X(N1BEG[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output108 (.A(net111),
    .X(N1BEG[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output109 (.A(net112),
    .X(N1BEG[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output110 (.A(net113),
    .X(N1BEG[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output111 (.A(net114),
    .X(N2BEG[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output112 (.A(net115),
    .X(N2BEG[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output113 (.A(net116),
    .X(N2BEG[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output114 (.A(net117),
    .X(N2BEG[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output115 (.A(net118),
    .X(N2BEG[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output116 (.A(net119),
    .X(N2BEG[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output117 (.A(net120),
    .X(N2BEG[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output118 (.A(net121),
    .X(N2BEG[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output119 (.A(net122),
    .X(N2BEGb[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output120 (.A(net123),
    .X(N2BEGb[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output121 (.A(net124),
    .X(N2BEGb[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output122 (.A(net125),
    .X(N2BEGb[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output123 (.A(net126),
    .X(N2BEGb[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output124 (.A(net127),
    .X(N2BEGb[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output125 (.A(net128),
    .X(N2BEGb[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output126 (.A(net129),
    .X(N2BEGb[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output127 (.A(net130),
    .X(N4BEG[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output128 (.A(net131),
    .X(N4BEG[10]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output129 (.A(net132),
    .X(N4BEG[11]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output130 (.A(net133),
    .X(N4BEG[12]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output131 (.A(net134),
    .X(N4BEG[13]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output132 (.A(net135),
    .X(N4BEG[14]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output133 (.A(net136),
    .X(N4BEG[15]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output134 (.A(net137),
    .X(N4BEG[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output135 (.A(net138),
    .X(N4BEG[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output136 (.A(net139),
    .X(N4BEG[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output137 (.A(net140),
    .X(N4BEG[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output138 (.A(net141),
    .X(N4BEG[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output139 (.A(net142),
    .X(N4BEG[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output140 (.A(net143),
    .X(N4BEG[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output141 (.A(net144),
    .X(N4BEG[8]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output142 (.A(net145),
    .X(N4BEG[9]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output143 (.A(net146),
    .X(NN4BEG[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output144 (.A(net147),
    .X(NN4BEG[10]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output145 (.A(net148),
    .X(NN4BEG[11]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output146 (.A(net149),
    .X(NN4BEG[12]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output147 (.A(net150),
    .X(NN4BEG[13]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output148 (.A(net151),
    .X(NN4BEG[14]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output149 (.A(net152),
    .X(NN4BEG[15]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output150 (.A(net153),
    .X(NN4BEG[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output151 (.A(net154),
    .X(NN4BEG[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output152 (.A(net155),
    .X(NN4BEG[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output153 (.A(net156),
    .X(NN4BEG[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output154 (.A(net157),
    .X(NN4BEG[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output155 (.A(net158),
    .X(NN4BEG[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output156 (.A(net159),
    .X(NN4BEG[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output157 (.A(net160),
    .X(NN4BEG[8]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output158 (.A(net161),
    .X(NN4BEG[9]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output159 (.A(net162),
    .X(SLOT_top0),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output160 (.A(net163),
    .X(SLOT_top1),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output161 (.A(net164),
    .X(SLOT_top2),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output162 (.A(net165),
    .X(SLOT_top3),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output163 (.A(net166),
    .X(UserCLKo),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_tielo S_WARMBOOT_164 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net167));
 sg13g2_antennanp ANTENNA_2 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[11]));
 sg13g2_antennanp ANTENNA_3 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[12]));
 sg13g2_antennanp ANTENNA_4 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[2]));
 sg13g2_antennanp ANTENNA_5 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[3]));
 sg13g2_antennanp ANTENNA_6 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[5]));
 sg13g2_antennanp ANTENNA_7 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[6]));
 sg13g2_antennanp ANTENNA_8 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[9]));
 sg13g2_antennanp ANTENNA_9 (.VDD(VPWR),
    .VSS(VGND),
    .A(net68));
 sg13g2_antennanp ANTENNA_10 (.VDD(VPWR),
    .VSS(VGND),
    .A(net79));
 sg13g2_antennanp ANTENNA_11 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[10]));
 sg13g2_antennanp ANTENNA_12 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[11]));
 sg13g2_antennanp ANTENNA_13 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[12]));
 sg13g2_antennanp ANTENNA_14 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[4]));
 sg13g2_antennanp ANTENNA_15 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[6]));
 sg13g2_antennanp ANTENNA_16 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[9]));
 sg13g2_antennanp ANTENNA_17 (.VDD(VPWR),
    .VSS(VGND),
    .A(net62));
 sg13g2_antennanp ANTENNA_18 (.VDD(VPWR),
    .VSS(VGND),
    .A(net68));
 sg13g2_antennanp ANTENNA_19 (.VDD(VPWR),
    .VSS(VGND),
    .A(net81));
 sg13g2_antennanp ANTENNA_20 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[0]));
 sg13g2_antennanp ANTENNA_21 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[10]));
 sg13g2_antennanp ANTENNA_22 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[11]));
 sg13g2_antennanp ANTENNA_23 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[6]));
 sg13g2_antennanp ANTENNA_24 (.VDD(VPWR),
    .VSS(VGND),
    .A(net62));
 sg13g2_antennanp ANTENNA_25 (.VDD(VPWR),
    .VSS(VGND),
    .A(net68));
 sg13g2_antennanp ANTENNA_26 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[0]));
 sg13g2_antennanp ANTENNA_27 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[10]));
 sg13g2_antennanp ANTENNA_28 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[11]));
 sg13g2_antennanp ANTENNA_29 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[6]));
 sg13g2_antennanp ANTENNA_30 (.VDD(VPWR),
    .VSS(VGND),
    .A(net62));
 sg13g2_antennanp ANTENNA_31 (.VDD(VPWR),
    .VSS(VGND),
    .A(net68));
 sg13g2_antennanp ANTENNA_32 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[10]));
 sg13g2_antennanp ANTENNA_33 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[11]));
 sg13g2_antennanp ANTENNA_34 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[6]));
 sg13g2_antennanp ANTENNA_35 (.VDD(VPWR),
    .VSS(VGND),
    .A(net62));
 sg13g2_antennanp ANTENNA_36 (.VDD(VPWR),
    .VSS(VGND),
    .A(net68));
 sg13g2_antennanp ANTENNA_37 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[10]));
 sg13g2_antennanp ANTENNA_38 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[11]));
 sg13g2_antennanp ANTENNA_39 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[6]));
 sg13g2_antennanp ANTENNA_40 (.VDD(VPWR),
    .VSS(VGND),
    .A(net62));
 sg13g2_antennanp ANTENNA_41 (.VDD(VPWR),
    .VSS(VGND),
    .A(net68));
 sg13g2_antennanp ANTENNA_42 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[10]));
 sg13g2_antennanp ANTENNA_43 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[11]));
 sg13g2_antennanp ANTENNA_44 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[6]));
 sg13g2_antennanp ANTENNA_45 (.VDD(VPWR),
    .VSS(VGND),
    .A(net62));
 sg13g2_antennanp ANTENNA_46 (.VDD(VPWR),
    .VSS(VGND),
    .A(net68));
 sg13g2_antennanp ANTENNA_47 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[10]));
 sg13g2_antennanp ANTENNA_48 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[11]));
 sg13g2_antennanp ANTENNA_49 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[4]));
 sg13g2_antennanp ANTENNA_50 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[6]));
 sg13g2_antennanp ANTENNA_51 (.VDD(VPWR),
    .VSS(VGND),
    .A(net68));
 sg13g2_antennanp ANTENNA_52 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[0]));
 sg13g2_antennanp ANTENNA_53 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[10]));
 sg13g2_antennanp ANTENNA_54 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[11]));
 sg13g2_antennanp ANTENNA_55 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[4]));
 sg13g2_antennanp ANTENNA_56 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[7]));
 sg13g2_antennanp ANTENNA_57 (.VDD(VPWR),
    .VSS(VGND),
    .A(net68));
 sg13g2_antennanp ANTENNA_58 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[0]));
 sg13g2_antennanp ANTENNA_59 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[10]));
 sg13g2_antennanp ANTENNA_60 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[11]));
 sg13g2_antennanp ANTENNA_61 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[4]));
 sg13g2_antennanp ANTENNA_62 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[7]));
 sg13g2_antennanp ANTENNA_63 (.VDD(VPWR),
    .VSS(VGND),
    .A(net68));
 sg13g2_decap_8 FILLER_0_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_17 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_24 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_44 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_65 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_97 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_227 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_265 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_293 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_370 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_426 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_433 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_426 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_414 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_370 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_426 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_433 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_12 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_19 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_26 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_440 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_15 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_22 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_29 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_36 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_43 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_50 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_79 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_15 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_22 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_29 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_36 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_43 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_50 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_64 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_71 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_78 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_107 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_12 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_37 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_44 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_51 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_58 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_65 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_79 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_86 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_136 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_178 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_16 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_23 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_30 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_37 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_44 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_51 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_58 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_65 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_79 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_86 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_397 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_24 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_31 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_38 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_45 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_52 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_59 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_66 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_73 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_80 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_227 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_414 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_435 (.VDD(VPWR),
    .VSS(VGND));
 assign Co = net167;
endmodule
