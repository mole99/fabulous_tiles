magic
tech ihp-sg13g2
magscale 1 2
timestamp 1743697575
<< metal1 >>
rect 1152 9848 52128 9872
rect 1152 9808 3688 9848
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 4056 9808 18808 9848
rect 18848 9808 18890 9848
rect 18930 9808 18972 9848
rect 19012 9808 19054 9848
rect 19094 9808 19136 9848
rect 19176 9808 33928 9848
rect 33968 9808 34010 9848
rect 34050 9808 34092 9848
rect 34132 9808 34174 9848
rect 34214 9808 34256 9848
rect 34296 9808 49048 9848
rect 49088 9808 49130 9848
rect 49170 9808 49212 9848
rect 49252 9808 49294 9848
rect 49334 9808 49376 9848
rect 49416 9808 52128 9848
rect 1152 9784 52128 9808
rect 2811 9680 2853 9689
rect 2811 9640 2812 9680
rect 2852 9640 2853 9680
rect 2811 9631 2853 9640
rect 3195 9680 3237 9689
rect 3195 9640 3196 9680
rect 3236 9640 3237 9680
rect 3195 9631 3237 9640
rect 3579 9680 3621 9689
rect 3579 9640 3580 9680
rect 3620 9640 3621 9680
rect 3579 9631 3621 9640
rect 3963 9680 4005 9689
rect 3963 9640 3964 9680
rect 4004 9640 4005 9680
rect 3963 9631 4005 9640
rect 4347 9680 4389 9689
rect 4347 9640 4348 9680
rect 4388 9640 4389 9680
rect 4347 9631 4389 9640
rect 4731 9680 4773 9689
rect 4731 9640 4732 9680
rect 4772 9640 4773 9680
rect 4731 9631 4773 9640
rect 5115 9680 5157 9689
rect 5115 9640 5116 9680
rect 5156 9640 5157 9680
rect 5115 9631 5157 9640
rect 5499 9680 5541 9689
rect 5499 9640 5500 9680
rect 5540 9640 5541 9680
rect 5499 9631 5541 9640
rect 5883 9680 5925 9689
rect 5883 9640 5884 9680
rect 5924 9640 5925 9680
rect 5883 9631 5925 9640
rect 6267 9680 6309 9689
rect 6267 9640 6268 9680
rect 6308 9640 6309 9680
rect 6267 9631 6309 9640
rect 6651 9680 6693 9689
rect 6651 9640 6652 9680
rect 6692 9640 6693 9680
rect 6651 9631 6693 9640
rect 7035 9680 7077 9689
rect 7035 9640 7036 9680
rect 7076 9640 7077 9680
rect 7035 9631 7077 9640
rect 7419 9680 7461 9689
rect 7419 9640 7420 9680
rect 7460 9640 7461 9680
rect 7419 9631 7461 9640
rect 7803 9680 7845 9689
rect 7803 9640 7804 9680
rect 7844 9640 7845 9680
rect 7803 9631 7845 9640
rect 8187 9680 8229 9689
rect 8187 9640 8188 9680
rect 8228 9640 8229 9680
rect 8187 9631 8229 9640
rect 8571 9680 8613 9689
rect 8571 9640 8572 9680
rect 8612 9640 8613 9680
rect 8571 9631 8613 9640
rect 8955 9680 8997 9689
rect 8955 9640 8956 9680
rect 8996 9640 8997 9680
rect 8955 9631 8997 9640
rect 9339 9680 9381 9689
rect 9339 9640 9340 9680
rect 9380 9640 9381 9680
rect 9339 9631 9381 9640
rect 9723 9680 9765 9689
rect 9723 9640 9724 9680
rect 9764 9640 9765 9680
rect 9723 9631 9765 9640
rect 10107 9680 10149 9689
rect 10107 9640 10108 9680
rect 10148 9640 10149 9680
rect 10107 9631 10149 9640
rect 10491 9680 10533 9689
rect 10491 9640 10492 9680
rect 10532 9640 10533 9680
rect 10491 9631 10533 9640
rect 10875 9680 10917 9689
rect 10875 9640 10876 9680
rect 10916 9640 10917 9680
rect 10875 9631 10917 9640
rect 11259 9680 11301 9689
rect 11259 9640 11260 9680
rect 11300 9640 11301 9680
rect 11259 9631 11301 9640
rect 11643 9680 11685 9689
rect 11643 9640 11644 9680
rect 11684 9640 11685 9680
rect 11643 9631 11685 9640
rect 12027 9680 12069 9689
rect 12027 9640 12028 9680
rect 12068 9640 12069 9680
rect 12027 9631 12069 9640
rect 12411 9680 12453 9689
rect 12411 9640 12412 9680
rect 12452 9640 12453 9680
rect 12411 9631 12453 9640
rect 12795 9680 12837 9689
rect 12795 9640 12796 9680
rect 12836 9640 12837 9680
rect 12795 9631 12837 9640
rect 13179 9680 13221 9689
rect 13179 9640 13180 9680
rect 13220 9640 13221 9680
rect 13179 9631 13221 9640
rect 13563 9680 13605 9689
rect 13563 9640 13564 9680
rect 13604 9640 13605 9680
rect 13563 9631 13605 9640
rect 13947 9680 13989 9689
rect 13947 9640 13948 9680
rect 13988 9640 13989 9680
rect 13947 9631 13989 9640
rect 14331 9680 14373 9689
rect 14331 9640 14332 9680
rect 14372 9640 14373 9680
rect 14331 9631 14373 9640
rect 14715 9680 14757 9689
rect 14715 9640 14716 9680
rect 14756 9640 14757 9680
rect 14715 9631 14757 9640
rect 15099 9680 15141 9689
rect 15099 9640 15100 9680
rect 15140 9640 15141 9680
rect 15099 9631 15141 9640
rect 15483 9680 15525 9689
rect 15483 9640 15484 9680
rect 15524 9640 15525 9680
rect 15483 9631 15525 9640
rect 15867 9680 15909 9689
rect 15867 9640 15868 9680
rect 15908 9640 15909 9680
rect 15867 9631 15909 9640
rect 16251 9680 16293 9689
rect 16251 9640 16252 9680
rect 16292 9640 16293 9680
rect 16251 9631 16293 9640
rect 16635 9680 16677 9689
rect 16635 9640 16636 9680
rect 16676 9640 16677 9680
rect 16635 9631 16677 9640
rect 17019 9680 17061 9689
rect 17019 9640 17020 9680
rect 17060 9640 17061 9680
rect 17019 9631 17061 9640
rect 17403 9680 17445 9689
rect 17403 9640 17404 9680
rect 17444 9640 17445 9680
rect 17403 9631 17445 9640
rect 17787 9680 17829 9689
rect 17787 9640 17788 9680
rect 17828 9640 17829 9680
rect 17787 9631 17829 9640
rect 18171 9680 18213 9689
rect 18171 9640 18172 9680
rect 18212 9640 18213 9680
rect 18171 9631 18213 9640
rect 18555 9680 18597 9689
rect 18555 9640 18556 9680
rect 18596 9640 18597 9680
rect 18555 9631 18597 9640
rect 19323 9680 19365 9689
rect 19323 9640 19324 9680
rect 19364 9640 19365 9680
rect 19323 9631 19365 9640
rect 19707 9680 19749 9689
rect 19707 9640 19708 9680
rect 19748 9640 19749 9680
rect 19707 9631 19749 9640
rect 20091 9680 20133 9689
rect 20091 9640 20092 9680
rect 20132 9640 20133 9680
rect 20091 9631 20133 9640
rect 20475 9680 20517 9689
rect 20475 9640 20476 9680
rect 20516 9640 20517 9680
rect 20475 9631 20517 9640
rect 20859 9680 20901 9689
rect 20859 9640 20860 9680
rect 20900 9640 20901 9680
rect 20859 9631 20901 9640
rect 21243 9680 21285 9689
rect 21243 9640 21244 9680
rect 21284 9640 21285 9680
rect 21243 9631 21285 9640
rect 21627 9680 21669 9689
rect 21627 9640 21628 9680
rect 21668 9640 21669 9680
rect 21627 9631 21669 9640
rect 22011 9680 22053 9689
rect 22011 9640 22012 9680
rect 22052 9640 22053 9680
rect 22011 9631 22053 9640
rect 22395 9680 22437 9689
rect 22395 9640 22396 9680
rect 22436 9640 22437 9680
rect 22395 9631 22437 9640
rect 42747 9680 42789 9689
rect 42747 9640 42748 9680
rect 42788 9640 42789 9680
rect 42747 9631 42789 9640
rect 43131 9680 43173 9689
rect 43131 9640 43132 9680
rect 43172 9640 43173 9680
rect 43131 9631 43173 9640
rect 43515 9680 43557 9689
rect 43515 9640 43516 9680
rect 43556 9640 43557 9680
rect 43515 9631 43557 9640
rect 43899 9680 43941 9689
rect 43899 9640 43900 9680
rect 43940 9640 43941 9680
rect 43899 9631 43941 9640
rect 44283 9680 44325 9689
rect 44283 9640 44284 9680
rect 44324 9640 44325 9680
rect 44283 9631 44325 9640
rect 44667 9680 44709 9689
rect 44667 9640 44668 9680
rect 44708 9640 44709 9680
rect 44667 9631 44709 9640
rect 45051 9680 45093 9689
rect 45051 9640 45052 9680
rect 45092 9640 45093 9680
rect 45051 9631 45093 9640
rect 45435 9680 45477 9689
rect 45435 9640 45436 9680
rect 45476 9640 45477 9680
rect 45435 9631 45477 9640
rect 45819 9680 45861 9689
rect 45819 9640 45820 9680
rect 45860 9640 45861 9680
rect 45819 9631 45861 9640
rect 46203 9680 46245 9689
rect 46203 9640 46204 9680
rect 46244 9640 46245 9680
rect 46203 9631 46245 9640
rect 46587 9680 46629 9689
rect 46587 9640 46588 9680
rect 46628 9640 46629 9680
rect 46587 9631 46629 9640
rect 46971 9680 47013 9689
rect 46971 9640 46972 9680
rect 47012 9640 47013 9680
rect 46971 9631 47013 9640
rect 47355 9680 47397 9689
rect 47355 9640 47356 9680
rect 47396 9640 47397 9680
rect 47355 9631 47397 9640
rect 47739 9680 47781 9689
rect 47739 9640 47740 9680
rect 47780 9640 47781 9680
rect 47739 9631 47781 9640
rect 48123 9680 48165 9689
rect 48123 9640 48124 9680
rect 48164 9640 48165 9680
rect 48123 9631 48165 9640
rect 48507 9680 48549 9689
rect 48507 9640 48508 9680
rect 48548 9640 48549 9680
rect 48507 9631 48549 9640
rect 48891 9680 48933 9689
rect 48891 9640 48892 9680
rect 48932 9640 48933 9680
rect 48891 9631 48933 9640
rect 49275 9680 49317 9689
rect 49275 9640 49276 9680
rect 49316 9640 49317 9680
rect 49275 9631 49317 9640
rect 50043 9680 50085 9689
rect 50043 9640 50044 9680
rect 50084 9640 50085 9680
rect 50043 9631 50085 9640
rect 50427 9680 50469 9689
rect 50427 9640 50428 9680
rect 50468 9640 50469 9680
rect 50427 9631 50469 9640
rect 18939 9596 18981 9605
rect 18939 9556 18940 9596
rect 18980 9556 18981 9596
rect 18939 9547 18981 9556
rect 49659 9596 49701 9605
rect 49659 9556 49660 9596
rect 49700 9556 49701 9596
rect 49659 9547 49701 9556
rect 3051 9512 3093 9521
rect 3051 9472 3052 9512
rect 3092 9472 3093 9512
rect 3051 9463 3093 9472
rect 3435 9512 3477 9521
rect 3435 9472 3436 9512
rect 3476 9472 3477 9512
rect 3435 9463 3477 9472
rect 3819 9512 3861 9521
rect 3819 9472 3820 9512
rect 3860 9472 3861 9512
rect 3819 9463 3861 9472
rect 4203 9512 4245 9521
rect 4203 9472 4204 9512
rect 4244 9472 4245 9512
rect 4203 9463 4245 9472
rect 4587 9512 4629 9521
rect 4587 9472 4588 9512
rect 4628 9472 4629 9512
rect 4587 9463 4629 9472
rect 4971 9512 5013 9521
rect 4971 9472 4972 9512
rect 5012 9472 5013 9512
rect 4971 9463 5013 9472
rect 5355 9512 5397 9521
rect 5355 9472 5356 9512
rect 5396 9472 5397 9512
rect 5355 9463 5397 9472
rect 5739 9512 5781 9521
rect 5739 9472 5740 9512
rect 5780 9472 5781 9512
rect 5739 9463 5781 9472
rect 6123 9512 6165 9521
rect 6123 9472 6124 9512
rect 6164 9472 6165 9512
rect 6123 9463 6165 9472
rect 6507 9512 6549 9521
rect 6507 9472 6508 9512
rect 6548 9472 6549 9512
rect 6507 9463 6549 9472
rect 6891 9512 6933 9521
rect 6891 9472 6892 9512
rect 6932 9472 6933 9512
rect 6891 9463 6933 9472
rect 7275 9512 7317 9521
rect 7275 9472 7276 9512
rect 7316 9472 7317 9512
rect 7275 9463 7317 9472
rect 7659 9512 7701 9521
rect 7659 9472 7660 9512
rect 7700 9472 7701 9512
rect 7659 9463 7701 9472
rect 8043 9512 8085 9521
rect 8043 9472 8044 9512
rect 8084 9472 8085 9512
rect 8043 9463 8085 9472
rect 8427 9512 8469 9521
rect 8427 9472 8428 9512
rect 8468 9472 8469 9512
rect 8427 9463 8469 9472
rect 8811 9512 8853 9521
rect 8811 9472 8812 9512
rect 8852 9472 8853 9512
rect 8811 9463 8853 9472
rect 9195 9512 9237 9521
rect 9195 9472 9196 9512
rect 9236 9472 9237 9512
rect 9195 9463 9237 9472
rect 9579 9512 9621 9521
rect 9579 9472 9580 9512
rect 9620 9472 9621 9512
rect 9579 9463 9621 9472
rect 9963 9512 10005 9521
rect 9963 9472 9964 9512
rect 10004 9472 10005 9512
rect 9963 9463 10005 9472
rect 10347 9512 10389 9521
rect 10347 9472 10348 9512
rect 10388 9472 10389 9512
rect 10347 9463 10389 9472
rect 10731 9512 10773 9521
rect 10731 9472 10732 9512
rect 10772 9472 10773 9512
rect 10731 9463 10773 9472
rect 11115 9512 11157 9521
rect 11115 9472 11116 9512
rect 11156 9472 11157 9512
rect 11115 9463 11157 9472
rect 11499 9512 11541 9521
rect 11499 9472 11500 9512
rect 11540 9472 11541 9512
rect 11499 9463 11541 9472
rect 11883 9512 11925 9521
rect 11883 9472 11884 9512
rect 11924 9472 11925 9512
rect 11883 9463 11925 9472
rect 12267 9512 12309 9521
rect 12267 9472 12268 9512
rect 12308 9472 12309 9512
rect 12267 9463 12309 9472
rect 12651 9512 12693 9521
rect 12651 9472 12652 9512
rect 12692 9472 12693 9512
rect 12651 9463 12693 9472
rect 13035 9512 13077 9521
rect 13035 9472 13036 9512
rect 13076 9472 13077 9512
rect 13035 9463 13077 9472
rect 13419 9512 13461 9521
rect 13419 9472 13420 9512
rect 13460 9472 13461 9512
rect 13419 9463 13461 9472
rect 13803 9512 13845 9521
rect 13803 9472 13804 9512
rect 13844 9472 13845 9512
rect 13803 9463 13845 9472
rect 14187 9512 14229 9521
rect 14187 9472 14188 9512
rect 14228 9472 14229 9512
rect 14187 9463 14229 9472
rect 14571 9512 14613 9521
rect 14571 9472 14572 9512
rect 14612 9472 14613 9512
rect 14571 9463 14613 9472
rect 14955 9512 14997 9521
rect 14955 9472 14956 9512
rect 14996 9472 14997 9512
rect 14955 9463 14997 9472
rect 15339 9512 15381 9521
rect 15339 9472 15340 9512
rect 15380 9472 15381 9512
rect 15339 9463 15381 9472
rect 15723 9512 15765 9521
rect 15723 9472 15724 9512
rect 15764 9472 15765 9512
rect 15723 9463 15765 9472
rect 16107 9512 16149 9521
rect 16107 9472 16108 9512
rect 16148 9472 16149 9512
rect 16107 9463 16149 9472
rect 16491 9512 16533 9521
rect 16491 9472 16492 9512
rect 16532 9472 16533 9512
rect 16491 9463 16533 9472
rect 16875 9512 16917 9521
rect 16875 9472 16876 9512
rect 16916 9472 16917 9512
rect 16875 9463 16917 9472
rect 17259 9512 17301 9521
rect 17259 9472 17260 9512
rect 17300 9472 17301 9512
rect 17259 9463 17301 9472
rect 17643 9512 17685 9521
rect 17643 9472 17644 9512
rect 17684 9472 17685 9512
rect 17643 9463 17685 9472
rect 18027 9512 18069 9521
rect 18027 9472 18028 9512
rect 18068 9472 18069 9512
rect 18027 9463 18069 9472
rect 18411 9512 18453 9521
rect 18411 9472 18412 9512
rect 18452 9472 18453 9512
rect 18411 9463 18453 9472
rect 18795 9512 18837 9521
rect 18795 9472 18796 9512
rect 18836 9472 18837 9512
rect 18795 9463 18837 9472
rect 19179 9512 19221 9521
rect 19179 9472 19180 9512
rect 19220 9472 19221 9512
rect 19179 9463 19221 9472
rect 19563 9512 19605 9521
rect 19563 9472 19564 9512
rect 19604 9472 19605 9512
rect 19563 9463 19605 9472
rect 19947 9512 19989 9521
rect 19947 9472 19948 9512
rect 19988 9472 19989 9512
rect 19947 9463 19989 9472
rect 20331 9512 20373 9521
rect 20331 9472 20332 9512
rect 20372 9472 20373 9512
rect 20331 9463 20373 9472
rect 20715 9512 20757 9521
rect 20715 9472 20716 9512
rect 20756 9472 20757 9512
rect 20715 9463 20757 9472
rect 21099 9512 21141 9521
rect 21099 9472 21100 9512
rect 21140 9472 21141 9512
rect 21099 9463 21141 9472
rect 21483 9512 21525 9521
rect 21483 9472 21484 9512
rect 21524 9472 21525 9512
rect 21483 9463 21525 9472
rect 21867 9512 21909 9521
rect 21867 9472 21868 9512
rect 21908 9472 21909 9512
rect 21867 9463 21909 9472
rect 22251 9512 22293 9521
rect 22251 9472 22252 9512
rect 22292 9472 22293 9512
rect 22251 9463 22293 9472
rect 22635 9512 22677 9521
rect 22635 9472 22636 9512
rect 22676 9472 22677 9512
rect 22635 9463 22677 9472
rect 42987 9512 43029 9521
rect 42987 9472 42988 9512
rect 43028 9472 43029 9512
rect 42987 9463 43029 9472
rect 43371 9512 43413 9521
rect 43371 9472 43372 9512
rect 43412 9472 43413 9512
rect 43371 9463 43413 9472
rect 43755 9512 43797 9521
rect 43755 9472 43756 9512
rect 43796 9472 43797 9512
rect 43755 9463 43797 9472
rect 44139 9512 44181 9521
rect 44139 9472 44140 9512
rect 44180 9472 44181 9512
rect 44139 9463 44181 9472
rect 44523 9512 44565 9521
rect 44523 9472 44524 9512
rect 44564 9472 44565 9512
rect 44523 9463 44565 9472
rect 44907 9512 44949 9521
rect 44907 9472 44908 9512
rect 44948 9472 44949 9512
rect 44907 9463 44949 9472
rect 45291 9512 45333 9521
rect 45291 9472 45292 9512
rect 45332 9472 45333 9512
rect 45291 9463 45333 9472
rect 45675 9512 45717 9521
rect 45675 9472 45676 9512
rect 45716 9472 45717 9512
rect 45675 9463 45717 9472
rect 46059 9512 46101 9521
rect 46059 9472 46060 9512
rect 46100 9472 46101 9512
rect 46059 9463 46101 9472
rect 46443 9512 46485 9521
rect 46443 9472 46444 9512
rect 46484 9472 46485 9512
rect 46443 9463 46485 9472
rect 46827 9512 46869 9521
rect 46827 9472 46828 9512
rect 46868 9472 46869 9512
rect 46827 9463 46869 9472
rect 47211 9512 47253 9521
rect 47211 9472 47212 9512
rect 47252 9472 47253 9512
rect 47211 9463 47253 9472
rect 47595 9512 47637 9521
rect 47595 9472 47596 9512
rect 47636 9472 47637 9512
rect 47595 9463 47637 9472
rect 47979 9512 48021 9521
rect 47979 9472 47980 9512
rect 48020 9472 48021 9512
rect 47979 9463 48021 9472
rect 48363 9512 48405 9521
rect 48363 9472 48364 9512
rect 48404 9472 48405 9512
rect 48363 9463 48405 9472
rect 48747 9512 48789 9521
rect 48747 9472 48748 9512
rect 48788 9472 48789 9512
rect 48747 9463 48789 9472
rect 49131 9512 49173 9521
rect 49131 9472 49132 9512
rect 49172 9472 49173 9512
rect 49131 9463 49173 9472
rect 49515 9512 49557 9521
rect 49515 9472 49516 9512
rect 49556 9472 49557 9512
rect 49515 9463 49557 9472
rect 49899 9512 49941 9521
rect 49899 9472 49900 9512
rect 49940 9472 49941 9512
rect 49899 9463 49941 9472
rect 50283 9512 50325 9521
rect 50283 9472 50284 9512
rect 50324 9472 50325 9512
rect 50283 9463 50325 9472
rect 50667 9512 50709 9521
rect 50667 9472 50668 9512
rect 50708 9472 50709 9512
rect 50667 9463 50709 9472
rect 51051 9512 51093 9521
rect 51051 9472 51052 9512
rect 51092 9472 51093 9512
rect 51051 9463 51093 9472
rect 51435 9512 51477 9521
rect 51435 9472 51436 9512
rect 51476 9472 51477 9512
rect 51435 9463 51477 9472
rect 51819 9512 51861 9521
rect 51819 9472 51820 9512
rect 51860 9472 51861 9512
rect 51819 9463 51861 9472
rect 51291 9344 51333 9353
rect 51291 9304 51292 9344
rect 51332 9304 51333 9344
rect 51291 9295 51333 9304
rect 51675 9260 51717 9269
rect 51675 9220 51676 9260
rect 51716 9220 51717 9260
rect 51675 9211 51717 9220
rect 52059 9260 52101 9269
rect 52059 9220 52060 9260
rect 52100 9220 52101 9260
rect 52059 9211 52101 9220
rect 1152 9092 52128 9116
rect 1152 9052 4928 9092
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 5296 9052 20048 9092
rect 20088 9052 20130 9092
rect 20170 9052 20212 9092
rect 20252 9052 20294 9092
rect 20334 9052 20376 9092
rect 20416 9052 35168 9092
rect 35208 9052 35250 9092
rect 35290 9052 35332 9092
rect 35372 9052 35414 9092
rect 35454 9052 35496 9092
rect 35536 9052 50288 9092
rect 50328 9052 50370 9092
rect 50410 9052 50452 9092
rect 50492 9052 50534 9092
rect 50574 9052 50616 9092
rect 50656 9052 52128 9092
rect 1152 9028 52128 9052
rect 21627 8924 21669 8933
rect 21627 8884 21628 8924
rect 21668 8884 21669 8924
rect 21627 8875 21669 8884
rect 23067 8924 23109 8933
rect 23067 8884 23068 8924
rect 23108 8884 23109 8924
rect 23067 8875 23109 8884
rect 23643 8924 23685 8933
rect 23643 8884 23644 8924
rect 23684 8884 23685 8924
rect 23643 8875 23685 8884
rect 27003 8924 27045 8933
rect 27003 8884 27004 8924
rect 27044 8884 27045 8924
rect 27003 8875 27045 8884
rect 28155 8924 28197 8933
rect 28155 8884 28156 8924
rect 28196 8884 28197 8924
rect 28155 8875 28197 8884
rect 28923 8924 28965 8933
rect 28923 8884 28924 8924
rect 28964 8884 28965 8924
rect 28923 8875 28965 8884
rect 29691 8924 29733 8933
rect 29691 8884 29692 8924
rect 29732 8884 29733 8924
rect 29691 8875 29733 8884
rect 50139 8924 50181 8933
rect 50139 8884 50140 8924
rect 50180 8884 50181 8924
rect 50139 8875 50181 8884
rect 50523 8924 50565 8933
rect 50523 8884 50524 8924
rect 50564 8884 50565 8924
rect 50523 8875 50565 8884
rect 50907 8924 50949 8933
rect 50907 8884 50908 8924
rect 50948 8884 50949 8924
rect 50907 8875 50949 8884
rect 51291 8924 51333 8933
rect 51291 8884 51292 8924
rect 51332 8884 51333 8924
rect 51291 8875 51333 8884
rect 29307 8840 29349 8849
rect 29307 8800 29308 8840
rect 29348 8800 29349 8840
rect 29307 8791 29349 8800
rect 21867 8672 21909 8681
rect 21867 8632 21868 8672
rect 21908 8632 21909 8672
rect 21867 8623 21909 8632
rect 22347 8672 22389 8681
rect 22347 8632 22348 8672
rect 22388 8632 22389 8672
rect 22347 8623 22389 8632
rect 22731 8672 22773 8681
rect 22731 8632 22732 8672
rect 22772 8632 22773 8672
rect 22731 8623 22773 8632
rect 23307 8672 23349 8681
rect 23307 8632 23308 8672
rect 23348 8632 23349 8672
rect 23307 8623 23349 8632
rect 23883 8672 23925 8681
rect 23883 8632 23884 8672
rect 23924 8632 23925 8672
rect 23883 8623 23925 8632
rect 26763 8672 26805 8681
rect 26763 8632 26764 8672
rect 26804 8632 26805 8672
rect 26763 8623 26805 8632
rect 27147 8672 27189 8681
rect 27147 8632 27148 8672
rect 27188 8632 27189 8672
rect 27147 8623 27189 8632
rect 27531 8672 27573 8681
rect 27531 8632 27532 8672
rect 27572 8632 27573 8672
rect 27531 8623 27573 8632
rect 27771 8672 27813 8681
rect 27771 8632 27772 8672
rect 27812 8632 27813 8672
rect 27771 8623 27813 8632
rect 27946 8672 28004 8673
rect 27946 8632 27955 8672
rect 27995 8632 28004 8672
rect 27946 8631 28004 8632
rect 28299 8672 28341 8681
rect 28299 8632 28300 8672
rect 28340 8632 28341 8672
rect 28299 8623 28341 8632
rect 28539 8672 28581 8681
rect 28539 8632 28540 8672
rect 28580 8632 28581 8672
rect 28539 8623 28581 8632
rect 28683 8672 28725 8681
rect 28683 8632 28684 8672
rect 28724 8632 28725 8672
rect 28683 8623 28725 8632
rect 29067 8672 29109 8681
rect 29067 8632 29068 8672
rect 29108 8632 29109 8672
rect 29067 8623 29109 8632
rect 29451 8672 29493 8681
rect 29451 8632 29452 8672
rect 29492 8632 29493 8672
rect 29451 8623 29493 8632
rect 31227 8672 31269 8681
rect 31227 8632 31228 8672
rect 31268 8632 31269 8672
rect 31227 8623 31269 8632
rect 31467 8672 31509 8681
rect 31467 8632 31468 8672
rect 31508 8632 31509 8672
rect 31467 8623 31509 8632
rect 49899 8672 49941 8681
rect 49899 8632 49900 8672
rect 49940 8632 49941 8672
rect 49899 8623 49941 8632
rect 50283 8672 50325 8681
rect 50283 8632 50284 8672
rect 50324 8632 50325 8672
rect 50283 8623 50325 8632
rect 50667 8672 50709 8681
rect 50667 8632 50668 8672
rect 50708 8632 50709 8672
rect 50667 8623 50709 8632
rect 51051 8672 51093 8681
rect 51051 8632 51052 8672
rect 51092 8632 51093 8672
rect 51051 8623 51093 8632
rect 51435 8672 51477 8681
rect 51435 8632 51436 8672
rect 51476 8632 51477 8672
rect 51435 8623 51477 8632
rect 51819 8672 51861 8681
rect 51819 8632 51820 8672
rect 51860 8632 51861 8672
rect 51819 8623 51861 8632
rect 27387 8588 27429 8597
rect 27387 8548 27388 8588
rect 27428 8548 27429 8588
rect 27387 8539 27429 8548
rect 22107 8504 22149 8513
rect 22107 8464 22108 8504
rect 22148 8464 22149 8504
rect 22107 8455 22149 8464
rect 22491 8504 22533 8513
rect 22491 8464 22492 8504
rect 22532 8464 22533 8504
rect 22491 8455 22533 8464
rect 51675 8504 51717 8513
rect 51675 8464 51676 8504
rect 51716 8464 51717 8504
rect 51675 8455 51717 8464
rect 52059 8504 52101 8513
rect 52059 8464 52060 8504
rect 52100 8464 52101 8504
rect 52059 8455 52101 8464
rect 1152 8336 52128 8360
rect 1152 8296 3688 8336
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 4056 8296 18808 8336
rect 18848 8296 18890 8336
rect 18930 8296 18972 8336
rect 19012 8296 19054 8336
rect 19094 8296 19136 8336
rect 19176 8296 33928 8336
rect 33968 8296 34010 8336
rect 34050 8296 34092 8336
rect 34132 8296 34174 8336
rect 34214 8296 34256 8336
rect 34296 8296 49048 8336
rect 49088 8296 49130 8336
rect 49170 8296 49212 8336
rect 49252 8296 49294 8336
rect 49334 8296 49376 8336
rect 49416 8296 52128 8336
rect 1152 8272 52128 8296
rect 3483 8168 3525 8177
rect 3483 8128 3484 8168
rect 3524 8128 3525 8168
rect 3483 8119 3525 8128
rect 4347 8168 4389 8177
rect 4347 8128 4348 8168
rect 4388 8128 4389 8168
rect 4347 8119 4389 8128
rect 6363 8168 6405 8177
rect 6363 8128 6364 8168
rect 6404 8128 6405 8168
rect 6363 8119 6405 8128
rect 7803 8168 7845 8177
rect 7803 8128 7804 8168
rect 7844 8128 7845 8168
rect 7803 8119 7845 8128
rect 10203 8168 10245 8177
rect 10203 8128 10204 8168
rect 10244 8128 10245 8168
rect 10203 8119 10245 8128
rect 15291 8168 15333 8177
rect 15291 8128 15292 8168
rect 15332 8128 15333 8168
rect 15291 8119 15333 8128
rect 15675 8168 15717 8177
rect 15675 8128 15676 8168
rect 15716 8128 15717 8168
rect 15675 8119 15717 8128
rect 16059 8168 16101 8177
rect 16059 8128 16060 8168
rect 16100 8128 16101 8168
rect 16059 8119 16101 8128
rect 16443 8168 16485 8177
rect 16443 8128 16444 8168
rect 16484 8128 16485 8168
rect 16443 8119 16485 8128
rect 16827 8168 16869 8177
rect 16827 8128 16828 8168
rect 16868 8128 16869 8168
rect 16827 8119 16869 8128
rect 17595 8168 17637 8177
rect 17595 8128 17596 8168
rect 17636 8128 17637 8168
rect 17595 8119 17637 8128
rect 17979 8168 18021 8177
rect 17979 8128 17980 8168
rect 18020 8128 18021 8168
rect 17979 8119 18021 8128
rect 18363 8168 18405 8177
rect 18363 8128 18364 8168
rect 18404 8128 18405 8168
rect 18363 8119 18405 8128
rect 19035 8168 19077 8177
rect 19035 8128 19036 8168
rect 19076 8128 19077 8168
rect 19035 8119 19077 8128
rect 20763 8168 20805 8177
rect 20763 8128 20764 8168
rect 20804 8128 20805 8168
rect 20763 8119 20805 8128
rect 32763 8168 32805 8177
rect 32763 8128 32764 8168
rect 32804 8128 32805 8168
rect 32763 8119 32805 8128
rect 37083 8168 37125 8177
rect 37083 8128 37084 8168
rect 37124 8128 37125 8168
rect 37083 8119 37125 8128
rect 37467 8168 37509 8177
rect 37467 8128 37468 8168
rect 37508 8128 37509 8168
rect 37467 8119 37509 8128
rect 38139 8168 38181 8177
rect 38139 8128 38140 8168
rect 38180 8128 38181 8168
rect 38139 8119 38181 8128
rect 51291 8168 51333 8177
rect 51291 8128 51292 8168
rect 51332 8128 51333 8168
rect 51291 8119 51333 8128
rect 5499 8084 5541 8093
rect 5499 8044 5500 8084
rect 5540 8044 5541 8084
rect 5499 8035 5541 8044
rect 11931 8084 11973 8093
rect 11931 8044 11932 8084
rect 11972 8044 11973 8084
rect 11931 8035 11973 8044
rect 17211 8084 17253 8093
rect 17211 8044 17212 8084
rect 17252 8044 17253 8084
rect 17211 8035 17253 8044
rect 19419 8084 19461 8093
rect 19419 8044 19420 8084
rect 19460 8044 19461 8084
rect 19419 8035 19461 8044
rect 20283 8084 20325 8093
rect 20283 8044 20284 8084
rect 20324 8044 20325 8084
rect 20283 8035 20325 8044
rect 28635 8084 28677 8093
rect 28635 8044 28636 8084
rect 28676 8044 28677 8084
rect 28635 8035 28677 8044
rect 35067 8084 35109 8093
rect 35067 8044 35068 8084
rect 35108 8044 35109 8084
rect 35067 8035 35109 8044
rect 39387 8084 39429 8093
rect 39387 8044 39388 8084
rect 39428 8044 39429 8084
rect 39387 8035 39429 8044
rect 3243 8000 3285 8009
rect 3243 7960 3244 8000
rect 3284 7960 3285 8000
rect 3243 7951 3285 7960
rect 4587 8000 4629 8009
rect 4587 7960 4588 8000
rect 4628 7960 4629 8000
rect 4587 7951 4629 7960
rect 5259 8000 5301 8009
rect 5259 7960 5260 8000
rect 5300 7960 5301 8000
rect 5259 7951 5301 7960
rect 6123 8000 6165 8009
rect 6123 7960 6124 8000
rect 6164 7960 6165 8000
rect 6123 7951 6165 7960
rect 8043 8000 8085 8009
rect 8043 7960 8044 8000
rect 8084 7960 8085 8000
rect 8043 7951 8085 7960
rect 8427 8000 8469 8009
rect 8427 7960 8428 8000
rect 8468 7960 8469 8000
rect 8427 7951 8469 7960
rect 10443 8000 10485 8009
rect 10443 7960 10444 8000
rect 10484 7960 10485 8000
rect 10443 7951 10485 7960
rect 10587 8000 10629 8009
rect 10587 7960 10588 8000
rect 10628 7960 10629 8000
rect 10587 7951 10629 7960
rect 10827 8000 10869 8009
rect 10827 7960 10828 8000
rect 10868 7960 10869 8000
rect 10827 7951 10869 7960
rect 12171 8000 12213 8009
rect 12171 7960 12172 8000
rect 12212 7960 12213 8000
rect 12171 7951 12213 7960
rect 15531 8000 15573 8009
rect 15531 7960 15532 8000
rect 15572 7960 15573 8000
rect 15531 7951 15573 7960
rect 15915 8000 15957 8009
rect 15915 7960 15916 8000
rect 15956 7960 15957 8000
rect 15915 7951 15957 7960
rect 16299 8000 16341 8009
rect 16299 7960 16300 8000
rect 16340 7960 16341 8000
rect 16299 7951 16341 7960
rect 16683 8000 16725 8009
rect 16683 7960 16684 8000
rect 16724 7960 16725 8000
rect 16683 7951 16725 7960
rect 17067 8000 17109 8009
rect 17067 7960 17068 8000
rect 17108 7960 17109 8000
rect 17067 7951 17109 7960
rect 17451 8000 17493 8009
rect 17451 7960 17452 8000
rect 17492 7960 17493 8000
rect 17451 7951 17493 7960
rect 17835 8000 17877 8009
rect 17835 7960 17836 8000
rect 17876 7960 17877 8000
rect 17835 7951 17877 7960
rect 18219 8000 18261 8009
rect 18219 7960 18220 8000
rect 18260 7960 18261 8000
rect 18219 7951 18261 7960
rect 18603 8000 18645 8009
rect 18603 7960 18604 8000
rect 18644 7960 18645 8000
rect 18603 7951 18645 7960
rect 19275 8000 19317 8009
rect 19275 7960 19276 8000
rect 19316 7960 19317 8000
rect 19275 7951 19317 7960
rect 19659 8000 19701 8009
rect 19659 7960 19660 8000
rect 19700 7960 19701 8000
rect 19659 7951 19701 7960
rect 20523 8000 20565 8009
rect 20523 7960 20524 8000
rect 20564 7960 20565 8000
rect 20523 7951 20565 7960
rect 21003 8000 21045 8009
rect 21003 7960 21004 8000
rect 21044 7960 21045 8000
rect 21003 7951 21045 7960
rect 28395 8000 28437 8009
rect 28395 7960 28396 8000
rect 28436 7960 28437 8000
rect 28395 7951 28437 7960
rect 33003 8000 33045 8009
rect 33003 7960 33004 8000
rect 33044 7960 33045 8000
rect 33003 7951 33045 7960
rect 33387 8000 33429 8009
rect 33387 7960 33388 8000
rect 33428 7960 33429 8000
rect 33387 7951 33429 7960
rect 33771 8000 33813 8009
rect 33771 7960 33772 8000
rect 33812 7960 33813 8000
rect 33771 7951 33813 7960
rect 34923 8000 34965 8009
rect 34923 7960 34924 8000
rect 34964 7960 34965 8000
rect 34923 7951 34965 7960
rect 35307 8000 35349 8009
rect 35307 7960 35308 8000
rect 35348 7960 35349 8000
rect 35307 7951 35349 7960
rect 35691 8000 35733 8009
rect 35691 7960 35692 8000
rect 35732 7960 35733 8000
rect 35691 7951 35733 7960
rect 36075 8000 36117 8009
rect 36075 7960 36076 8000
rect 36116 7960 36117 8000
rect 36075 7951 36117 7960
rect 36363 8000 36405 8009
rect 36363 7960 36364 8000
rect 36404 7960 36405 8000
rect 36363 7951 36405 7960
rect 36747 8000 36789 8009
rect 36747 7960 36748 8000
rect 36788 7960 36789 8000
rect 36747 7951 36789 7960
rect 37323 8000 37365 8009
rect 37323 7960 37324 8000
rect 37364 7960 37365 8000
rect 37323 7951 37365 7960
rect 37707 8000 37749 8009
rect 37707 7960 37708 8000
rect 37748 7960 37749 8000
rect 37707 7951 37749 7960
rect 37899 8000 37941 8009
rect 37899 7960 37900 8000
rect 37940 7960 37941 8000
rect 37899 7951 37941 7960
rect 38235 8000 38277 8009
rect 38235 7960 38236 8000
rect 38276 7960 38277 8000
rect 38235 7951 38277 7960
rect 38475 8000 38517 8009
rect 38475 7960 38476 8000
rect 38516 7960 38517 8000
rect 38475 7951 38517 7960
rect 38859 8000 38901 8009
rect 38859 7960 38860 8000
rect 38900 7960 38901 8000
rect 38859 7951 38901 7960
rect 39243 8000 39285 8009
rect 39243 7960 39244 8000
rect 39284 7960 39285 8000
rect 39243 7951 39285 7960
rect 39627 8000 39669 8009
rect 39627 7960 39628 8000
rect 39668 7960 39669 8000
rect 39627 7951 39669 7960
rect 40011 8000 40053 8009
rect 40011 7960 40012 8000
rect 40052 7960 40053 8000
rect 40011 7951 40053 7960
rect 51051 8000 51093 8009
rect 51051 7960 51052 8000
rect 51092 7960 51093 8000
rect 51051 7951 51093 7960
rect 51435 8000 51477 8009
rect 51435 7960 51436 8000
rect 51476 7960 51477 8000
rect 51435 7951 51477 7960
rect 51819 8000 51861 8009
rect 51819 7960 51820 8000
rect 51860 7960 51861 8000
rect 51819 7951 51861 7960
rect 8187 7832 8229 7841
rect 8187 7792 8188 7832
rect 8228 7792 8229 7832
rect 8187 7783 8229 7792
rect 33147 7832 33189 7841
rect 33147 7792 33148 7832
rect 33188 7792 33189 7832
rect 33147 7783 33189 7792
rect 35451 7832 35493 7841
rect 35451 7792 35452 7832
rect 35492 7792 35493 7832
rect 35451 7783 35493 7792
rect 36987 7832 37029 7841
rect 36987 7792 36988 7832
rect 37028 7792 37029 7832
rect 36987 7783 37029 7792
rect 33531 7748 33573 7757
rect 33531 7708 33532 7748
rect 33572 7708 33573 7748
rect 33531 7699 33573 7708
rect 34683 7748 34725 7757
rect 34683 7708 34684 7748
rect 34724 7708 34725 7748
rect 34683 7699 34725 7708
rect 35835 7748 35877 7757
rect 35835 7708 35836 7748
rect 35876 7708 35877 7748
rect 35835 7699 35877 7708
rect 36603 7748 36645 7757
rect 36603 7708 36604 7748
rect 36644 7708 36645 7748
rect 36603 7699 36645 7708
rect 38619 7748 38661 7757
rect 38619 7708 38620 7748
rect 38660 7708 38661 7748
rect 38619 7699 38661 7708
rect 39003 7748 39045 7757
rect 39003 7708 39004 7748
rect 39044 7708 39045 7748
rect 39003 7699 39045 7708
rect 39771 7748 39813 7757
rect 39771 7708 39772 7748
rect 39812 7708 39813 7748
rect 39771 7699 39813 7708
rect 51675 7748 51717 7757
rect 51675 7708 51676 7748
rect 51716 7708 51717 7748
rect 51675 7699 51717 7708
rect 52059 7748 52101 7757
rect 52059 7708 52060 7748
rect 52100 7708 52101 7748
rect 52059 7699 52101 7708
rect 1152 7580 52128 7604
rect 1152 7540 4928 7580
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 5296 7540 20048 7580
rect 20088 7540 20130 7580
rect 20170 7540 20212 7580
rect 20252 7540 20294 7580
rect 20334 7540 20376 7580
rect 20416 7540 35168 7580
rect 35208 7540 35250 7580
rect 35290 7540 35332 7580
rect 35372 7540 35414 7580
rect 35454 7540 35496 7580
rect 35536 7540 50288 7580
rect 50328 7540 50370 7580
rect 50410 7540 50452 7580
rect 50492 7540 50534 7580
rect 50574 7540 50616 7580
rect 50656 7540 52128 7580
rect 1152 7516 52128 7540
rect 10875 7160 10917 7169
rect 10875 7120 10876 7160
rect 10916 7120 10917 7160
rect 10875 7111 10917 7120
rect 11115 7160 11157 7169
rect 11115 7120 11116 7160
rect 11156 7120 11157 7160
rect 11115 7111 11157 7120
rect 11499 7160 11541 7169
rect 11499 7120 11500 7160
rect 11540 7120 11541 7160
rect 11499 7111 11541 7120
rect 11979 7160 12021 7169
rect 11979 7120 11980 7160
rect 12020 7120 12021 7160
rect 11979 7111 12021 7120
rect 12651 7160 12693 7169
rect 12651 7120 12652 7160
rect 12692 7120 12693 7160
rect 12651 7111 12693 7120
rect 13611 7160 13653 7169
rect 13611 7120 13612 7160
rect 13652 7120 13653 7160
rect 13611 7111 13653 7120
rect 13995 7160 14037 7169
rect 13995 7120 13996 7160
rect 14036 7120 14037 7160
rect 13995 7111 14037 7120
rect 14859 7160 14901 7169
rect 14859 7120 14860 7160
rect 14900 7120 14901 7160
rect 14859 7111 14901 7120
rect 15003 7160 15045 7169
rect 15003 7120 15004 7160
rect 15044 7120 15045 7160
rect 15003 7111 15045 7120
rect 15243 7160 15285 7169
rect 15243 7120 15244 7160
rect 15284 7120 15285 7160
rect 15243 7111 15285 7120
rect 17163 7160 17205 7169
rect 17163 7120 17164 7160
rect 17204 7120 17205 7160
rect 17163 7111 17205 7120
rect 27051 7160 27093 7169
rect 27051 7120 27052 7160
rect 27092 7120 27093 7160
rect 27051 7111 27093 7120
rect 27435 7160 27477 7169
rect 27435 7120 27436 7160
rect 27476 7120 27477 7160
rect 27435 7111 27477 7120
rect 28779 7160 28821 7169
rect 28779 7120 28780 7160
rect 28820 7120 28821 7160
rect 28779 7111 28821 7120
rect 37371 7160 37413 7169
rect 37371 7120 37372 7160
rect 37412 7120 37413 7160
rect 37371 7111 37413 7120
rect 37659 7160 37701 7169
rect 37659 7120 37660 7160
rect 37700 7120 37701 7160
rect 37659 7111 37701 7120
rect 38091 7160 38133 7169
rect 38091 7120 38092 7160
rect 38132 7120 38133 7160
rect 38091 7111 38133 7120
rect 38907 7160 38949 7169
rect 38907 7120 38908 7160
rect 38948 7120 38949 7160
rect 38907 7111 38949 7120
rect 39082 7160 39140 7161
rect 39082 7120 39091 7160
rect 39131 7120 39140 7160
rect 39082 7119 39140 7120
rect 51435 7160 51477 7169
rect 51435 7120 51436 7160
rect 51476 7120 51477 7160
rect 51435 7111 51477 7120
rect 51819 7160 51861 7169
rect 51819 7120 51820 7160
rect 51860 7120 51861 7160
rect 51819 7111 51861 7120
rect 11259 7076 11301 7085
rect 11259 7036 11260 7076
rect 11300 7036 11301 7076
rect 11259 7027 11301 7036
rect 11739 6992 11781 7001
rect 11739 6952 11740 6992
rect 11780 6952 11781 6992
rect 11739 6943 11781 6952
rect 12411 6992 12453 7001
rect 12411 6952 12412 6992
rect 12452 6952 12453 6992
rect 12411 6943 12453 6952
rect 13371 6992 13413 7001
rect 13371 6952 13372 6992
rect 13412 6952 13413 6992
rect 13371 6943 13413 6952
rect 13755 6992 13797 7001
rect 13755 6952 13756 6992
rect 13796 6952 13797 6992
rect 13755 6943 13797 6952
rect 14619 6992 14661 7001
rect 14619 6952 14620 6992
rect 14660 6952 14661 6992
rect 14619 6943 14661 6952
rect 16923 6992 16965 7001
rect 16923 6952 16924 6992
rect 16964 6952 16965 6992
rect 16923 6943 16965 6952
rect 27291 6992 27333 7001
rect 27291 6952 27292 6992
rect 27332 6952 27333 6992
rect 27291 6943 27333 6952
rect 27675 6992 27717 7001
rect 27675 6952 27676 6992
rect 27716 6952 27717 6992
rect 27675 6943 27717 6952
rect 29019 6992 29061 7001
rect 29019 6952 29020 6992
rect 29060 6952 29061 6992
rect 29019 6943 29061 6952
rect 38331 6992 38373 7001
rect 38331 6952 38332 6992
rect 38372 6952 38373 6992
rect 38331 6943 38373 6952
rect 51675 6992 51717 7001
rect 51675 6952 51676 6992
rect 51716 6952 51717 6992
rect 51675 6943 51717 6952
rect 52059 6992 52101 7001
rect 52059 6952 52060 6992
rect 52100 6952 52101 6992
rect 52059 6943 52101 6952
rect 1152 6824 52128 6848
rect 1152 6784 3688 6824
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 4056 6784 18808 6824
rect 18848 6784 18890 6824
rect 18930 6784 18972 6824
rect 19012 6784 19054 6824
rect 19094 6784 19136 6824
rect 19176 6784 33928 6824
rect 33968 6784 34010 6824
rect 34050 6784 34092 6824
rect 34132 6784 34174 6824
rect 34214 6784 34256 6824
rect 34296 6784 49048 6824
rect 49088 6784 49130 6824
rect 49170 6784 49212 6824
rect 49252 6784 49294 6824
rect 49334 6784 49376 6824
rect 49416 6784 52128 6824
rect 1152 6760 52128 6784
rect 23451 6656 23493 6665
rect 23451 6616 23452 6656
rect 23492 6616 23493 6656
rect 23451 6607 23493 6616
rect 39867 6656 39909 6665
rect 39867 6616 39868 6656
rect 39908 6616 39909 6656
rect 39867 6607 39909 6616
rect 49563 6656 49605 6665
rect 49563 6616 49564 6656
rect 49604 6616 49605 6656
rect 49563 6607 49605 6616
rect 25851 6572 25893 6581
rect 25851 6532 25852 6572
rect 25892 6532 25893 6572
rect 25851 6523 25893 6532
rect 42555 6572 42597 6581
rect 42555 6532 42556 6572
rect 42596 6532 42597 6572
rect 42555 6523 42597 6532
rect 23211 6488 23253 6497
rect 23211 6448 23212 6488
rect 23252 6448 23253 6488
rect 23211 6439 23253 6448
rect 23595 6488 23637 6497
rect 23595 6448 23596 6488
rect 23636 6448 23637 6488
rect 23595 6439 23637 6448
rect 25035 6488 25077 6497
rect 25035 6448 25036 6488
rect 25076 6448 25077 6488
rect 25035 6439 25077 6448
rect 25275 6488 25317 6497
rect 25275 6448 25276 6488
rect 25316 6448 25317 6488
rect 25275 6439 25317 6448
rect 25611 6488 25653 6497
rect 25611 6448 25612 6488
rect 25652 6448 25653 6488
rect 25611 6439 25653 6448
rect 34827 6488 34869 6497
rect 34827 6448 34828 6488
rect 34868 6448 34869 6488
rect 34827 6439 34869 6448
rect 39627 6488 39669 6497
rect 39627 6448 39628 6488
rect 39668 6448 39669 6488
rect 39627 6439 39669 6448
rect 42315 6488 42357 6497
rect 42315 6448 42316 6488
rect 42356 6448 42357 6488
rect 42315 6439 42357 6448
rect 49323 6488 49365 6497
rect 49323 6448 49324 6488
rect 49364 6448 49365 6488
rect 49323 6439 49365 6448
rect 51435 6488 51477 6497
rect 51435 6448 51436 6488
rect 51476 6448 51477 6488
rect 51435 6439 51477 6448
rect 51819 6488 51861 6497
rect 51819 6448 51820 6488
rect 51860 6448 51861 6488
rect 51819 6439 51861 6448
rect 23835 6320 23877 6329
rect 23835 6280 23836 6320
rect 23876 6280 23877 6320
rect 23835 6271 23877 6280
rect 35067 6320 35109 6329
rect 35067 6280 35068 6320
rect 35108 6280 35109 6320
rect 35067 6271 35109 6280
rect 52059 6320 52101 6329
rect 52059 6280 52060 6320
rect 52100 6280 52101 6320
rect 52059 6271 52101 6280
rect 51675 6236 51717 6245
rect 51675 6196 51676 6236
rect 51716 6196 51717 6236
rect 51675 6187 51717 6196
rect 1152 6068 52128 6092
rect 1152 6028 4928 6068
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 5296 6028 20048 6068
rect 20088 6028 20130 6068
rect 20170 6028 20212 6068
rect 20252 6028 20294 6068
rect 20334 6028 20376 6068
rect 20416 6028 35168 6068
rect 35208 6028 35250 6068
rect 35290 6028 35332 6068
rect 35372 6028 35414 6068
rect 35454 6028 35496 6068
rect 35536 6028 50288 6068
rect 50328 6028 50370 6068
rect 50410 6028 50452 6068
rect 50492 6028 50534 6068
rect 50574 6028 50616 6068
rect 50656 6028 52128 6068
rect 1152 6004 52128 6028
rect 26763 5648 26805 5657
rect 26763 5608 26764 5648
rect 26804 5608 26805 5648
rect 26763 5599 26805 5608
rect 27627 5648 27669 5657
rect 27627 5608 27628 5648
rect 27668 5608 27669 5648
rect 27627 5599 27669 5608
rect 29835 5648 29877 5657
rect 29835 5608 29836 5648
rect 29876 5608 29877 5648
rect 29835 5599 29877 5608
rect 31659 5648 31701 5657
rect 31659 5608 31660 5648
rect 31700 5608 31701 5648
rect 31659 5599 31701 5608
rect 31899 5648 31941 5657
rect 31899 5608 31900 5648
rect 31940 5608 31941 5648
rect 31899 5599 31941 5608
rect 33099 5648 33141 5657
rect 33099 5608 33100 5648
rect 33140 5608 33141 5648
rect 33099 5599 33141 5608
rect 46443 5648 46485 5657
rect 46443 5608 46444 5648
rect 46484 5608 46485 5648
rect 46443 5599 46485 5608
rect 46683 5648 46725 5657
rect 46683 5608 46684 5648
rect 46724 5608 46725 5648
rect 46683 5599 46725 5608
rect 49227 5648 49269 5657
rect 49227 5608 49228 5648
rect 49268 5608 49269 5648
rect 49227 5599 49269 5608
rect 49467 5648 49509 5657
rect 49467 5608 49468 5648
rect 49508 5608 49509 5648
rect 49467 5599 49509 5608
rect 51435 5648 51477 5657
rect 51435 5608 51436 5648
rect 51476 5608 51477 5648
rect 51435 5599 51477 5608
rect 51819 5648 51861 5657
rect 51819 5608 51820 5648
rect 51860 5608 51861 5648
rect 51819 5599 51861 5608
rect 52059 5648 52101 5657
rect 52059 5608 52060 5648
rect 52100 5608 52101 5648
rect 52059 5599 52101 5608
rect 27003 5564 27045 5573
rect 27003 5524 27004 5564
rect 27044 5524 27045 5564
rect 27003 5515 27045 5524
rect 27867 5480 27909 5489
rect 27867 5440 27868 5480
rect 27908 5440 27909 5480
rect 27867 5431 27909 5440
rect 30075 5480 30117 5489
rect 30075 5440 30076 5480
rect 30116 5440 30117 5480
rect 30075 5431 30117 5440
rect 33339 5480 33381 5489
rect 33339 5440 33340 5480
rect 33380 5440 33381 5480
rect 33339 5431 33381 5440
rect 51675 5480 51717 5489
rect 51675 5440 51676 5480
rect 51716 5440 51717 5480
rect 51675 5431 51717 5440
rect 1152 5312 52128 5336
rect 1152 5272 3688 5312
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 4056 5272 18808 5312
rect 18848 5272 18890 5312
rect 18930 5272 18972 5312
rect 19012 5272 19054 5312
rect 19094 5272 19136 5312
rect 19176 5272 33928 5312
rect 33968 5272 34010 5312
rect 34050 5272 34092 5312
rect 34132 5272 34174 5312
rect 34214 5272 34256 5312
rect 34296 5272 49048 5312
rect 49088 5272 49130 5312
rect 49170 5272 49212 5312
rect 49252 5272 49294 5312
rect 49334 5272 49376 5312
rect 49416 5272 52128 5312
rect 1152 5248 52128 5272
rect 31995 5060 32037 5069
rect 31995 5020 31996 5060
rect 32036 5020 32037 5060
rect 31995 5011 32037 5020
rect 31755 4976 31797 4985
rect 31755 4936 31756 4976
rect 31796 4936 31797 4976
rect 31755 4927 31797 4936
rect 32427 4976 32469 4985
rect 32427 4936 32428 4976
rect 32468 4936 32469 4976
rect 32427 4927 32469 4936
rect 51435 4976 51477 4985
rect 51435 4936 51436 4976
rect 51476 4936 51477 4976
rect 51435 4927 51477 4936
rect 51819 4976 51861 4985
rect 51819 4936 51820 4976
rect 51860 4936 51861 4976
rect 51819 4927 51861 4936
rect 52059 4976 52101 4985
rect 52059 4936 52060 4976
rect 52100 4936 52101 4976
rect 52059 4927 52101 4936
rect 32667 4724 32709 4733
rect 32667 4684 32668 4724
rect 32708 4684 32709 4724
rect 32667 4675 32709 4684
rect 51675 4724 51717 4733
rect 51675 4684 51676 4724
rect 51716 4684 51717 4724
rect 51675 4675 51717 4684
rect 1152 4556 52128 4580
rect 1152 4516 4928 4556
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 5296 4516 20048 4556
rect 20088 4516 20130 4556
rect 20170 4516 20212 4556
rect 20252 4516 20294 4556
rect 20334 4516 20376 4556
rect 20416 4516 35168 4556
rect 35208 4516 35250 4556
rect 35290 4516 35332 4556
rect 35372 4516 35414 4556
rect 35454 4516 35496 4556
rect 35536 4516 50288 4556
rect 50328 4516 50370 4556
rect 50410 4516 50452 4556
rect 50492 4516 50534 4556
rect 50574 4516 50616 4556
rect 50656 4516 52128 4556
rect 1152 4492 52128 4516
rect 25467 4304 25509 4313
rect 25467 4264 25468 4304
rect 25508 4264 25509 4304
rect 25467 4255 25509 4264
rect 52059 4304 52101 4313
rect 52059 4264 52060 4304
rect 52100 4264 52101 4304
rect 52059 4255 52101 4264
rect 20619 4136 20661 4145
rect 20619 4096 20620 4136
rect 20660 4096 20661 4136
rect 20619 4087 20661 4096
rect 21675 4136 21717 4145
rect 21675 4096 21676 4136
rect 21716 4096 21717 4136
rect 21675 4087 21717 4096
rect 22059 4136 22101 4145
rect 22059 4096 22060 4136
rect 22100 4096 22101 4136
rect 22059 4087 22101 4096
rect 22539 4136 22581 4145
rect 22539 4096 22540 4136
rect 22580 4096 22581 4136
rect 22539 4087 22581 4096
rect 22923 4136 22965 4145
rect 22923 4096 22924 4136
rect 22964 4096 22965 4136
rect 22923 4087 22965 4096
rect 23307 4136 23349 4145
rect 23307 4096 23308 4136
rect 23348 4096 23349 4136
rect 23307 4087 23349 4096
rect 24075 4136 24117 4145
rect 24075 4096 24076 4136
rect 24116 4096 24117 4136
rect 24075 4087 24117 4096
rect 24459 4136 24501 4145
rect 24459 4096 24460 4136
rect 24500 4096 24501 4136
rect 24459 4087 24501 4096
rect 24843 4136 24885 4145
rect 24843 4096 24844 4136
rect 24884 4096 24885 4136
rect 24843 4087 24885 4096
rect 25227 4136 25269 4145
rect 25227 4096 25228 4136
rect 25268 4096 25269 4136
rect 25227 4087 25269 4096
rect 25611 4136 25653 4145
rect 25611 4096 25612 4136
rect 25652 4096 25653 4136
rect 25611 4087 25653 4096
rect 25995 4136 26037 4145
rect 25995 4096 25996 4136
rect 26036 4096 26037 4136
rect 25995 4087 26037 4096
rect 26235 4136 26277 4145
rect 26235 4096 26236 4136
rect 26276 4096 26277 4136
rect 26235 4087 26277 4096
rect 51435 4136 51477 4145
rect 51435 4096 51436 4136
rect 51476 4096 51477 4136
rect 51435 4087 51477 4096
rect 51819 4136 51861 4145
rect 51819 4096 51820 4136
rect 51860 4096 51861 4136
rect 51819 4087 51861 4096
rect 22299 4052 22341 4061
rect 22299 4012 22300 4052
rect 22340 4012 22341 4052
rect 22299 4003 22341 4012
rect 25083 4052 25125 4061
rect 25083 4012 25084 4052
rect 25124 4012 25125 4052
rect 25083 4003 25125 4012
rect 51675 4052 51717 4061
rect 51675 4012 51676 4052
rect 51716 4012 51717 4052
rect 51675 4003 51717 4012
rect 20859 3968 20901 3977
rect 20859 3928 20860 3968
rect 20900 3928 20901 3968
rect 20859 3919 20901 3928
rect 21915 3968 21957 3977
rect 21915 3928 21916 3968
rect 21956 3928 21957 3968
rect 21915 3919 21957 3928
rect 22779 3968 22821 3977
rect 22779 3928 22780 3968
rect 22820 3928 22821 3968
rect 22779 3919 22821 3928
rect 23163 3968 23205 3977
rect 23163 3928 23164 3968
rect 23204 3928 23205 3968
rect 23163 3919 23205 3928
rect 23547 3968 23589 3977
rect 23547 3928 23548 3968
rect 23588 3928 23589 3968
rect 23547 3919 23589 3928
rect 24315 3968 24357 3977
rect 24315 3928 24316 3968
rect 24356 3928 24357 3968
rect 24315 3919 24357 3928
rect 24699 3968 24741 3977
rect 24699 3928 24700 3968
rect 24740 3928 24741 3968
rect 24699 3919 24741 3928
rect 25851 3968 25893 3977
rect 25851 3928 25852 3968
rect 25892 3928 25893 3968
rect 25851 3919 25893 3928
rect 1152 3800 52128 3824
rect 1152 3760 3688 3800
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 4056 3760 18808 3800
rect 18848 3760 18890 3800
rect 18930 3760 18972 3800
rect 19012 3760 19054 3800
rect 19094 3760 19136 3800
rect 19176 3760 33928 3800
rect 33968 3760 34010 3800
rect 34050 3760 34092 3800
rect 34132 3760 34174 3800
rect 34214 3760 34256 3800
rect 34296 3760 49048 3800
rect 49088 3760 49130 3800
rect 49170 3760 49212 3800
rect 49252 3760 49294 3800
rect 49334 3760 49376 3800
rect 49416 3760 52128 3800
rect 1152 3736 52128 3760
rect 22011 3632 22053 3641
rect 22011 3592 22012 3632
rect 22052 3592 22053 3632
rect 22011 3583 22053 3592
rect 23355 3632 23397 3641
rect 23355 3592 23356 3632
rect 23396 3592 23397 3632
rect 23355 3583 23397 3592
rect 24507 3632 24549 3641
rect 24507 3592 24508 3632
rect 24548 3592 24549 3632
rect 24507 3583 24549 3592
rect 25467 3632 25509 3641
rect 25467 3592 25468 3632
rect 25508 3592 25509 3632
rect 25467 3583 25509 3592
rect 28539 3632 28581 3641
rect 28539 3592 28540 3632
rect 28580 3592 28581 3632
rect 28539 3583 28581 3592
rect 52059 3632 52101 3641
rect 52059 3592 52060 3632
rect 52100 3592 52101 3632
rect 52059 3583 52101 3592
rect 21771 3464 21813 3473
rect 21771 3424 21772 3464
rect 21812 3424 21813 3464
rect 21771 3415 21813 3424
rect 23115 3464 23157 3473
rect 23115 3424 23116 3464
rect 23156 3424 23157 3464
rect 23115 3415 23157 3424
rect 24267 3464 24309 3473
rect 24267 3424 24268 3464
rect 24308 3424 24309 3464
rect 24267 3415 24309 3424
rect 24843 3464 24885 3473
rect 24843 3424 24844 3464
rect 24884 3424 24885 3464
rect 24843 3415 24885 3424
rect 25227 3464 25269 3473
rect 25227 3424 25228 3464
rect 25268 3424 25269 3464
rect 25227 3415 25269 3424
rect 28299 3464 28341 3473
rect 28299 3424 28300 3464
rect 28340 3424 28341 3464
rect 28299 3415 28341 3424
rect 51435 3464 51477 3473
rect 51435 3424 51436 3464
rect 51476 3424 51477 3464
rect 51435 3415 51477 3424
rect 51819 3464 51861 3473
rect 51819 3424 51820 3464
rect 51860 3424 51861 3464
rect 51819 3415 51861 3424
rect 51675 3296 51717 3305
rect 51675 3256 51676 3296
rect 51716 3256 51717 3296
rect 51675 3247 51717 3256
rect 25083 3212 25125 3221
rect 25083 3172 25084 3212
rect 25124 3172 25125 3212
rect 25083 3163 25125 3172
rect 1152 3044 52128 3068
rect 1152 3004 4928 3044
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 5296 3004 20048 3044
rect 20088 3004 20130 3044
rect 20170 3004 20212 3044
rect 20252 3004 20294 3044
rect 20334 3004 20376 3044
rect 20416 3004 35168 3044
rect 35208 3004 35250 3044
rect 35290 3004 35332 3044
rect 35372 3004 35414 3044
rect 35454 3004 35496 3044
rect 35536 3004 50288 3044
rect 50328 3004 50370 3044
rect 50410 3004 50452 3044
rect 50492 3004 50534 3044
rect 50574 3004 50616 3044
rect 50656 3004 52128 3044
rect 1152 2980 52128 3004
rect 25467 2876 25509 2885
rect 25467 2836 25468 2876
rect 25508 2836 25509 2876
rect 25467 2827 25509 2836
rect 52059 2876 52101 2885
rect 52059 2836 52060 2876
rect 52100 2836 52101 2876
rect 52059 2827 52101 2836
rect 25227 2624 25269 2633
rect 25227 2584 25228 2624
rect 25268 2584 25269 2624
rect 25227 2575 25269 2584
rect 51051 2624 51093 2633
rect 51051 2584 51052 2624
rect 51092 2584 51093 2624
rect 51051 2575 51093 2584
rect 51435 2624 51477 2633
rect 51435 2584 51436 2624
rect 51476 2584 51477 2624
rect 51435 2575 51477 2584
rect 51819 2624 51861 2633
rect 51819 2584 51820 2624
rect 51860 2584 51861 2624
rect 51819 2575 51861 2584
rect 51675 2540 51717 2549
rect 51675 2500 51676 2540
rect 51716 2500 51717 2540
rect 51675 2491 51717 2500
rect 51291 2456 51333 2465
rect 51291 2416 51292 2456
rect 51332 2416 51333 2456
rect 51291 2407 51333 2416
rect 1152 2288 52128 2312
rect 1152 2248 3688 2288
rect 3728 2248 3770 2288
rect 3810 2248 3852 2288
rect 3892 2248 3934 2288
rect 3974 2248 4016 2288
rect 4056 2248 18808 2288
rect 18848 2248 18890 2288
rect 18930 2248 18972 2288
rect 19012 2248 19054 2288
rect 19094 2248 19136 2288
rect 19176 2248 33928 2288
rect 33968 2248 34010 2288
rect 34050 2248 34092 2288
rect 34132 2248 34174 2288
rect 34214 2248 34256 2288
rect 34296 2248 49048 2288
rect 49088 2248 49130 2288
rect 49170 2248 49212 2288
rect 49252 2248 49294 2288
rect 49334 2248 49376 2288
rect 49416 2248 52128 2288
rect 1152 2224 52128 2248
rect 52059 2120 52101 2129
rect 52059 2080 52060 2120
rect 52100 2080 52101 2120
rect 52059 2071 52101 2080
rect 50314 1952 50372 1953
rect 50314 1912 50323 1952
rect 50363 1912 50372 1952
rect 50314 1911 50372 1912
rect 50667 1952 50709 1961
rect 50667 1912 50668 1952
rect 50708 1912 50709 1952
rect 50667 1903 50709 1912
rect 51051 1952 51093 1961
rect 51051 1912 51052 1952
rect 51092 1912 51093 1952
rect 51051 1903 51093 1912
rect 51291 1952 51333 1961
rect 51291 1912 51292 1952
rect 51332 1912 51333 1952
rect 51291 1903 51333 1912
rect 51435 1952 51477 1961
rect 51435 1912 51436 1952
rect 51476 1912 51477 1952
rect 51435 1903 51477 1912
rect 51819 1952 51861 1961
rect 51819 1912 51820 1952
rect 51860 1912 51861 1952
rect 51819 1903 51861 1912
rect 50907 1784 50949 1793
rect 50907 1744 50908 1784
rect 50948 1744 50949 1784
rect 50907 1735 50949 1744
rect 50523 1700 50565 1709
rect 50523 1660 50524 1700
rect 50564 1660 50565 1700
rect 50523 1651 50565 1660
rect 51675 1700 51717 1709
rect 51675 1660 51676 1700
rect 51716 1660 51717 1700
rect 51675 1651 51717 1660
rect 1152 1532 52128 1556
rect 1152 1492 4928 1532
rect 4968 1492 5010 1532
rect 5050 1492 5092 1532
rect 5132 1492 5174 1532
rect 5214 1492 5256 1532
rect 5296 1492 20048 1532
rect 20088 1492 20130 1532
rect 20170 1492 20212 1532
rect 20252 1492 20294 1532
rect 20334 1492 20376 1532
rect 20416 1492 35168 1532
rect 35208 1492 35250 1532
rect 35290 1492 35332 1532
rect 35372 1492 35414 1532
rect 35454 1492 35496 1532
rect 35536 1492 50288 1532
rect 50328 1492 50370 1532
rect 50410 1492 50452 1532
rect 50492 1492 50534 1532
rect 50574 1492 50616 1532
rect 50656 1492 52128 1532
rect 1152 1468 52128 1492
<< via1 >>
rect 3688 9808 3728 9848
rect 3770 9808 3810 9848
rect 3852 9808 3892 9848
rect 3934 9808 3974 9848
rect 4016 9808 4056 9848
rect 18808 9808 18848 9848
rect 18890 9808 18930 9848
rect 18972 9808 19012 9848
rect 19054 9808 19094 9848
rect 19136 9808 19176 9848
rect 33928 9808 33968 9848
rect 34010 9808 34050 9848
rect 34092 9808 34132 9848
rect 34174 9808 34214 9848
rect 34256 9808 34296 9848
rect 49048 9808 49088 9848
rect 49130 9808 49170 9848
rect 49212 9808 49252 9848
rect 49294 9808 49334 9848
rect 49376 9808 49416 9848
rect 2812 9640 2852 9680
rect 3196 9640 3236 9680
rect 3580 9640 3620 9680
rect 3964 9640 4004 9680
rect 4348 9640 4388 9680
rect 4732 9640 4772 9680
rect 5116 9640 5156 9680
rect 5500 9640 5540 9680
rect 5884 9640 5924 9680
rect 6268 9640 6308 9680
rect 6652 9640 6692 9680
rect 7036 9640 7076 9680
rect 7420 9640 7460 9680
rect 7804 9640 7844 9680
rect 8188 9640 8228 9680
rect 8572 9640 8612 9680
rect 8956 9640 8996 9680
rect 9340 9640 9380 9680
rect 9724 9640 9764 9680
rect 10108 9640 10148 9680
rect 10492 9640 10532 9680
rect 10876 9640 10916 9680
rect 11260 9640 11300 9680
rect 11644 9640 11684 9680
rect 12028 9640 12068 9680
rect 12412 9640 12452 9680
rect 12796 9640 12836 9680
rect 13180 9640 13220 9680
rect 13564 9640 13604 9680
rect 13948 9640 13988 9680
rect 14332 9640 14372 9680
rect 14716 9640 14756 9680
rect 15100 9640 15140 9680
rect 15484 9640 15524 9680
rect 15868 9640 15908 9680
rect 16252 9640 16292 9680
rect 16636 9640 16676 9680
rect 17020 9640 17060 9680
rect 17404 9640 17444 9680
rect 17788 9640 17828 9680
rect 18172 9640 18212 9680
rect 18556 9640 18596 9680
rect 19324 9640 19364 9680
rect 19708 9640 19748 9680
rect 20092 9640 20132 9680
rect 20476 9640 20516 9680
rect 20860 9640 20900 9680
rect 21244 9640 21284 9680
rect 21628 9640 21668 9680
rect 22012 9640 22052 9680
rect 22396 9640 22436 9680
rect 42748 9640 42788 9680
rect 43132 9640 43172 9680
rect 43516 9640 43556 9680
rect 43900 9640 43940 9680
rect 44284 9640 44324 9680
rect 44668 9640 44708 9680
rect 45052 9640 45092 9680
rect 45436 9640 45476 9680
rect 45820 9640 45860 9680
rect 46204 9640 46244 9680
rect 46588 9640 46628 9680
rect 46972 9640 47012 9680
rect 47356 9640 47396 9680
rect 47740 9640 47780 9680
rect 48124 9640 48164 9680
rect 48508 9640 48548 9680
rect 48892 9640 48932 9680
rect 49276 9640 49316 9680
rect 50044 9640 50084 9680
rect 50428 9640 50468 9680
rect 18940 9556 18980 9596
rect 49660 9556 49700 9596
rect 3052 9472 3092 9512
rect 3436 9472 3476 9512
rect 3820 9472 3860 9512
rect 4204 9472 4244 9512
rect 4588 9472 4628 9512
rect 4972 9472 5012 9512
rect 5356 9472 5396 9512
rect 5740 9472 5780 9512
rect 6124 9472 6164 9512
rect 6508 9472 6548 9512
rect 6892 9472 6932 9512
rect 7276 9472 7316 9512
rect 7660 9472 7700 9512
rect 8044 9472 8084 9512
rect 8428 9472 8468 9512
rect 8812 9472 8852 9512
rect 9196 9472 9236 9512
rect 9580 9472 9620 9512
rect 9964 9472 10004 9512
rect 10348 9472 10388 9512
rect 10732 9472 10772 9512
rect 11116 9472 11156 9512
rect 11500 9472 11540 9512
rect 11884 9472 11924 9512
rect 12268 9472 12308 9512
rect 12652 9472 12692 9512
rect 13036 9472 13076 9512
rect 13420 9472 13460 9512
rect 13804 9472 13844 9512
rect 14188 9472 14228 9512
rect 14572 9472 14612 9512
rect 14956 9472 14996 9512
rect 15340 9472 15380 9512
rect 15724 9472 15764 9512
rect 16108 9472 16148 9512
rect 16492 9472 16532 9512
rect 16876 9472 16916 9512
rect 17260 9472 17300 9512
rect 17644 9472 17684 9512
rect 18028 9472 18068 9512
rect 18412 9472 18452 9512
rect 18796 9472 18836 9512
rect 19180 9472 19220 9512
rect 19564 9472 19604 9512
rect 19948 9472 19988 9512
rect 20332 9472 20372 9512
rect 20716 9472 20756 9512
rect 21100 9472 21140 9512
rect 21484 9472 21524 9512
rect 21868 9472 21908 9512
rect 22252 9472 22292 9512
rect 22636 9472 22676 9512
rect 42988 9472 43028 9512
rect 43372 9472 43412 9512
rect 43756 9472 43796 9512
rect 44140 9472 44180 9512
rect 44524 9472 44564 9512
rect 44908 9472 44948 9512
rect 45292 9472 45332 9512
rect 45676 9472 45716 9512
rect 46060 9472 46100 9512
rect 46444 9472 46484 9512
rect 46828 9472 46868 9512
rect 47212 9472 47252 9512
rect 47596 9472 47636 9512
rect 47980 9472 48020 9512
rect 48364 9472 48404 9512
rect 48748 9472 48788 9512
rect 49132 9472 49172 9512
rect 49516 9472 49556 9512
rect 49900 9472 49940 9512
rect 50284 9472 50324 9512
rect 50668 9472 50708 9512
rect 51052 9472 51092 9512
rect 51436 9472 51476 9512
rect 51820 9472 51860 9512
rect 51292 9304 51332 9344
rect 51676 9220 51716 9260
rect 52060 9220 52100 9260
rect 4928 9052 4968 9092
rect 5010 9052 5050 9092
rect 5092 9052 5132 9092
rect 5174 9052 5214 9092
rect 5256 9052 5296 9092
rect 20048 9052 20088 9092
rect 20130 9052 20170 9092
rect 20212 9052 20252 9092
rect 20294 9052 20334 9092
rect 20376 9052 20416 9092
rect 35168 9052 35208 9092
rect 35250 9052 35290 9092
rect 35332 9052 35372 9092
rect 35414 9052 35454 9092
rect 35496 9052 35536 9092
rect 50288 9052 50328 9092
rect 50370 9052 50410 9092
rect 50452 9052 50492 9092
rect 50534 9052 50574 9092
rect 50616 9052 50656 9092
rect 21628 8884 21668 8924
rect 23068 8884 23108 8924
rect 23644 8884 23684 8924
rect 27004 8884 27044 8924
rect 28156 8884 28196 8924
rect 28924 8884 28964 8924
rect 29692 8884 29732 8924
rect 50140 8884 50180 8924
rect 50524 8884 50564 8924
rect 50908 8884 50948 8924
rect 51292 8884 51332 8924
rect 29308 8800 29348 8840
rect 21868 8632 21908 8672
rect 22348 8632 22388 8672
rect 22732 8632 22772 8672
rect 23308 8632 23348 8672
rect 23884 8632 23924 8672
rect 26764 8632 26804 8672
rect 27148 8632 27188 8672
rect 27532 8632 27572 8672
rect 27772 8632 27812 8672
rect 27955 8632 27995 8672
rect 28300 8632 28340 8672
rect 28540 8632 28580 8672
rect 28684 8632 28724 8672
rect 29068 8632 29108 8672
rect 29452 8632 29492 8672
rect 31228 8632 31268 8672
rect 31468 8632 31508 8672
rect 49900 8632 49940 8672
rect 50284 8632 50324 8672
rect 50668 8632 50708 8672
rect 51052 8632 51092 8672
rect 51436 8632 51476 8672
rect 51820 8632 51860 8672
rect 27388 8548 27428 8588
rect 22108 8464 22148 8504
rect 22492 8464 22532 8504
rect 51676 8464 51716 8504
rect 52060 8464 52100 8504
rect 3688 8296 3728 8336
rect 3770 8296 3810 8336
rect 3852 8296 3892 8336
rect 3934 8296 3974 8336
rect 4016 8296 4056 8336
rect 18808 8296 18848 8336
rect 18890 8296 18930 8336
rect 18972 8296 19012 8336
rect 19054 8296 19094 8336
rect 19136 8296 19176 8336
rect 33928 8296 33968 8336
rect 34010 8296 34050 8336
rect 34092 8296 34132 8336
rect 34174 8296 34214 8336
rect 34256 8296 34296 8336
rect 49048 8296 49088 8336
rect 49130 8296 49170 8336
rect 49212 8296 49252 8336
rect 49294 8296 49334 8336
rect 49376 8296 49416 8336
rect 3484 8128 3524 8168
rect 4348 8128 4388 8168
rect 6364 8128 6404 8168
rect 7804 8128 7844 8168
rect 10204 8128 10244 8168
rect 15292 8128 15332 8168
rect 15676 8128 15716 8168
rect 16060 8128 16100 8168
rect 16444 8128 16484 8168
rect 16828 8128 16868 8168
rect 17596 8128 17636 8168
rect 17980 8128 18020 8168
rect 18364 8128 18404 8168
rect 19036 8128 19076 8168
rect 20764 8128 20804 8168
rect 32764 8128 32804 8168
rect 37084 8128 37124 8168
rect 37468 8128 37508 8168
rect 38140 8128 38180 8168
rect 51292 8128 51332 8168
rect 5500 8044 5540 8084
rect 11932 8044 11972 8084
rect 17212 8044 17252 8084
rect 19420 8044 19460 8084
rect 20284 8044 20324 8084
rect 28636 8044 28676 8084
rect 35068 8044 35108 8084
rect 39388 8044 39428 8084
rect 3244 7960 3284 8000
rect 4588 7960 4628 8000
rect 5260 7960 5300 8000
rect 6124 7960 6164 8000
rect 8044 7960 8084 8000
rect 8428 7960 8468 8000
rect 10444 7960 10484 8000
rect 10588 7960 10628 8000
rect 10828 7960 10868 8000
rect 12172 7960 12212 8000
rect 15532 7960 15572 8000
rect 15916 7960 15956 8000
rect 16300 7960 16340 8000
rect 16684 7960 16724 8000
rect 17068 7960 17108 8000
rect 17452 7960 17492 8000
rect 17836 7960 17876 8000
rect 18220 7960 18260 8000
rect 18604 7960 18644 8000
rect 19276 7960 19316 8000
rect 19660 7960 19700 8000
rect 20524 7960 20564 8000
rect 21004 7960 21044 8000
rect 28396 7960 28436 8000
rect 33004 7960 33044 8000
rect 33388 7960 33428 8000
rect 33772 7960 33812 8000
rect 34924 7960 34964 8000
rect 35308 7960 35348 8000
rect 35692 7960 35732 8000
rect 36076 7960 36116 8000
rect 36364 7960 36404 8000
rect 36748 7960 36788 8000
rect 37324 7960 37364 8000
rect 37708 7960 37748 8000
rect 37900 7960 37940 8000
rect 38236 7960 38276 8000
rect 38476 7960 38516 8000
rect 38860 7960 38900 8000
rect 39244 7960 39284 8000
rect 39628 7960 39668 8000
rect 40012 7960 40052 8000
rect 51052 7960 51092 8000
rect 51436 7960 51476 8000
rect 51820 7960 51860 8000
rect 8188 7792 8228 7832
rect 33148 7792 33188 7832
rect 35452 7792 35492 7832
rect 36988 7792 37028 7832
rect 33532 7708 33572 7748
rect 34684 7708 34724 7748
rect 35836 7708 35876 7748
rect 36604 7708 36644 7748
rect 38620 7708 38660 7748
rect 39004 7708 39044 7748
rect 39772 7708 39812 7748
rect 51676 7708 51716 7748
rect 52060 7708 52100 7748
rect 4928 7540 4968 7580
rect 5010 7540 5050 7580
rect 5092 7540 5132 7580
rect 5174 7540 5214 7580
rect 5256 7540 5296 7580
rect 20048 7540 20088 7580
rect 20130 7540 20170 7580
rect 20212 7540 20252 7580
rect 20294 7540 20334 7580
rect 20376 7540 20416 7580
rect 35168 7540 35208 7580
rect 35250 7540 35290 7580
rect 35332 7540 35372 7580
rect 35414 7540 35454 7580
rect 35496 7540 35536 7580
rect 50288 7540 50328 7580
rect 50370 7540 50410 7580
rect 50452 7540 50492 7580
rect 50534 7540 50574 7580
rect 50616 7540 50656 7580
rect 10876 7120 10916 7160
rect 11116 7120 11156 7160
rect 11500 7120 11540 7160
rect 11980 7120 12020 7160
rect 12652 7120 12692 7160
rect 13612 7120 13652 7160
rect 13996 7120 14036 7160
rect 14860 7120 14900 7160
rect 15004 7120 15044 7160
rect 15244 7120 15284 7160
rect 17164 7120 17204 7160
rect 27052 7120 27092 7160
rect 27436 7120 27476 7160
rect 28780 7120 28820 7160
rect 37372 7120 37412 7160
rect 37660 7120 37700 7160
rect 38092 7120 38132 7160
rect 38908 7120 38948 7160
rect 39091 7120 39131 7160
rect 51436 7120 51476 7160
rect 51820 7120 51860 7160
rect 11260 7036 11300 7076
rect 11740 6952 11780 6992
rect 12412 6952 12452 6992
rect 13372 6952 13412 6992
rect 13756 6952 13796 6992
rect 14620 6952 14660 6992
rect 16924 6952 16964 6992
rect 27292 6952 27332 6992
rect 27676 6952 27716 6992
rect 29020 6952 29060 6992
rect 38332 6952 38372 6992
rect 51676 6952 51716 6992
rect 52060 6952 52100 6992
rect 3688 6784 3728 6824
rect 3770 6784 3810 6824
rect 3852 6784 3892 6824
rect 3934 6784 3974 6824
rect 4016 6784 4056 6824
rect 18808 6784 18848 6824
rect 18890 6784 18930 6824
rect 18972 6784 19012 6824
rect 19054 6784 19094 6824
rect 19136 6784 19176 6824
rect 33928 6784 33968 6824
rect 34010 6784 34050 6824
rect 34092 6784 34132 6824
rect 34174 6784 34214 6824
rect 34256 6784 34296 6824
rect 49048 6784 49088 6824
rect 49130 6784 49170 6824
rect 49212 6784 49252 6824
rect 49294 6784 49334 6824
rect 49376 6784 49416 6824
rect 23452 6616 23492 6656
rect 39868 6616 39908 6656
rect 49564 6616 49604 6656
rect 25852 6532 25892 6572
rect 42556 6532 42596 6572
rect 23212 6448 23252 6488
rect 23596 6448 23636 6488
rect 25036 6448 25076 6488
rect 25276 6448 25316 6488
rect 25612 6448 25652 6488
rect 34828 6448 34868 6488
rect 39628 6448 39668 6488
rect 42316 6448 42356 6488
rect 49324 6448 49364 6488
rect 51436 6448 51476 6488
rect 51820 6448 51860 6488
rect 23836 6280 23876 6320
rect 35068 6280 35108 6320
rect 52060 6280 52100 6320
rect 51676 6196 51716 6236
rect 4928 6028 4968 6068
rect 5010 6028 5050 6068
rect 5092 6028 5132 6068
rect 5174 6028 5214 6068
rect 5256 6028 5296 6068
rect 20048 6028 20088 6068
rect 20130 6028 20170 6068
rect 20212 6028 20252 6068
rect 20294 6028 20334 6068
rect 20376 6028 20416 6068
rect 35168 6028 35208 6068
rect 35250 6028 35290 6068
rect 35332 6028 35372 6068
rect 35414 6028 35454 6068
rect 35496 6028 35536 6068
rect 50288 6028 50328 6068
rect 50370 6028 50410 6068
rect 50452 6028 50492 6068
rect 50534 6028 50574 6068
rect 50616 6028 50656 6068
rect 26764 5608 26804 5648
rect 27628 5608 27668 5648
rect 29836 5608 29876 5648
rect 31660 5608 31700 5648
rect 31900 5608 31940 5648
rect 33100 5608 33140 5648
rect 46444 5608 46484 5648
rect 46684 5608 46724 5648
rect 49228 5608 49268 5648
rect 49468 5608 49508 5648
rect 51436 5608 51476 5648
rect 51820 5608 51860 5648
rect 52060 5608 52100 5648
rect 27004 5524 27044 5564
rect 27868 5440 27908 5480
rect 30076 5440 30116 5480
rect 33340 5440 33380 5480
rect 51676 5440 51716 5480
rect 3688 5272 3728 5312
rect 3770 5272 3810 5312
rect 3852 5272 3892 5312
rect 3934 5272 3974 5312
rect 4016 5272 4056 5312
rect 18808 5272 18848 5312
rect 18890 5272 18930 5312
rect 18972 5272 19012 5312
rect 19054 5272 19094 5312
rect 19136 5272 19176 5312
rect 33928 5272 33968 5312
rect 34010 5272 34050 5312
rect 34092 5272 34132 5312
rect 34174 5272 34214 5312
rect 34256 5272 34296 5312
rect 49048 5272 49088 5312
rect 49130 5272 49170 5312
rect 49212 5272 49252 5312
rect 49294 5272 49334 5312
rect 49376 5272 49416 5312
rect 31996 5020 32036 5060
rect 31756 4936 31796 4976
rect 32428 4936 32468 4976
rect 51436 4936 51476 4976
rect 51820 4936 51860 4976
rect 52060 4936 52100 4976
rect 32668 4684 32708 4724
rect 51676 4684 51716 4724
rect 4928 4516 4968 4556
rect 5010 4516 5050 4556
rect 5092 4516 5132 4556
rect 5174 4516 5214 4556
rect 5256 4516 5296 4556
rect 20048 4516 20088 4556
rect 20130 4516 20170 4556
rect 20212 4516 20252 4556
rect 20294 4516 20334 4556
rect 20376 4516 20416 4556
rect 35168 4516 35208 4556
rect 35250 4516 35290 4556
rect 35332 4516 35372 4556
rect 35414 4516 35454 4556
rect 35496 4516 35536 4556
rect 50288 4516 50328 4556
rect 50370 4516 50410 4556
rect 50452 4516 50492 4556
rect 50534 4516 50574 4556
rect 50616 4516 50656 4556
rect 25468 4264 25508 4304
rect 52060 4264 52100 4304
rect 20620 4096 20660 4136
rect 21676 4096 21716 4136
rect 22060 4096 22100 4136
rect 22540 4096 22580 4136
rect 22924 4096 22964 4136
rect 23308 4096 23348 4136
rect 24076 4096 24116 4136
rect 24460 4096 24500 4136
rect 24844 4096 24884 4136
rect 25228 4096 25268 4136
rect 25612 4096 25652 4136
rect 25996 4096 26036 4136
rect 26236 4096 26276 4136
rect 51436 4096 51476 4136
rect 51820 4096 51860 4136
rect 22300 4012 22340 4052
rect 25084 4012 25124 4052
rect 51676 4012 51716 4052
rect 20860 3928 20900 3968
rect 21916 3928 21956 3968
rect 22780 3928 22820 3968
rect 23164 3928 23204 3968
rect 23548 3928 23588 3968
rect 24316 3928 24356 3968
rect 24700 3928 24740 3968
rect 25852 3928 25892 3968
rect 3688 3760 3728 3800
rect 3770 3760 3810 3800
rect 3852 3760 3892 3800
rect 3934 3760 3974 3800
rect 4016 3760 4056 3800
rect 18808 3760 18848 3800
rect 18890 3760 18930 3800
rect 18972 3760 19012 3800
rect 19054 3760 19094 3800
rect 19136 3760 19176 3800
rect 33928 3760 33968 3800
rect 34010 3760 34050 3800
rect 34092 3760 34132 3800
rect 34174 3760 34214 3800
rect 34256 3760 34296 3800
rect 49048 3760 49088 3800
rect 49130 3760 49170 3800
rect 49212 3760 49252 3800
rect 49294 3760 49334 3800
rect 49376 3760 49416 3800
rect 22012 3592 22052 3632
rect 23356 3592 23396 3632
rect 24508 3592 24548 3632
rect 25468 3592 25508 3632
rect 28540 3592 28580 3632
rect 52060 3592 52100 3632
rect 21772 3424 21812 3464
rect 23116 3424 23156 3464
rect 24268 3424 24308 3464
rect 24844 3424 24884 3464
rect 25228 3424 25268 3464
rect 28300 3424 28340 3464
rect 51436 3424 51476 3464
rect 51820 3424 51860 3464
rect 51676 3256 51716 3296
rect 25084 3172 25124 3212
rect 4928 3004 4968 3044
rect 5010 3004 5050 3044
rect 5092 3004 5132 3044
rect 5174 3004 5214 3044
rect 5256 3004 5296 3044
rect 20048 3004 20088 3044
rect 20130 3004 20170 3044
rect 20212 3004 20252 3044
rect 20294 3004 20334 3044
rect 20376 3004 20416 3044
rect 35168 3004 35208 3044
rect 35250 3004 35290 3044
rect 35332 3004 35372 3044
rect 35414 3004 35454 3044
rect 35496 3004 35536 3044
rect 50288 3004 50328 3044
rect 50370 3004 50410 3044
rect 50452 3004 50492 3044
rect 50534 3004 50574 3044
rect 50616 3004 50656 3044
rect 25468 2836 25508 2876
rect 52060 2836 52100 2876
rect 25228 2584 25268 2624
rect 51052 2584 51092 2624
rect 51436 2584 51476 2624
rect 51820 2584 51860 2624
rect 51676 2500 51716 2540
rect 51292 2416 51332 2456
rect 3688 2248 3728 2288
rect 3770 2248 3810 2288
rect 3852 2248 3892 2288
rect 3934 2248 3974 2288
rect 4016 2248 4056 2288
rect 18808 2248 18848 2288
rect 18890 2248 18930 2288
rect 18972 2248 19012 2288
rect 19054 2248 19094 2288
rect 19136 2248 19176 2288
rect 33928 2248 33968 2288
rect 34010 2248 34050 2288
rect 34092 2248 34132 2288
rect 34174 2248 34214 2288
rect 34256 2248 34296 2288
rect 49048 2248 49088 2288
rect 49130 2248 49170 2288
rect 49212 2248 49252 2288
rect 49294 2248 49334 2288
rect 49376 2248 49416 2288
rect 52060 2080 52100 2120
rect 50323 1912 50363 1952
rect 50668 1912 50708 1952
rect 51052 1912 51092 1952
rect 51292 1912 51332 1952
rect 51436 1912 51476 1952
rect 51820 1912 51860 1952
rect 50908 1744 50948 1784
rect 50524 1660 50564 1700
rect 51676 1660 51716 1700
rect 4928 1492 4968 1532
rect 5010 1492 5050 1532
rect 5092 1492 5132 1532
rect 5174 1492 5214 1532
rect 5256 1492 5296 1532
rect 20048 1492 20088 1532
rect 20130 1492 20170 1532
rect 20212 1492 20252 1532
rect 20294 1492 20334 1532
rect 20376 1492 20416 1532
rect 35168 1492 35208 1532
rect 35250 1492 35290 1532
rect 35332 1492 35372 1532
rect 35414 1492 35454 1532
rect 35496 1492 35536 1532
rect 50288 1492 50328 1532
rect 50370 1492 50410 1532
rect 50452 1492 50492 1532
rect 50534 1492 50574 1532
rect 50616 1492 50656 1532
<< metal2 >>
rect 17155 11740 17164 11780
rect 17204 11740 31948 11780
rect 31988 11740 31997 11780
rect 17251 11656 17260 11696
rect 17300 11656 31564 11696
rect 31604 11656 31613 11696
rect 19363 11572 19372 11612
rect 19412 11572 32716 11612
rect 32756 11572 32765 11612
rect 19555 11488 19564 11528
rect 19604 11488 31180 11528
rect 31220 11488 31229 11528
rect 19843 11404 19852 11444
rect 19892 11404 30796 11444
rect 30836 11404 30845 11444
rect 16675 11152 16684 11192
rect 16724 11152 25036 11192
rect 25076 11152 25085 11192
rect 0 11024 90 11044
rect 53190 11024 53280 11044
rect 0 10984 748 11024
rect 788 10984 797 11024
rect 50851 10984 50860 11024
rect 50900 10984 53280 11024
rect 0 10964 90 10984
rect 53190 10964 53280 10984
rect 0 10688 90 10708
rect 53190 10688 53280 10708
rect 0 10648 556 10688
rect 596 10648 605 10688
rect 50755 10648 50764 10688
rect 50804 10648 53280 10688
rect 0 10628 90 10648
rect 53190 10628 53280 10648
rect 0 10352 90 10372
rect 53190 10352 53280 10372
rect 0 10312 1228 10352
rect 1268 10312 1277 10352
rect 52291 10312 52300 10352
rect 52340 10312 53280 10352
rect 0 10292 90 10312
rect 53190 10292 53280 10312
rect 18019 10228 18028 10268
rect 18068 10228 24652 10268
rect 24692 10228 24701 10268
rect 22828 10144 23116 10184
rect 23156 10144 23165 10184
rect 22828 10100 22868 10144
rect 10732 10060 22868 10100
rect 23299 10060 23308 10100
rect 23348 10060 35788 10100
rect 35828 10060 35837 10100
rect 0 10016 90 10036
rect 0 9976 1420 10016
rect 1460 9976 1469 10016
rect 1996 9976 8620 10016
rect 8660 9976 8669 10016
rect 0 9956 90 9976
rect 0 9680 90 9700
rect 1996 9680 2036 9976
rect 3679 9808 3688 9848
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 4056 9808 4065 9848
rect 3052 9724 10636 9764
rect 10676 9724 10685 9764
rect 0 9640 2036 9680
rect 2755 9640 2764 9680
rect 2804 9640 2812 9680
rect 2852 9640 2935 9680
rect 0 9620 90 9640
rect 3052 9512 3092 9724
rect 3139 9640 3148 9680
rect 3188 9640 3196 9680
rect 3236 9640 3319 9680
rect 3523 9640 3532 9680
rect 3572 9640 3580 9680
rect 3620 9640 3703 9680
rect 3955 9640 3964 9680
rect 4004 9640 4108 9680
rect 4148 9640 4157 9680
rect 4291 9640 4300 9680
rect 4340 9640 4348 9680
rect 4388 9640 4471 9680
rect 4675 9640 4684 9680
rect 4724 9640 4732 9680
rect 4772 9640 4855 9680
rect 5059 9640 5068 9680
rect 5108 9640 5116 9680
rect 5156 9640 5239 9680
rect 5443 9640 5452 9680
rect 5492 9640 5500 9680
rect 5540 9640 5623 9680
rect 5827 9640 5836 9680
rect 5876 9640 5884 9680
rect 5924 9640 6007 9680
rect 6211 9640 6220 9680
rect 6260 9640 6268 9680
rect 6308 9640 6391 9680
rect 6595 9640 6604 9680
rect 6644 9640 6652 9680
rect 6692 9640 6775 9680
rect 6979 9640 6988 9680
rect 7028 9640 7036 9680
rect 7076 9640 7159 9680
rect 7363 9640 7372 9680
rect 7412 9640 7420 9680
rect 7460 9640 7543 9680
rect 7747 9640 7756 9680
rect 7796 9640 7804 9680
rect 7844 9640 7927 9680
rect 8131 9640 8140 9680
rect 8180 9640 8188 9680
rect 8228 9640 8311 9680
rect 8515 9640 8524 9680
rect 8564 9640 8572 9680
rect 8612 9640 8695 9680
rect 8899 9640 8908 9680
rect 8948 9640 8956 9680
rect 8996 9640 9079 9680
rect 9283 9640 9292 9680
rect 9332 9640 9340 9680
rect 9380 9640 9463 9680
rect 9667 9640 9676 9680
rect 9716 9640 9724 9680
rect 9764 9640 9847 9680
rect 10051 9640 10060 9680
rect 10100 9640 10108 9680
rect 10148 9640 10231 9680
rect 10435 9640 10444 9680
rect 10484 9640 10492 9680
rect 10532 9640 10615 9680
rect 3436 9556 7180 9596
rect 7220 9556 7229 9596
rect 3436 9512 3476 9556
rect 10732 9512 10772 10060
rect 53190 10016 53280 10036
rect 11116 9976 16012 10016
rect 16052 9976 16061 10016
rect 16291 9976 16300 10016
rect 16340 9976 19468 10016
rect 19508 9976 19517 10016
rect 28579 9976 28588 10016
rect 28628 9976 50956 10016
rect 50996 9976 51005 10016
rect 51139 9976 51148 10016
rect 51188 9976 53280 10016
rect 10819 9640 10828 9680
rect 10868 9640 10876 9680
rect 10916 9640 10999 9680
rect 11116 9596 11156 9976
rect 53190 9956 53280 9976
rect 11500 9892 13228 9932
rect 13268 9892 13277 9932
rect 13324 9892 13804 9932
rect 13844 9892 13853 9932
rect 14179 9892 14188 9932
rect 14228 9892 22828 9932
rect 22868 9892 22877 9932
rect 25507 9892 25516 9932
rect 25556 9892 44564 9932
rect 11203 9640 11212 9680
rect 11252 9640 11260 9680
rect 11300 9640 11383 9680
rect 11020 9556 11156 9596
rect 3043 9472 3052 9512
rect 3092 9472 3101 9512
rect 3427 9472 3436 9512
rect 3476 9472 3485 9512
rect 3811 9472 3820 9512
rect 3860 9472 3869 9512
rect 4073 9472 4108 9512
rect 4148 9472 4204 9512
rect 4244 9472 4253 9512
rect 4457 9472 4588 9512
rect 4628 9472 4637 9512
rect 4963 9472 4972 9512
rect 5012 9472 5021 9512
rect 5225 9472 5356 9512
rect 5396 9472 5405 9512
rect 5731 9472 5740 9512
rect 5780 9472 6068 9512
rect 6115 9472 6124 9512
rect 6164 9472 6173 9512
rect 6499 9472 6508 9512
rect 6548 9472 6557 9512
rect 6761 9472 6892 9512
rect 6932 9472 6941 9512
rect 7075 9472 7084 9512
rect 7124 9472 7276 9512
rect 7316 9472 7325 9512
rect 7651 9472 7660 9512
rect 7700 9472 7988 9512
rect 8035 9472 8044 9512
rect 8084 9472 8215 9512
rect 8419 9472 8428 9512
rect 8468 9472 8599 9512
rect 8681 9472 8812 9512
rect 8852 9472 8861 9512
rect 9065 9472 9196 9512
rect 9236 9472 9245 9512
rect 9449 9472 9580 9512
rect 9620 9472 9629 9512
rect 9833 9472 9964 9512
rect 10004 9472 10013 9512
rect 10217 9472 10348 9512
rect 10388 9472 10397 9512
rect 10723 9472 10732 9512
rect 10772 9472 10781 9512
rect 3820 9428 3860 9472
rect 4972 9428 5012 9472
rect 6028 9428 6068 9472
rect 3820 9388 4300 9428
rect 4340 9388 4349 9428
rect 4972 9388 5644 9428
rect 5684 9388 5693 9428
rect 6019 9388 6028 9428
rect 6068 9388 6077 9428
rect 0 9344 90 9364
rect 6124 9344 6164 9472
rect 6508 9428 6548 9472
rect 7948 9428 7988 9472
rect 11020 9428 11060 9556
rect 11500 9512 11540 9892
rect 13324 9848 13364 9892
rect 11884 9808 13364 9848
rect 13420 9808 18412 9848
rect 18452 9808 18461 9848
rect 18799 9808 18808 9848
rect 18848 9808 18890 9848
rect 18930 9808 18972 9848
rect 19012 9808 19054 9848
rect 19094 9808 19136 9848
rect 19176 9808 19185 9848
rect 19459 9808 19468 9848
rect 19508 9808 22444 9848
rect 22484 9808 22493 9848
rect 22540 9808 31180 9848
rect 31220 9808 31229 9848
rect 33919 9808 33928 9848
rect 33968 9808 34010 9848
rect 34050 9808 34092 9848
rect 34132 9808 34174 9848
rect 34214 9808 34256 9848
rect 34296 9808 34305 9848
rect 11587 9640 11596 9680
rect 11636 9640 11644 9680
rect 11684 9640 11767 9680
rect 11884 9512 11924 9808
rect 11971 9640 11980 9680
rect 12020 9640 12028 9680
rect 12068 9640 12151 9680
rect 12355 9640 12364 9680
rect 12404 9640 12412 9680
rect 12452 9640 12535 9680
rect 12739 9640 12748 9680
rect 12788 9640 12796 9680
rect 12836 9640 12919 9680
rect 13123 9640 13132 9680
rect 13172 9640 13180 9680
rect 13220 9640 13303 9680
rect 12268 9556 13324 9596
rect 13364 9556 13373 9596
rect 12268 9512 12308 9556
rect 13420 9512 13460 9808
rect 22540 9764 22580 9808
rect 13804 9724 18316 9764
rect 18356 9724 18365 9764
rect 19084 9724 20140 9764
rect 20180 9724 20189 9764
rect 20323 9724 20332 9764
rect 20372 9724 22580 9764
rect 23020 9724 34636 9764
rect 34676 9724 34685 9764
rect 13507 9640 13516 9680
rect 13556 9640 13564 9680
rect 13604 9640 13687 9680
rect 13804 9512 13844 9724
rect 13891 9640 13900 9680
rect 13940 9640 13948 9680
rect 13988 9640 14071 9680
rect 14275 9640 14284 9680
rect 14324 9640 14332 9680
rect 14372 9640 14455 9680
rect 14659 9640 14668 9680
rect 14708 9640 14716 9680
rect 14756 9640 14839 9680
rect 15043 9640 15052 9680
rect 15092 9640 15100 9680
rect 15140 9640 15223 9680
rect 15427 9640 15436 9680
rect 15476 9640 15484 9680
rect 15524 9640 15607 9680
rect 15811 9640 15820 9680
rect 15860 9640 15868 9680
rect 15908 9640 15991 9680
rect 16195 9640 16204 9680
rect 16244 9640 16252 9680
rect 16292 9640 16375 9680
rect 16579 9640 16588 9680
rect 16628 9640 16636 9680
rect 16676 9640 16759 9680
rect 16963 9640 16972 9680
rect 17012 9640 17020 9680
rect 17060 9640 17143 9680
rect 17347 9640 17356 9680
rect 17396 9640 17404 9680
rect 17444 9640 17527 9680
rect 17731 9640 17740 9680
rect 17780 9640 17788 9680
rect 17828 9640 17911 9680
rect 18115 9640 18124 9680
rect 18164 9640 18172 9680
rect 18212 9640 18295 9680
rect 18499 9640 18508 9680
rect 18548 9640 18556 9680
rect 18596 9640 18679 9680
rect 16108 9556 17932 9596
rect 17972 9556 17981 9596
rect 18691 9556 18700 9596
rect 18740 9556 18940 9596
rect 18980 9556 18989 9596
rect 16108 9512 16148 9556
rect 19084 9512 19124 9724
rect 23020 9680 23060 9724
rect 19267 9640 19276 9680
rect 19316 9640 19324 9680
rect 19364 9640 19447 9680
rect 19651 9640 19660 9680
rect 19700 9640 19708 9680
rect 19748 9640 19831 9680
rect 20035 9640 20044 9680
rect 20084 9640 20092 9680
rect 20132 9640 20215 9680
rect 20419 9640 20428 9680
rect 20468 9640 20476 9680
rect 20516 9640 20599 9680
rect 20803 9640 20812 9680
rect 20852 9640 20860 9680
rect 20900 9640 20983 9680
rect 21187 9640 21196 9680
rect 21236 9640 21244 9680
rect 21284 9640 21367 9680
rect 21571 9640 21580 9680
rect 21620 9640 21628 9680
rect 21668 9640 21751 9680
rect 21955 9640 21964 9680
rect 22004 9640 22012 9680
rect 22052 9640 22135 9680
rect 22339 9640 22348 9680
rect 22388 9640 22396 9680
rect 22436 9640 22519 9680
rect 22627 9640 22636 9680
rect 22676 9640 23060 9680
rect 23875 9640 23884 9680
rect 23924 9640 36172 9680
rect 36212 9640 36221 9680
rect 42691 9640 42700 9680
rect 42740 9640 42748 9680
rect 42788 9640 42871 9680
rect 43001 9640 43084 9680
rect 43124 9640 43132 9680
rect 43172 9640 43181 9680
rect 43459 9640 43468 9680
rect 43508 9640 43516 9680
rect 43556 9640 43639 9680
rect 43843 9640 43852 9680
rect 43892 9640 43900 9680
rect 43940 9640 44023 9680
rect 44227 9640 44236 9680
rect 44276 9640 44284 9680
rect 44324 9640 44407 9680
rect 19564 9556 20620 9596
rect 20660 9556 20669 9596
rect 20716 9556 21772 9596
rect 21812 9556 21821 9596
rect 21868 9556 28780 9596
rect 28820 9556 28829 9596
rect 19564 9512 19604 9556
rect 20716 9512 20756 9556
rect 21868 9512 21908 9556
rect 44524 9512 44564 9892
rect 49039 9808 49048 9848
rect 49088 9808 49130 9848
rect 49170 9808 49212 9848
rect 49252 9808 49294 9848
rect 49334 9808 49376 9848
rect 49416 9808 49425 9848
rect 47107 9724 47116 9764
rect 47156 9724 51860 9764
rect 44611 9640 44620 9680
rect 44660 9640 44668 9680
rect 44708 9640 44791 9680
rect 44995 9640 45004 9680
rect 45044 9640 45052 9680
rect 45092 9640 45175 9680
rect 45379 9640 45388 9680
rect 45428 9640 45436 9680
rect 45476 9640 45559 9680
rect 45763 9640 45772 9680
rect 45812 9640 45820 9680
rect 45860 9640 45943 9680
rect 46147 9640 46156 9680
rect 46196 9640 46204 9680
rect 46244 9640 46327 9680
rect 46531 9640 46540 9680
rect 46580 9640 46588 9680
rect 46628 9640 46711 9680
rect 46915 9640 46924 9680
rect 46964 9640 46972 9680
rect 47012 9640 47095 9680
rect 47299 9640 47308 9680
rect 47348 9640 47356 9680
rect 47396 9640 47479 9680
rect 47683 9640 47692 9680
rect 47732 9640 47740 9680
rect 47780 9640 47863 9680
rect 48067 9640 48076 9680
rect 48116 9640 48124 9680
rect 48164 9640 48247 9680
rect 48451 9640 48460 9680
rect 48500 9640 48508 9680
rect 48548 9640 48631 9680
rect 48835 9640 48844 9680
rect 48884 9640 48892 9680
rect 48932 9640 49015 9680
rect 49267 9640 49276 9680
rect 49316 9640 49516 9680
rect 49556 9640 49565 9680
rect 49987 9640 49996 9680
rect 50036 9640 50044 9680
rect 50084 9640 50167 9680
rect 50371 9640 50380 9680
rect 50420 9640 50428 9680
rect 50468 9640 50551 9680
rect 49603 9556 49612 9596
rect 49652 9556 49660 9596
rect 49700 9556 49783 9596
rect 50764 9556 51476 9596
rect 11107 9472 11116 9512
rect 11156 9472 11287 9512
rect 11491 9472 11500 9512
rect 11540 9472 11549 9512
rect 11875 9472 11884 9512
rect 11924 9472 11933 9512
rect 12259 9472 12268 9512
rect 12308 9472 12317 9512
rect 12521 9472 12652 9512
rect 12692 9472 12701 9512
rect 13027 9472 13036 9512
rect 13076 9472 13228 9512
rect 13268 9472 13277 9512
rect 13411 9472 13420 9512
rect 13460 9472 13469 9512
rect 13795 9472 13804 9512
rect 13844 9472 13853 9512
rect 14179 9472 14188 9512
rect 14228 9472 14237 9512
rect 14563 9472 14572 9512
rect 14612 9472 14621 9512
rect 14947 9472 14956 9512
rect 14996 9472 15148 9512
rect 15188 9472 15197 9512
rect 15331 9472 15340 9512
rect 15380 9472 15389 9512
rect 15715 9472 15724 9512
rect 15764 9472 15916 9512
rect 15956 9472 15965 9512
rect 16099 9472 16108 9512
rect 16148 9472 16157 9512
rect 16483 9472 16492 9512
rect 16532 9472 16541 9512
rect 16867 9472 16876 9512
rect 16916 9472 16925 9512
rect 17251 9472 17260 9512
rect 17300 9472 17309 9512
rect 17635 9472 17644 9512
rect 17684 9472 17972 9512
rect 18019 9472 18028 9512
rect 18068 9472 18356 9512
rect 18403 9472 18412 9512
rect 18452 9472 18604 9512
rect 18644 9472 18653 9512
rect 18787 9472 18796 9512
rect 18836 9472 19124 9512
rect 19171 9472 19180 9512
rect 19220 9472 19229 9512
rect 19555 9472 19564 9512
rect 19604 9472 19613 9512
rect 19817 9472 19948 9512
rect 19988 9472 19997 9512
rect 20323 9472 20332 9512
rect 20372 9472 20524 9512
rect 20564 9472 20573 9512
rect 20707 9472 20716 9512
rect 20756 9472 20765 9512
rect 21091 9472 21100 9512
rect 21140 9472 21292 9512
rect 21332 9472 21341 9512
rect 21475 9472 21484 9512
rect 21524 9472 21676 9512
rect 21716 9472 21725 9512
rect 21859 9472 21868 9512
rect 21908 9472 21917 9512
rect 22243 9472 22252 9512
rect 22292 9472 22348 9512
rect 22388 9472 22423 9512
rect 22627 9472 22636 9512
rect 22676 9472 23020 9512
rect 23060 9472 23069 9512
rect 24748 9472 36940 9512
rect 36980 9472 36989 9512
rect 40291 9472 40300 9512
rect 40340 9472 42988 9512
rect 43028 9472 43037 9512
rect 43084 9472 43372 9512
rect 43412 9472 43421 9512
rect 43747 9472 43756 9512
rect 43796 9472 43805 9512
rect 44131 9472 44140 9512
rect 44180 9472 44189 9512
rect 44515 9472 44524 9512
rect 44564 9472 44573 9512
rect 44899 9472 44908 9512
rect 44948 9472 44957 9512
rect 45283 9472 45292 9512
rect 45332 9472 45341 9512
rect 45667 9472 45676 9512
rect 45716 9472 45725 9512
rect 45929 9472 46060 9512
rect 46100 9472 46109 9512
rect 46313 9472 46444 9512
rect 46484 9472 46493 9512
rect 46697 9472 46828 9512
rect 46868 9472 46877 9512
rect 47081 9472 47212 9512
rect 47252 9472 47261 9512
rect 47395 9472 47404 9512
rect 47444 9472 47596 9512
rect 47636 9472 47645 9512
rect 47849 9472 47980 9512
rect 48020 9472 48029 9512
rect 48233 9472 48364 9512
rect 48404 9472 48413 9512
rect 48617 9472 48748 9512
rect 48788 9472 48797 9512
rect 49001 9472 49036 9512
rect 49076 9472 49132 9512
rect 49172 9472 49181 9512
rect 49228 9472 49516 9512
rect 49556 9472 49565 9512
rect 49891 9472 49900 9512
rect 49940 9472 49949 9512
rect 50083 9472 50092 9512
rect 50132 9472 50284 9512
rect 50324 9472 50333 9512
rect 50659 9472 50668 9512
rect 50708 9472 50717 9512
rect 6508 9388 7756 9428
rect 7796 9388 7805 9428
rect 7948 9388 11060 9428
rect 0 9304 268 9344
rect 308 9304 317 9344
rect 6124 9304 10156 9344
rect 10196 9304 10205 9344
rect 0 9284 90 9304
rect 14188 9176 14228 9472
rect 14572 9344 14612 9472
rect 15340 9428 15380 9472
rect 15340 9388 16396 9428
rect 16436 9388 16445 9428
rect 14572 9304 16300 9344
rect 16340 9304 16349 9344
rect 16492 9176 16532 9472
rect 16876 9260 16916 9472
rect 17260 9428 17300 9472
rect 17260 9388 17836 9428
rect 17876 9388 17885 9428
rect 17932 9344 17972 9472
rect 18316 9428 18356 9472
rect 18316 9388 19084 9428
rect 19124 9388 19133 9428
rect 19180 9344 19220 9472
rect 19267 9388 19276 9428
rect 19316 9388 22252 9428
rect 22292 9388 22301 9428
rect 24748 9344 24788 9472
rect 43084 9428 43124 9472
rect 43756 9428 43796 9472
rect 24931 9388 24940 9428
rect 24980 9388 32716 9428
rect 32756 9388 32765 9428
rect 40579 9388 40588 9428
rect 40628 9388 43124 9428
rect 43171 9388 43180 9428
rect 43220 9388 43796 9428
rect 44140 9344 44180 9472
rect 44908 9428 44948 9472
rect 44227 9388 44236 9428
rect 44276 9388 44948 9428
rect 17932 9304 18988 9344
rect 19028 9304 19037 9344
rect 19180 9304 22156 9344
rect 22196 9304 22205 9344
rect 22339 9304 22348 9344
rect 22388 9304 24788 9344
rect 24835 9304 24844 9344
rect 24884 9304 35020 9344
rect 35060 9304 35069 9344
rect 40483 9304 40492 9344
rect 40532 9304 44180 9344
rect 45292 9260 45332 9472
rect 16876 9220 20140 9260
rect 20180 9220 20189 9260
rect 20284 9220 22924 9260
rect 22964 9220 22973 9260
rect 23020 9220 35404 9260
rect 35444 9220 35453 9260
rect 41731 9220 41740 9260
rect 41780 9220 45332 9260
rect 20284 9176 20324 9220
rect 23020 9176 23060 9220
rect 45676 9176 45716 9472
rect 49228 9428 49268 9472
rect 8035 9136 8044 9176
rect 8084 9136 12940 9176
rect 12980 9136 12989 9176
rect 14188 9136 16436 9176
rect 16492 9136 18700 9176
rect 18740 9136 18749 9176
rect 19075 9136 19084 9176
rect 19124 9136 19660 9176
rect 19700 9136 19709 9176
rect 19939 9136 19948 9176
rect 19988 9136 20324 9176
rect 22723 9136 22732 9176
rect 22772 9136 23060 9176
rect 27715 9136 27724 9176
rect 27764 9136 31468 9176
rect 31508 9136 31517 9176
rect 41827 9136 41836 9176
rect 41876 9136 45716 9176
rect 46348 9388 49268 9428
rect 16396 9092 16436 9136
rect 46348 9092 46388 9388
rect 49900 9344 49940 9472
rect 50668 9428 50708 9472
rect 49987 9388 49996 9428
rect 50036 9388 50708 9428
rect 46723 9304 46732 9344
rect 46772 9304 49940 9344
rect 50764 9176 50804 9556
rect 51436 9512 51476 9556
rect 51820 9512 51860 9724
rect 53190 9680 53280 9700
rect 51916 9640 53280 9680
rect 51043 9472 51052 9512
rect 51092 9472 51223 9512
rect 51427 9472 51436 9512
rect 51476 9472 51485 9512
rect 51811 9472 51820 9512
rect 51860 9472 51869 9512
rect 51916 9428 51956 9640
rect 53190 9620 53280 9640
rect 4919 9052 4928 9092
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 5296 9052 5305 9092
rect 6019 9052 6028 9092
rect 6068 9052 11500 9092
rect 11540 9052 11549 9092
rect 11692 9052 15052 9092
rect 15092 9052 15101 9092
rect 16396 9052 17548 9092
rect 17588 9052 17597 9092
rect 17644 9052 19988 9092
rect 20039 9052 20048 9092
rect 20088 9052 20130 9092
rect 20170 9052 20212 9092
rect 20252 9052 20294 9092
rect 20334 9052 20376 9092
rect 20416 9052 20425 9092
rect 20611 9052 20620 9092
rect 20660 9052 24172 9092
rect 24212 9052 24221 9092
rect 30211 9052 30220 9092
rect 30260 9052 31084 9092
rect 31124 9052 31133 9092
rect 35159 9052 35168 9092
rect 35208 9052 35250 9092
rect 35290 9052 35332 9092
rect 35372 9052 35414 9092
rect 35454 9052 35496 9092
rect 35536 9052 35545 9092
rect 37987 9052 37996 9092
rect 38036 9052 42316 9092
rect 42356 9052 42365 9092
rect 42595 9052 42604 9092
rect 42644 9052 46388 9092
rect 47308 9136 50804 9176
rect 51148 9388 51956 9428
rect 0 9008 90 9028
rect 0 8968 11596 9008
rect 11636 8968 11645 9008
rect 0 8948 90 8968
rect 11692 8924 11732 9052
rect 11779 8968 11788 9008
rect 11828 8968 17452 9008
rect 17492 8968 17501 9008
rect 17644 8924 17684 9052
rect 19948 9008 19988 9052
rect 47308 9008 47348 9136
rect 18595 8968 18604 9008
rect 18644 8968 19756 9008
rect 19796 8968 19805 9008
rect 19948 8968 21484 9008
rect 21524 8968 21533 9008
rect 23107 8968 23116 9008
rect 23156 8968 23348 9008
rect 23308 8924 23348 8968
rect 28012 8968 29356 9008
rect 29396 8968 29405 9008
rect 29548 8968 30988 9008
rect 31028 8968 31037 9008
rect 31363 8968 31372 9008
rect 31412 8968 47348 9008
rect 47404 9052 50188 9092
rect 50228 9052 50237 9092
rect 50279 9052 50288 9092
rect 50328 9052 50370 9092
rect 50410 9052 50452 9092
rect 50492 9052 50534 9092
rect 50574 9052 50616 9092
rect 50656 9052 50665 9092
rect 28012 8924 28052 8968
rect 29548 8924 29588 8968
rect 47404 8924 47444 9052
rect 5635 8884 5644 8924
rect 5684 8884 11732 8924
rect 12940 8884 13708 8924
rect 13748 8884 13757 8924
rect 13891 8884 13900 8924
rect 13940 8884 17684 8924
rect 17740 8884 20236 8924
rect 20276 8884 20285 8924
rect 20707 8884 20716 8924
rect 20756 8884 21628 8924
rect 21668 8884 21677 8924
rect 22147 8884 22156 8924
rect 22196 8884 22636 8924
rect 22676 8884 22685 8924
rect 22819 8884 22828 8924
rect 22868 8884 23068 8924
rect 23108 8884 23117 8924
rect 23308 8884 23644 8924
rect 23684 8884 23693 8924
rect 26995 8884 27004 8924
rect 27044 8884 28052 8924
rect 28147 8884 28156 8924
rect 28196 8884 28820 8924
rect 28915 8884 28924 8924
rect 28964 8884 29588 8924
rect 29683 8884 29692 8924
rect 29732 8884 31276 8924
rect 31316 8884 31325 8924
rect 31459 8884 31468 8924
rect 31508 8884 47444 8924
rect 50092 8968 50860 9008
rect 50900 8968 50909 9008
rect 50092 8924 50132 8968
rect 51148 8924 51188 9388
rect 53190 9344 53280 9364
rect 51283 9304 51292 9344
rect 51332 9304 53280 9344
rect 53190 9284 53280 9304
rect 51667 9220 51676 9260
rect 51716 9220 51725 9260
rect 52051 9220 52060 9260
rect 52100 9220 52684 9260
rect 52724 9220 52733 9260
rect 51676 8924 51716 9220
rect 53190 9008 53280 9028
rect 53164 8948 53280 9008
rect 53164 8924 53204 8948
rect 50092 8884 50140 8924
rect 50180 8884 50189 8924
rect 50515 8884 50524 8924
rect 50564 8884 50764 8924
rect 50804 8884 50813 8924
rect 50899 8884 50908 8924
rect 50948 8884 51052 8924
rect 51092 8884 51101 8924
rect 51148 8884 51292 8924
rect 51332 8884 51341 8924
rect 51676 8884 53204 8924
rect 12940 8840 12980 8884
rect 17740 8840 17780 8884
rect 5347 8800 5356 8840
rect 5396 8800 12980 8840
rect 13315 8800 13324 8840
rect 13364 8800 17780 8840
rect 17827 8800 17836 8840
rect 17876 8800 20276 8840
rect 20236 8756 20276 8800
rect 20476 8800 28724 8840
rect 20476 8756 20516 8800
rect 13219 8716 13228 8756
rect 13268 8716 20140 8756
rect 20180 8716 20189 8756
rect 20236 8716 20516 8756
rect 22348 8716 24844 8756
rect 24884 8716 24893 8756
rect 25027 8716 25036 8756
rect 25076 8716 28340 8756
rect 28579 8716 28588 8756
rect 28628 8716 28637 8756
rect 0 8672 90 8692
rect 22348 8672 22388 8716
rect 28300 8672 28340 8716
rect 28588 8672 28628 8716
rect 28684 8672 28724 8800
rect 28780 8756 28820 8884
rect 29299 8800 29308 8840
rect 29348 8800 47116 8840
rect 47156 8800 47165 8840
rect 47395 8800 47404 8840
rect 47444 8800 51860 8840
rect 28780 8716 50036 8756
rect 0 8632 1420 8672
rect 1460 8632 1469 8672
rect 12643 8632 12652 8672
rect 12692 8632 20716 8672
rect 20756 8632 20765 8672
rect 21737 8632 21868 8672
rect 21908 8632 21917 8672
rect 22339 8632 22348 8672
rect 22388 8632 22397 8672
rect 22601 8632 22732 8672
rect 22772 8632 22781 8672
rect 23177 8632 23308 8672
rect 23348 8632 23357 8672
rect 23753 8632 23884 8672
rect 23924 8632 23933 8672
rect 26633 8632 26764 8672
rect 26804 8632 26813 8672
rect 27017 8632 27148 8672
rect 27188 8632 27197 8672
rect 27401 8632 27532 8672
rect 27572 8632 27581 8672
rect 27715 8632 27724 8672
rect 27764 8632 27772 8672
rect 27812 8632 27895 8672
rect 27946 8632 27955 8672
rect 27995 8632 28012 8672
rect 28052 8632 28135 8672
rect 28291 8632 28300 8672
rect 28340 8632 28349 8672
rect 28531 8632 28540 8672
rect 28580 8632 28628 8672
rect 28675 8632 28684 8672
rect 28724 8632 28733 8672
rect 28937 8632 29068 8672
rect 29108 8632 29117 8672
rect 29321 8632 29452 8672
rect 29492 8632 29501 8672
rect 31171 8632 31180 8672
rect 31220 8632 31228 8672
rect 31268 8632 31351 8672
rect 31459 8632 31468 8672
rect 31508 8632 37996 8672
rect 38036 8632 38045 8672
rect 38179 8632 38188 8672
rect 38228 8632 49900 8672
rect 49940 8632 49949 8672
rect 0 8612 90 8632
rect 49996 8588 50036 8716
rect 51820 8672 51860 8800
rect 53190 8672 53280 8692
rect 50153 8632 50284 8672
rect 50324 8632 50333 8672
rect 50380 8632 50668 8672
rect 50708 8632 50717 8672
rect 50921 8632 50956 8672
rect 50996 8632 51052 8672
rect 51092 8632 51101 8672
rect 51305 8632 51436 8672
rect 51476 8632 51485 8672
rect 51811 8632 51820 8672
rect 51860 8632 51869 8672
rect 52675 8632 52684 8672
rect 52724 8632 53280 8672
rect 50380 8588 50420 8632
rect 53190 8612 53280 8632
rect 6115 8548 6124 8588
rect 6164 8548 18028 8588
rect 18068 8548 18077 8588
rect 18595 8548 18604 8588
rect 18644 8548 25228 8588
rect 25268 8548 25277 8588
rect 27379 8548 27388 8588
rect 27428 8548 30220 8588
rect 30260 8548 30269 8588
rect 30316 8548 35252 8588
rect 35299 8548 35308 8588
rect 35348 8548 40396 8588
rect 40436 8548 40445 8588
rect 49996 8548 50420 8588
rect 30316 8504 30356 8548
rect 35212 8504 35252 8548
rect 172 8464 15820 8504
rect 15860 8464 15869 8504
rect 15916 8464 17068 8504
rect 17108 8464 17117 8504
rect 18211 8464 18220 8504
rect 18260 8464 19852 8504
rect 19892 8464 19901 8504
rect 20035 8464 20044 8504
rect 20084 8464 20332 8504
rect 20372 8464 20381 8504
rect 21475 8464 21484 8504
rect 21524 8464 22108 8504
rect 22148 8464 22157 8504
rect 22435 8464 22444 8504
rect 22484 8464 22492 8504
rect 22532 8464 22615 8504
rect 22915 8464 22924 8504
rect 22964 8464 30356 8504
rect 31075 8464 31084 8504
rect 31124 8464 32908 8504
rect 32948 8464 32957 8504
rect 35212 8464 37132 8504
rect 37172 8464 37181 8504
rect 37603 8464 37612 8504
rect 37652 8464 40012 8504
rect 40052 8464 40061 8504
rect 51667 8464 51676 8504
rect 51716 8464 51956 8504
rect 52051 8464 52060 8504
rect 52100 8464 52684 8504
rect 52724 8464 52733 8504
rect 0 8336 90 8356
rect 172 8336 212 8464
rect 15916 8420 15956 8464
rect 4588 8380 10060 8420
rect 10100 8380 10109 8420
rect 15907 8380 15916 8420
rect 15956 8380 15965 8420
rect 16291 8380 16300 8420
rect 16340 8380 16780 8420
rect 16820 8380 16829 8420
rect 16876 8380 23500 8420
rect 23540 8380 23549 8420
rect 24163 8380 24172 8420
rect 24212 8380 32812 8420
rect 32852 8380 32861 8420
rect 37795 8380 37804 8420
rect 37844 8380 39628 8420
rect 39668 8380 39677 8420
rect 0 8296 212 8336
rect 3679 8296 3688 8336
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 4056 8296 4065 8336
rect 0 8276 90 8296
rect 3475 8128 3484 8168
rect 3524 8128 4108 8168
rect 4148 8128 4157 8168
rect 4291 8128 4300 8168
rect 4340 8128 4348 8168
rect 4388 8128 4471 8168
rect 0 8000 90 8020
rect 4588 8000 4628 8380
rect 16876 8336 16916 8380
rect 51916 8336 51956 8464
rect 53190 8336 53280 8356
rect 9964 8296 10100 8336
rect 10243 8296 10252 8336
rect 10292 8296 16916 8336
rect 18799 8296 18808 8336
rect 18848 8296 18890 8336
rect 18930 8296 18972 8336
rect 19012 8296 19054 8336
rect 19094 8296 19136 8336
rect 19176 8296 19185 8336
rect 19660 8296 20140 8336
rect 20180 8296 20189 8336
rect 20323 8296 20332 8336
rect 20372 8296 31852 8336
rect 31892 8296 31901 8336
rect 33919 8296 33928 8336
rect 33968 8296 34010 8336
rect 34050 8296 34092 8336
rect 34132 8296 34174 8336
rect 34214 8296 34256 8336
rect 34296 8296 34305 8336
rect 37699 8296 37708 8336
rect 37748 8296 39052 8336
rect 39092 8296 39101 8336
rect 39331 8296 39340 8336
rect 39380 8296 41548 8336
rect 41588 8296 41597 8336
rect 49039 8296 49048 8336
rect 49088 8296 49130 8336
rect 49170 8296 49212 8336
rect 49252 8296 49294 8336
rect 49334 8296 49376 8336
rect 49416 8296 49425 8336
rect 51916 8296 53280 8336
rect 6355 8128 6364 8168
rect 6404 8128 6892 8168
rect 6932 8128 6941 8168
rect 7747 8128 7756 8168
rect 7796 8128 7804 8168
rect 7844 8128 7927 8168
rect 9964 8084 10004 8296
rect 5491 8044 5500 8084
rect 5540 8044 7084 8084
rect 7124 8044 7133 8084
rect 8428 8044 10004 8084
rect 10060 8084 10100 8296
rect 10147 8128 10156 8168
rect 10196 8128 10204 8168
rect 10244 8128 10327 8168
rect 10444 8128 12844 8168
rect 12884 8128 12893 8168
rect 13027 8128 13036 8168
rect 13076 8128 15292 8168
rect 15332 8128 15341 8168
rect 15619 8128 15628 8168
rect 15668 8128 15676 8168
rect 15716 8128 15799 8168
rect 16003 8128 16012 8168
rect 16052 8128 16060 8168
rect 16100 8128 16183 8168
rect 16387 8128 16396 8168
rect 16436 8128 16444 8168
rect 16484 8128 16567 8168
rect 16697 8128 16780 8168
rect 16820 8128 16828 8168
rect 16868 8128 16877 8168
rect 16972 8128 17260 8168
rect 17300 8128 17309 8168
rect 17539 8128 17548 8168
rect 17588 8128 17596 8168
rect 17636 8128 17719 8168
rect 17923 8128 17932 8168
rect 17972 8128 17980 8168
rect 18020 8128 18103 8168
rect 18307 8128 18316 8168
rect 18356 8128 18364 8168
rect 18404 8128 18487 8168
rect 18691 8128 18700 8168
rect 18740 8128 19036 8168
rect 19076 8128 19085 8168
rect 10060 8044 10252 8084
rect 10292 8044 10301 8084
rect 8428 8000 8468 8044
rect 10444 8000 10484 8128
rect 11491 8044 11500 8084
rect 11540 8044 11932 8084
rect 11972 8044 11981 8084
rect 12163 8044 12172 8084
rect 12212 8044 15860 8084
rect 0 7960 1228 8000
rect 1268 7960 1277 8000
rect 3235 7960 3244 8000
rect 3284 7960 3293 8000
rect 4579 7960 4588 8000
rect 4628 7960 4637 8000
rect 5251 7960 5260 8000
rect 5300 7960 5836 8000
rect 5876 7960 5885 8000
rect 5993 7960 6124 8000
rect 6164 7960 6173 8000
rect 8035 7960 8044 8000
rect 8084 7960 8093 8000
rect 8419 7960 8428 8000
rect 8468 7960 8477 8000
rect 10435 7960 10444 8000
rect 10484 7960 10493 8000
rect 10579 7960 10588 8000
rect 10628 7960 10636 8000
rect 10676 7960 10759 8000
rect 10819 7960 10828 8000
rect 10868 7960 12116 8000
rect 12163 7960 12172 8000
rect 12212 7960 15340 8000
rect 15380 7960 15389 8000
rect 15523 7960 15532 8000
rect 15572 7960 15581 8000
rect 0 7940 90 7960
rect 0 7664 90 7684
rect 3244 7664 3284 7960
rect 8044 7916 8084 7960
rect 12076 7916 12116 7960
rect 8044 7876 10060 7916
rect 10100 7876 10109 7916
rect 12076 7876 15436 7916
rect 15476 7876 15485 7916
rect 7171 7792 7180 7832
rect 7220 7792 8188 7832
rect 8228 7792 8237 7832
rect 15532 7664 15572 7960
rect 15820 7748 15860 8044
rect 16972 8000 17012 8128
rect 17059 8044 17068 8084
rect 17108 8044 17212 8084
rect 17252 8044 17261 8084
rect 18403 8044 18412 8084
rect 18452 8044 19420 8084
rect 19460 8044 19469 8084
rect 19660 8000 19700 8296
rect 53190 8276 53280 8296
rect 20044 8212 25132 8252
rect 25172 8212 25181 8252
rect 25315 8212 25324 8252
rect 25364 8212 35404 8252
rect 35444 8212 35453 8252
rect 38764 8212 47980 8252
rect 48020 8212 48029 8252
rect 15907 7960 15916 8000
rect 15956 7960 16108 8000
rect 16148 7960 16157 8000
rect 16291 7960 16300 8000
rect 16340 7960 16349 8000
rect 16675 7960 16684 8000
rect 16724 7960 17012 8000
rect 17059 7960 17068 8000
rect 17108 7960 17117 8000
rect 17321 7960 17452 8000
rect 17492 7960 17501 8000
rect 17705 7960 17836 8000
rect 17876 7960 17885 8000
rect 18089 7960 18220 8000
rect 18260 7960 18269 8000
rect 18473 7960 18604 8000
rect 18644 7960 18653 8000
rect 19145 7960 19276 8000
rect 19316 7960 19325 8000
rect 19651 7960 19660 8000
rect 19700 7960 19709 8000
rect 16300 7832 16340 7960
rect 17068 7916 17108 7960
rect 20044 7916 20084 8212
rect 38764 8168 38804 8212
rect 20707 8128 20716 8168
rect 20756 8128 20764 8168
rect 20804 8128 20887 8168
rect 25027 8128 25036 8168
rect 25076 8128 30028 8168
rect 30068 8128 30077 8168
rect 32707 8128 32716 8168
rect 32756 8128 32764 8168
rect 32804 8128 32887 8168
rect 35692 8128 36556 8168
rect 36596 8128 36605 8168
rect 36931 8128 36940 8168
rect 36980 8128 37084 8168
rect 37124 8128 37133 8168
rect 37411 8128 37420 8168
rect 37460 8128 37468 8168
rect 37508 8128 37591 8168
rect 37891 8128 37900 8168
rect 37940 8128 37949 8168
rect 38131 8128 38140 8168
rect 38180 8128 38804 8168
rect 38851 8128 38860 8168
rect 38900 8128 39668 8168
rect 51283 8128 51292 8168
rect 51332 8128 52300 8168
rect 52340 8128 52349 8168
rect 20227 8044 20236 8084
rect 20276 8044 20284 8084
rect 20324 8044 20407 8084
rect 20524 8044 28492 8084
rect 28532 8044 28541 8084
rect 28588 8044 28636 8084
rect 28676 8044 28685 8084
rect 30220 8044 33292 8084
rect 33332 8044 33341 8084
rect 33475 8044 33484 8084
rect 33524 8044 35068 8084
rect 35108 8044 35117 8084
rect 20524 8000 20564 8044
rect 28588 8000 28628 8044
rect 30220 8000 30260 8044
rect 35692 8000 35732 8128
rect 36076 8044 37612 8084
rect 37652 8044 37661 8084
rect 37795 8044 37804 8084
rect 37844 8044 37853 8084
rect 36076 8000 36116 8044
rect 37804 8000 37844 8044
rect 37900 8000 37940 8128
rect 38860 8044 39244 8084
rect 39284 8044 39293 8084
rect 39379 8044 39388 8084
rect 39428 8044 39436 8084
rect 39476 8044 39559 8084
rect 38860 8000 38900 8044
rect 39628 8000 39668 8128
rect 39715 8044 39724 8084
rect 39764 8044 41932 8084
rect 41972 8044 41981 8084
rect 47491 8044 47500 8084
rect 47540 8044 51476 8084
rect 51436 8000 51476 8044
rect 53190 8000 53280 8020
rect 20515 7960 20524 8000
rect 20564 7960 20573 8000
rect 20873 7960 21004 8000
rect 21044 7960 21053 8000
rect 21187 7960 21196 8000
rect 21236 7960 22540 8000
rect 22580 7960 22589 8000
rect 22723 7960 22732 8000
rect 22772 7960 25268 8000
rect 28265 7960 28396 8000
rect 28436 7960 28445 8000
rect 28579 7960 28588 8000
rect 28628 7960 28637 8000
rect 28963 7960 28972 8000
rect 29012 7960 30260 8000
rect 32995 7960 33004 8000
rect 33044 7960 33196 8000
rect 33236 7960 33245 8000
rect 33379 7960 33388 8000
rect 33428 7960 33580 8000
rect 33620 7960 33629 8000
rect 33763 7960 33772 8000
rect 33812 7960 34636 8000
rect 34676 7960 34685 8000
rect 34793 7960 34924 8000
rect 34964 7960 34973 8000
rect 35177 7960 35308 8000
rect 35348 7960 35357 8000
rect 35683 7960 35692 8000
rect 35732 7960 35741 8000
rect 36067 7960 36076 8000
rect 36116 7960 36125 8000
rect 36355 7960 36364 8000
rect 36404 7960 36556 8000
rect 36596 7960 36605 8000
rect 36739 7960 36748 8000
rect 36788 7960 36919 8000
rect 37193 7960 37228 8000
rect 37268 7960 37324 8000
rect 37364 7960 37373 8000
rect 37699 7960 37708 8000
rect 37748 7960 37844 8000
rect 37891 7960 37900 8000
rect 37940 7960 37949 8000
rect 37996 7960 38236 8000
rect 38276 7960 38285 8000
rect 38371 7960 38380 8000
rect 38420 7960 38476 8000
rect 38516 7960 38551 8000
rect 38851 7960 38860 8000
rect 38900 7960 38909 8000
rect 39043 7960 39052 8000
rect 39092 7960 39244 8000
rect 39284 7960 39293 8000
rect 39619 7960 39628 8000
rect 39668 7960 39677 8000
rect 40003 7960 40012 8000
rect 40052 7960 40061 8000
rect 51043 7960 51052 8000
rect 51092 7960 51101 8000
rect 51427 7960 51436 8000
rect 51476 7960 51485 8000
rect 51811 7960 51820 8000
rect 51860 7960 51916 8000
rect 51956 7960 51991 8000
rect 52675 7960 52684 8000
rect 52724 7960 53280 8000
rect 17068 7876 20084 7916
rect 20140 7876 25036 7916
rect 25076 7876 25085 7916
rect 20140 7832 20180 7876
rect 25228 7832 25268 7960
rect 37996 7916 38036 7960
rect 40012 7916 40052 7960
rect 28771 7876 28780 7916
rect 28820 7876 38036 7916
rect 38380 7876 39628 7916
rect 39668 7876 39677 7916
rect 39724 7876 40052 7916
rect 38380 7832 38420 7876
rect 39724 7832 39764 7876
rect 16300 7792 20180 7832
rect 20236 7792 23212 7832
rect 23252 7792 23261 7832
rect 25228 7792 28052 7832
rect 28099 7792 28108 7832
rect 28148 7792 33148 7832
rect 33188 7792 33197 7832
rect 33283 7792 33292 7832
rect 33332 7792 35452 7832
rect 35492 7792 35501 7832
rect 36979 7792 36988 7832
rect 37028 7792 38420 7832
rect 38467 7792 38476 7832
rect 38516 7792 39764 7832
rect 39811 7792 39820 7832
rect 39860 7792 48748 7832
rect 48788 7792 48797 7832
rect 20236 7748 20276 7792
rect 28012 7748 28052 7792
rect 15820 7708 17644 7748
rect 17684 7708 17693 7748
rect 17827 7708 17836 7748
rect 17876 7708 19372 7748
rect 19412 7708 19421 7748
rect 19555 7708 19564 7748
rect 19604 7708 20276 7748
rect 20323 7708 20332 7748
rect 20372 7708 22540 7748
rect 22580 7708 22589 7748
rect 22723 7708 22732 7748
rect 22772 7708 22781 7748
rect 23971 7708 23980 7748
rect 24020 7708 27916 7748
rect 27956 7708 27965 7748
rect 28012 7708 29644 7748
rect 29684 7708 29693 7748
rect 29827 7708 29836 7748
rect 29876 7708 33532 7748
rect 33572 7708 33581 7748
rect 33859 7708 33868 7748
rect 33908 7708 34684 7748
rect 34724 7708 34733 7748
rect 35596 7708 35836 7748
rect 35876 7708 35885 7748
rect 36595 7708 36604 7748
rect 36644 7708 36980 7748
rect 37315 7708 37324 7748
rect 37364 7708 38620 7748
rect 38660 7708 38669 7748
rect 38851 7708 38860 7748
rect 38900 7708 39004 7748
rect 39044 7708 39053 7748
rect 39523 7708 39532 7748
rect 39572 7708 39772 7748
rect 39812 7708 39821 7748
rect 22732 7664 22772 7708
rect 35596 7664 35636 7708
rect 0 7624 2900 7664
rect 3244 7624 12172 7664
rect 12212 7624 12221 7664
rect 15532 7624 22772 7664
rect 28108 7624 35636 7664
rect 36940 7664 36980 7708
rect 36940 7624 48364 7664
rect 48404 7624 48413 7664
rect 0 7604 90 7624
rect 0 7328 90 7348
rect 0 7288 1132 7328
rect 1172 7288 1181 7328
rect 0 7268 90 7288
rect 2860 7244 2900 7624
rect 28108 7580 28148 7624
rect 4919 7540 4928 7580
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 5296 7540 5305 7580
rect 17443 7540 17452 7580
rect 17492 7540 19468 7580
rect 19508 7540 19517 7580
rect 20039 7540 20048 7580
rect 20088 7540 20130 7580
rect 20170 7540 20212 7580
rect 20252 7540 20294 7580
rect 20334 7540 20376 7580
rect 20416 7540 20425 7580
rect 20524 7540 22636 7580
rect 22676 7540 22685 7580
rect 23011 7540 23020 7580
rect 23060 7540 24268 7580
rect 24308 7540 24317 7580
rect 24547 7540 24556 7580
rect 24596 7540 28148 7580
rect 28204 7540 32332 7580
rect 32372 7540 32381 7580
rect 35159 7540 35168 7580
rect 35208 7540 35250 7580
rect 35290 7540 35332 7580
rect 35372 7540 35414 7580
rect 35454 7540 35496 7580
rect 35536 7540 35545 7580
rect 36739 7540 36748 7580
rect 36788 7540 39052 7580
rect 39092 7540 39101 7580
rect 50279 7540 50288 7580
rect 50328 7540 50370 7580
rect 50410 7540 50452 7580
rect 50492 7540 50534 7580
rect 50574 7540 50616 7580
rect 50656 7540 50665 7580
rect 20524 7496 20564 7540
rect 28204 7496 28244 7540
rect 5827 7456 5836 7496
rect 5876 7456 15284 7496
rect 15244 7328 15284 7456
rect 15436 7456 20564 7496
rect 25123 7456 25132 7496
rect 25172 7456 28244 7496
rect 30019 7456 30028 7496
rect 30068 7456 33140 7496
rect 34531 7456 34540 7496
rect 34580 7456 37900 7496
rect 37940 7456 37949 7496
rect 37996 7456 41164 7496
rect 41204 7456 41213 7496
rect 15436 7328 15476 7456
rect 33100 7412 33140 7456
rect 37996 7412 38036 7456
rect 15523 7372 15532 7412
rect 15572 7372 20908 7412
rect 20948 7372 20957 7412
rect 22924 7372 26956 7412
rect 26996 7372 27005 7412
rect 27907 7372 27916 7412
rect 27956 7372 30412 7412
rect 30452 7372 30461 7412
rect 33100 7372 33772 7412
rect 33812 7372 33821 7412
rect 34627 7372 34636 7412
rect 34676 7372 38036 7412
rect 38947 7372 38956 7412
rect 38996 7372 40780 7412
rect 40820 7372 40829 7412
rect 22924 7328 22964 7372
rect 51052 7328 51092 7960
rect 53190 7940 53280 7960
rect 51667 7708 51676 7748
rect 51716 7708 51725 7748
rect 52051 7708 52060 7748
rect 52100 7708 52684 7748
rect 52724 7708 52733 7748
rect 51676 7664 51716 7708
rect 53190 7664 53280 7684
rect 51676 7624 53280 7664
rect 53190 7604 53280 7624
rect 53190 7328 53280 7348
rect 15244 7288 15476 7328
rect 16099 7288 16108 7328
rect 16148 7288 22964 7328
rect 23011 7288 23020 7328
rect 23060 7288 33868 7328
rect 33908 7288 33917 7328
rect 38956 7288 51092 7328
rect 52675 7288 52684 7328
rect 52724 7288 53280 7328
rect 38956 7244 38996 7288
rect 53190 7268 53280 7288
rect 2860 7204 18740 7244
rect 19267 7204 19276 7244
rect 19316 7204 23980 7244
rect 24020 7204 24029 7244
rect 28492 7204 28916 7244
rect 30211 7204 30220 7244
rect 30260 7204 38996 7244
rect 39100 7204 39148 7244
rect 39188 7204 39197 7244
rect 18700 7160 18740 7204
rect 28492 7160 28532 7204
rect 28876 7160 28916 7204
rect 39100 7160 39140 7204
rect 10339 7120 10348 7160
rect 10388 7120 10876 7160
rect 10916 7120 10925 7160
rect 11107 7120 11116 7160
rect 11156 7120 11287 7160
rect 11491 7120 11500 7160
rect 11540 7120 11788 7160
rect 11828 7120 11837 7160
rect 11971 7120 11980 7160
rect 12020 7120 12029 7160
rect 12521 7120 12652 7160
rect 12692 7120 12701 7160
rect 13481 7120 13612 7160
rect 13652 7120 13661 7160
rect 13987 7120 13996 7160
rect 14036 7120 14045 7160
rect 14729 7120 14860 7160
rect 14900 7120 14909 7160
rect 14995 7120 15004 7160
rect 15044 7120 15052 7160
rect 15092 7120 15175 7160
rect 15235 7120 15244 7160
rect 15284 7120 16972 7160
rect 17012 7120 17021 7160
rect 17155 7120 17164 7160
rect 17204 7120 17335 7160
rect 18700 7120 27052 7160
rect 27092 7120 27101 7160
rect 27235 7120 27244 7160
rect 27284 7120 27436 7160
rect 27476 7120 27485 7160
rect 27532 7120 28532 7160
rect 28649 7120 28780 7160
rect 28820 7120 28829 7160
rect 28876 7120 37228 7160
rect 37268 7120 37277 7160
rect 37324 7120 37372 7160
rect 37412 7120 37421 7160
rect 37651 7120 37660 7160
rect 37700 7120 37804 7160
rect 37844 7120 37853 7160
rect 37961 7120 38092 7160
rect 38132 7120 38141 7160
rect 38188 7120 38908 7160
rect 38948 7120 38957 7160
rect 39082 7120 39091 7160
rect 39131 7120 39140 7160
rect 39235 7120 39244 7160
rect 39284 7120 51436 7160
rect 51476 7120 51485 7160
rect 51689 7120 51820 7160
rect 51860 7120 51869 7160
rect 11980 7076 12020 7120
rect 13996 7076 14036 7120
rect 27532 7076 27572 7120
rect 37324 7076 37364 7120
rect 38188 7076 38228 7120
rect 9955 7036 9964 7076
rect 10004 7036 11260 7076
rect 11300 7036 11309 7076
rect 11980 7036 13652 7076
rect 13996 7036 26092 7076
rect 26132 7036 26141 7076
rect 26275 7036 26284 7076
rect 26324 7036 27572 7076
rect 28012 7036 34580 7076
rect 37315 7036 37324 7076
rect 37364 7036 37373 7076
rect 37660 7036 38228 7076
rect 38380 7036 38956 7076
rect 38996 7036 39005 7076
rect 39331 7036 39340 7076
rect 39380 7036 40972 7076
rect 41012 7036 41021 7076
rect 0 6992 90 7012
rect 0 6952 652 6992
rect 692 6952 701 6992
rect 9571 6952 9580 6992
rect 9620 6952 11740 6992
rect 11780 6952 11789 6992
rect 11884 6952 12412 6992
rect 12452 6952 12461 6992
rect 12940 6952 13372 6992
rect 13412 6952 13421 6992
rect 0 6932 90 6952
rect 11884 6908 11924 6952
rect 9187 6868 9196 6908
rect 9236 6868 11404 6908
rect 11444 6868 11453 6908
rect 11587 6868 11596 6908
rect 11636 6868 11924 6908
rect 12940 6824 12980 6952
rect 13612 6908 13652 7036
rect 13699 6952 13708 6992
rect 13748 6952 13756 6992
rect 13796 6952 13879 6992
rect 14083 6952 14092 6992
rect 14132 6952 14620 6992
rect 14660 6952 14669 6992
rect 15139 6952 15148 6992
rect 15188 6952 16924 6992
rect 16964 6952 16973 6992
rect 17059 6952 17068 6992
rect 17108 6952 26572 6992
rect 26612 6952 26621 6992
rect 27283 6952 27292 6992
rect 27332 6952 27532 6992
rect 27572 6952 27581 6992
rect 27667 6952 27676 6992
rect 27716 6952 27916 6992
rect 27956 6952 27965 6992
rect 28012 6908 28052 7036
rect 29011 6952 29020 6992
rect 29060 6952 31028 6992
rect 13612 6868 19412 6908
rect 21571 6868 21580 6908
rect 21620 6868 28052 6908
rect 3679 6784 3688 6824
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 4056 6784 4065 6824
rect 8803 6784 8812 6824
rect 8852 6784 12980 6824
rect 14851 6784 14860 6824
rect 14900 6784 18700 6824
rect 18740 6784 18749 6824
rect 18799 6784 18808 6824
rect 18848 6784 18890 6824
rect 18930 6784 18972 6824
rect 19012 6784 19054 6824
rect 19094 6784 19136 6824
rect 19176 6784 19185 6824
rect 19372 6740 19412 6868
rect 19459 6784 19468 6824
rect 19508 6784 27628 6824
rect 27668 6784 27677 6824
rect 30988 6740 31028 6952
rect 34540 6908 34580 7036
rect 37660 6908 37700 7036
rect 38380 6992 38420 7036
rect 53190 6992 53280 7012
rect 38323 6952 38332 6992
rect 38372 6952 38420 6992
rect 41155 6952 41164 6992
rect 41204 6952 47308 6992
rect 47348 6952 47357 6992
rect 51667 6952 51676 6992
rect 51716 6952 51725 6992
rect 52051 6952 52060 6992
rect 52100 6952 53280 6992
rect 34540 6868 37700 6908
rect 37795 6868 37804 6908
rect 37844 6868 47212 6908
rect 47252 6868 47261 6908
rect 33919 6784 33928 6824
rect 33968 6784 34010 6824
rect 34050 6784 34092 6824
rect 34132 6784 34174 6824
rect 34214 6784 34256 6824
rect 34296 6784 34305 6824
rect 38092 6784 47404 6824
rect 47444 6784 47453 6824
rect 49039 6784 49048 6824
rect 49088 6784 49130 6824
rect 49170 6784 49212 6824
rect 49252 6784 49294 6824
rect 49334 6784 49376 6824
rect 49416 6784 49425 6824
rect 38092 6740 38132 6784
rect 13603 6700 13612 6740
rect 13652 6700 19316 6740
rect 19372 6700 27820 6740
rect 27860 6700 27869 6740
rect 28972 6700 29260 6740
rect 29300 6700 29309 6740
rect 30988 6700 38132 6740
rect 38188 6700 40492 6740
rect 40532 6700 40541 6740
rect 0 6656 90 6676
rect 19276 6656 19316 6700
rect 28972 6656 29012 6700
rect 38188 6656 38228 6700
rect 51676 6656 51716 6952
rect 53190 6932 53280 6952
rect 53190 6656 53280 6676
rect 0 6616 940 6656
rect 980 6616 989 6656
rect 11779 6616 11788 6656
rect 11828 6616 19180 6656
rect 19220 6616 19229 6656
rect 19276 6616 23308 6656
rect 23348 6616 23357 6656
rect 23443 6616 23452 6656
rect 23492 6616 25516 6656
rect 25556 6616 25565 6656
rect 25699 6616 25708 6656
rect 25748 6616 29012 6656
rect 29059 6616 29068 6656
rect 29108 6616 37324 6656
rect 37364 6616 37373 6656
rect 38092 6616 38228 6656
rect 39859 6616 39868 6656
rect 39908 6616 48940 6656
rect 48980 6616 48989 6656
rect 49555 6616 49564 6656
rect 49604 6616 50092 6656
rect 50132 6616 50141 6656
rect 51676 6616 53280 6656
rect 0 6596 90 6616
rect 38092 6572 38132 6616
rect 53190 6596 53280 6616
rect 8419 6532 8428 6572
rect 8468 6532 14092 6572
rect 14132 6532 14141 6572
rect 15235 6532 15244 6572
rect 15284 6532 20524 6572
rect 20564 6532 20573 6572
rect 20620 6532 23404 6572
rect 23444 6532 23453 6572
rect 23500 6532 25076 6572
rect 20620 6488 20660 6532
rect 4099 6448 4108 6488
rect 4148 6448 17972 6488
rect 18691 6448 18700 6488
rect 18740 6448 20660 6488
rect 23081 6448 23212 6488
rect 23252 6448 23261 6488
rect 17932 6404 17972 6448
rect 23500 6404 23540 6532
rect 25036 6488 25076 6532
rect 25132 6532 25652 6572
rect 25843 6532 25852 6572
rect 25892 6532 38132 6572
rect 42473 6532 42556 6572
rect 42596 6532 42604 6572
rect 42644 6532 42653 6572
rect 47299 6532 47308 6572
rect 47348 6532 51476 6572
rect 23587 6448 23596 6488
rect 23636 6448 23645 6488
rect 25027 6448 25036 6488
rect 25076 6448 25085 6488
rect 17932 6364 23540 6404
rect 0 6320 90 6340
rect 23596 6320 23636 6448
rect 25132 6404 25172 6532
rect 25612 6488 25652 6532
rect 51436 6488 51476 6532
rect 25267 6448 25276 6488
rect 25316 6448 25556 6488
rect 25603 6448 25612 6488
rect 25652 6448 25661 6488
rect 26371 6448 26380 6488
rect 26420 6448 28204 6488
rect 28244 6448 28253 6488
rect 28387 6448 28396 6488
rect 28436 6448 28876 6488
rect 28916 6448 28925 6488
rect 34819 6448 34828 6488
rect 34868 6448 34877 6488
rect 39619 6448 39628 6488
rect 39668 6448 41548 6488
rect 41588 6448 41597 6488
rect 42307 6448 42316 6488
rect 42356 6448 44044 6488
rect 44084 6448 44093 6488
rect 48931 6448 48940 6488
rect 48980 6448 49324 6488
rect 49364 6448 49373 6488
rect 51427 6448 51436 6488
rect 51476 6448 51485 6488
rect 51811 6448 51820 6488
rect 51860 6448 51869 6488
rect 0 6280 1420 6320
rect 1460 6280 1469 6320
rect 6595 6280 6604 6320
rect 6644 6280 23636 6320
rect 23692 6364 25172 6404
rect 25516 6404 25556 6448
rect 25516 6364 34732 6404
rect 34772 6364 34781 6404
rect 0 6260 90 6280
rect 9091 6196 9100 6236
rect 9140 6196 23348 6236
rect 23308 6152 23348 6196
rect 23692 6152 23732 6364
rect 23827 6280 23836 6320
rect 23876 6280 33140 6320
rect 33100 6236 33140 6280
rect 25699 6196 25708 6236
rect 25748 6196 28972 6236
rect 29012 6196 29021 6236
rect 33100 6196 34732 6236
rect 34772 6196 34781 6236
rect 34828 6152 34868 6448
rect 51820 6404 51860 6448
rect 1123 6112 1132 6152
rect 1172 6112 7892 6152
rect 11587 6112 11596 6152
rect 11636 6112 23212 6152
rect 23252 6112 23261 6152
rect 23308 6112 23732 6152
rect 23779 6112 23788 6152
rect 23828 6112 26380 6152
rect 26420 6112 26429 6152
rect 26563 6112 26572 6152
rect 26612 6112 34868 6152
rect 34924 6364 51860 6404
rect 7852 6068 7892 6112
rect 34924 6068 34964 6364
rect 53190 6320 53280 6340
rect 35059 6280 35068 6320
rect 35108 6280 46828 6320
rect 46868 6280 46877 6320
rect 52051 6280 52060 6320
rect 52100 6280 53280 6320
rect 53190 6260 53280 6280
rect 35107 6196 35116 6236
rect 35156 6196 43084 6236
rect 43124 6196 43133 6236
rect 51667 6196 51676 6236
rect 51716 6196 51725 6236
rect 51676 6152 51716 6196
rect 35011 6112 35020 6152
rect 35060 6112 40588 6152
rect 40628 6112 40637 6152
rect 51676 6112 53108 6152
rect 4919 6028 4928 6068
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 5296 6028 5305 6068
rect 7852 6028 15476 6068
rect 20039 6028 20048 6068
rect 20088 6028 20130 6068
rect 20170 6028 20212 6068
rect 20252 6028 20294 6068
rect 20334 6028 20376 6068
rect 20416 6028 20425 6068
rect 20515 6028 20524 6068
rect 20564 6028 23116 6068
rect 23156 6028 23165 6068
rect 23299 6028 23308 6068
rect 23348 6028 28396 6068
rect 28436 6028 28445 6068
rect 28579 6028 28588 6068
rect 28628 6028 34964 6068
rect 35159 6028 35168 6068
rect 35208 6028 35250 6068
rect 35290 6028 35332 6068
rect 35372 6028 35414 6068
rect 35454 6028 35496 6068
rect 35536 6028 35545 6068
rect 50279 6028 50288 6068
rect 50328 6028 50370 6068
rect 50410 6028 50452 6068
rect 50492 6028 50534 6068
rect 50574 6028 50616 6068
rect 50656 6028 50665 6068
rect 0 5984 90 6004
rect 15436 5984 15476 6028
rect 53068 5984 53108 6112
rect 53190 5984 53280 6004
rect 0 5944 1036 5984
rect 1076 5944 1085 5984
rect 1219 5944 1228 5984
rect 1268 5944 15380 5984
rect 15436 5944 27244 5984
rect 27284 5944 27293 5984
rect 27523 5944 27532 5984
rect 27572 5944 47500 5984
rect 47540 5944 47549 5984
rect 47596 5944 51916 5984
rect 51956 5944 51965 5984
rect 53068 5944 53280 5984
rect 0 5924 90 5944
rect 15340 5900 15380 5944
rect 12643 5860 12652 5900
rect 12692 5860 15244 5900
rect 15284 5860 15293 5900
rect 15340 5860 28780 5900
rect 28820 5860 28829 5900
rect 28963 5860 28972 5900
rect 29012 5860 47308 5900
rect 47348 5860 47357 5900
rect 47596 5816 47636 5944
rect 53190 5924 53280 5944
rect 11107 5776 11116 5816
rect 11156 5776 27436 5816
rect 27476 5776 27485 5816
rect 27907 5776 27916 5816
rect 27956 5776 47636 5816
rect 49132 5776 51820 5816
rect 51860 5776 51869 5816
rect 49132 5732 49172 5776
rect 26371 5692 26380 5732
rect 26420 5692 29876 5732
rect 0 5648 90 5668
rect 29836 5648 29876 5692
rect 32524 5692 35444 5732
rect 38083 5692 38092 5732
rect 38132 5692 49172 5732
rect 49228 5692 51532 5732
rect 51572 5692 51581 5732
rect 32524 5648 32564 5692
rect 35404 5648 35444 5692
rect 49228 5648 49268 5692
rect 53190 5648 53280 5668
rect 0 5608 212 5648
rect 1603 5608 1612 5648
rect 1652 5608 26764 5648
rect 26804 5608 26813 5648
rect 27497 5608 27628 5648
rect 27668 5608 27677 5648
rect 29827 5608 29836 5648
rect 29876 5608 29885 5648
rect 30019 5608 30028 5648
rect 30068 5608 31660 5648
rect 31700 5608 31709 5648
rect 31891 5608 31900 5648
rect 31940 5608 32564 5648
rect 33091 5608 33100 5648
rect 33140 5608 33292 5648
rect 33332 5608 33341 5648
rect 35404 5608 41740 5648
rect 41780 5608 41789 5648
rect 46435 5608 46444 5648
rect 46484 5608 46540 5648
rect 46580 5608 46615 5648
rect 46675 5608 46684 5648
rect 46724 5608 46732 5648
rect 46772 5608 46855 5648
rect 49219 5608 49228 5648
rect 49268 5608 49277 5648
rect 49459 5608 49468 5648
rect 49508 5608 49996 5648
rect 50036 5608 50045 5648
rect 51427 5608 51436 5648
rect 51476 5608 51485 5648
rect 51689 5608 51820 5648
rect 51860 5608 51869 5648
rect 52051 5608 52060 5648
rect 52100 5608 53280 5648
rect 0 5588 90 5608
rect 172 5480 212 5608
rect 51436 5564 51476 5608
rect 53190 5588 53280 5608
rect 26995 5524 27004 5564
rect 27044 5524 40300 5564
rect 40340 5524 40349 5564
rect 40483 5524 40492 5564
rect 40532 5524 51476 5564
rect 172 5440 21964 5480
rect 22004 5440 22013 5480
rect 27859 5440 27868 5480
rect 27908 5440 29972 5480
rect 30067 5440 30076 5480
rect 30116 5440 31604 5480
rect 33091 5440 33100 5480
rect 33140 5440 33149 5480
rect 33331 5440 33340 5480
rect 33380 5440 46444 5480
rect 46484 5440 46493 5480
rect 51667 5440 51676 5480
rect 51716 5440 53108 5480
rect 76 5356 2900 5396
rect 16579 5356 16588 5396
rect 16628 5356 29836 5396
rect 29876 5356 29885 5396
rect 76 5332 116 5356
rect 0 5272 116 5332
rect 0 5252 90 5272
rect 2860 5144 2900 5356
rect 3679 5272 3688 5312
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 4056 5272 4065 5312
rect 18799 5272 18808 5312
rect 18848 5272 18890 5312
rect 18930 5272 18972 5312
rect 19012 5272 19054 5312
rect 19094 5272 19136 5312
rect 19176 5272 19185 5312
rect 29932 5228 29972 5440
rect 31564 5396 31604 5440
rect 33100 5396 33140 5440
rect 31564 5356 33140 5396
rect 53068 5312 53108 5440
rect 53190 5312 53280 5332
rect 30115 5272 30124 5312
rect 30164 5272 33292 5312
rect 33332 5272 33341 5312
rect 33919 5272 33928 5312
rect 33968 5272 34010 5312
rect 34050 5272 34092 5312
rect 34132 5272 34174 5312
rect 34214 5272 34256 5312
rect 34296 5272 34305 5312
rect 49039 5272 49048 5312
rect 49088 5272 49130 5312
rect 49170 5272 49212 5312
rect 49252 5272 49294 5312
rect 49334 5272 49376 5312
rect 49416 5272 49425 5312
rect 53068 5272 53280 5312
rect 53190 5252 53280 5272
rect 14083 5188 14092 5228
rect 14132 5188 26380 5228
rect 26420 5188 26429 5228
rect 29932 5188 38092 5228
rect 38132 5188 38141 5228
rect 2860 5104 21772 5144
rect 21812 5104 21821 5144
rect 22051 5104 22060 5144
rect 22100 5104 26764 5144
rect 26804 5104 26813 5144
rect 33187 5104 33196 5144
rect 33236 5104 44236 5144
rect 44276 5104 44285 5144
rect 643 5020 652 5060
rect 692 5020 27628 5060
rect 27668 5020 27677 5060
rect 31987 5020 31996 5060
rect 32036 5020 41836 5060
rect 41876 5020 41885 5060
rect 43180 5020 51860 5060
rect 0 4976 90 4996
rect 43180 4976 43220 5020
rect 51820 4976 51860 5020
rect 53190 4976 53280 4996
rect 0 4936 21580 4976
rect 21620 4936 21629 4976
rect 23020 4936 31756 4976
rect 31796 4936 31805 4976
rect 32297 4936 32428 4976
rect 32468 4936 32477 4976
rect 32611 4936 32620 4976
rect 32660 4936 43220 4976
rect 51427 4936 51436 4976
rect 51476 4936 51485 4976
rect 51811 4936 51820 4976
rect 51860 4936 51869 4976
rect 52051 4936 52060 4976
rect 52100 4936 53280 4976
rect 0 4916 90 4936
rect 23020 4808 23060 4936
rect 51436 4892 51476 4936
rect 53190 4916 53280 4936
rect 25507 4852 25516 4892
rect 25556 4852 51476 4892
rect 19267 4768 19276 4808
rect 19316 4768 23060 4808
rect 26755 4768 26764 4808
rect 26804 4768 40492 4808
rect 40532 4768 40541 4808
rect 47500 4768 51820 4808
rect 51860 4768 51869 4808
rect 23971 4684 23980 4724
rect 24020 4684 30124 4724
rect 30164 4684 30173 4724
rect 32659 4684 32668 4724
rect 32708 4684 46060 4724
rect 46100 4684 46109 4724
rect 0 4640 90 4660
rect 47500 4640 47540 4768
rect 51667 4684 51676 4724
rect 51716 4684 51725 4724
rect 0 4600 22348 4640
rect 22388 4600 22397 4640
rect 33100 4600 47540 4640
rect 51676 4640 51716 4684
rect 53190 4640 53280 4660
rect 51676 4600 53280 4640
rect 0 4580 90 4600
rect 4919 4516 4928 4556
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 5296 4516 5305 4556
rect 20039 4516 20048 4556
rect 20088 4516 20130 4556
rect 20170 4516 20212 4556
rect 20252 4516 20294 4556
rect 20334 4516 20376 4556
rect 20416 4516 20425 4556
rect 21667 4516 21676 4556
rect 21716 4516 32428 4556
rect 32468 4516 32477 4556
rect 33100 4472 33140 4600
rect 53190 4580 53280 4600
rect 35159 4516 35168 4556
rect 35208 4516 35250 4556
rect 35290 4516 35332 4556
rect 35372 4516 35414 4556
rect 35454 4516 35496 4556
rect 35536 4516 35545 4556
rect 50279 4516 50288 4556
rect 50328 4516 50370 4556
rect 50410 4516 50452 4556
rect 50492 4516 50534 4556
rect 50574 4516 50616 4556
rect 50656 4516 50665 4556
rect 23491 4432 23500 4472
rect 23540 4432 33140 4472
rect 24739 4348 24748 4388
rect 24788 4348 32620 4388
rect 32660 4348 32669 4388
rect 0 4304 90 4324
rect 53190 4304 53280 4324
rect 0 4264 24500 4304
rect 25459 4264 25468 4304
rect 25508 4264 31316 4304
rect 52051 4264 52060 4304
rect 52100 4264 53280 4304
rect 0 4244 90 4264
rect 19843 4180 19852 4220
rect 19892 4180 22964 4220
rect 22924 4136 22964 4180
rect 24460 4136 24500 4264
rect 24940 4180 31180 4220
rect 31220 4180 31229 4220
rect 17923 4096 17932 4136
rect 17972 4096 20620 4136
rect 20660 4096 20669 4136
rect 21667 4096 21676 4136
rect 21716 4096 21725 4136
rect 22051 4096 22060 4136
rect 22100 4096 22109 4136
rect 22156 4096 22540 4136
rect 22580 4096 22589 4136
rect 22915 4096 22924 4136
rect 22964 4096 22973 4136
rect 23177 4096 23308 4136
rect 23348 4096 23357 4136
rect 23945 4096 24076 4136
rect 24116 4096 24125 4136
rect 24451 4096 24460 4136
rect 24500 4096 24509 4136
rect 24643 4096 24652 4136
rect 24692 4096 24844 4136
rect 24884 4096 24893 4136
rect 21676 4052 21716 4096
rect 19459 4012 19468 4052
rect 19508 4012 21716 4052
rect 0 3968 90 3988
rect 0 3928 7852 3968
rect 7892 3928 7901 3968
rect 20851 3928 20860 3968
rect 20900 3928 21484 3968
rect 21524 3928 21533 3968
rect 21785 3928 21868 3968
rect 21908 3928 21916 3968
rect 21956 3928 21965 3968
rect 0 3908 90 3928
rect 22060 3884 22100 4096
rect 2860 3844 22100 3884
rect 0 3632 90 3652
rect 2860 3632 2900 3844
rect 3679 3760 3688 3800
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 4056 3760 4065 3800
rect 18799 3760 18808 3800
rect 18848 3760 18890 3800
rect 18930 3760 18972 3800
rect 19012 3760 19054 3800
rect 19094 3760 19136 3800
rect 19176 3760 19185 3800
rect 22156 3716 22196 4096
rect 24940 4052 24980 4180
rect 31276 4136 31316 4264
rect 53190 4244 53280 4264
rect 31363 4180 31372 4220
rect 31412 4180 51820 4220
rect 51860 4180 51869 4220
rect 25097 4096 25228 4136
rect 25268 4096 25277 4136
rect 25481 4096 25612 4136
rect 25652 4096 25661 4136
rect 25865 4096 25996 4136
rect 26036 4096 26045 4136
rect 26153 4096 26236 4136
rect 26276 4096 26284 4136
rect 26324 4096 26333 4136
rect 31276 4096 47308 4136
rect 47348 4096 47357 4136
rect 51427 4096 51436 4136
rect 51476 4096 51485 4136
rect 51532 4096 51820 4136
rect 51860 4096 51869 4136
rect 51436 4052 51476 4096
rect 22291 4012 22300 4052
rect 22340 4012 24980 4052
rect 25075 4012 25084 4052
rect 25124 4012 51476 4052
rect 22771 3928 22780 3968
rect 22820 3928 22924 3968
rect 22964 3928 22973 3968
rect 23155 3928 23164 3968
rect 23204 3928 23404 3968
rect 23444 3928 23453 3968
rect 23539 3928 23548 3968
rect 23588 3928 24172 3968
rect 24212 3928 24221 3968
rect 24307 3928 24316 3968
rect 24356 3928 24460 3968
rect 24500 3928 24509 3968
rect 24691 3928 24700 3968
rect 24740 3928 25364 3968
rect 25843 3928 25852 3968
rect 25892 3928 25900 3968
rect 25940 3928 26023 3968
rect 25324 3884 25364 3928
rect 51532 3884 51572 4096
rect 51667 4012 51676 4052
rect 51716 4012 52628 4052
rect 52588 3968 52628 4012
rect 53190 3968 53280 3988
rect 52588 3928 53280 3968
rect 53190 3908 53280 3928
rect 25324 3844 51572 3884
rect 33919 3760 33928 3800
rect 33968 3760 34010 3800
rect 34050 3760 34092 3800
rect 34132 3760 34174 3800
rect 34214 3760 34256 3800
rect 34296 3760 34305 3800
rect 49039 3760 49048 3800
rect 49088 3760 49130 3800
rect 49170 3760 49212 3800
rect 49252 3760 49294 3800
rect 49334 3760 49376 3800
rect 49416 3760 49425 3800
rect 18115 3676 18124 3716
rect 18164 3676 22196 3716
rect 23203 3676 23212 3716
rect 23252 3676 25228 3716
rect 25268 3676 25277 3716
rect 53190 3632 53280 3652
rect 0 3592 2900 3632
rect 21929 3592 22012 3632
rect 22052 3592 22060 3632
rect 22100 3592 22109 3632
rect 23347 3592 23356 3632
rect 23396 3592 23500 3632
rect 23540 3592 23549 3632
rect 24499 3592 24508 3632
rect 24548 3592 24748 3632
rect 24788 3592 24797 3632
rect 25385 3592 25468 3632
rect 25508 3592 25516 3632
rect 25556 3592 25565 3632
rect 28457 3592 28540 3632
rect 28580 3592 28588 3632
rect 28628 3592 28637 3632
rect 52051 3592 52060 3632
rect 52100 3592 53280 3632
rect 0 3572 90 3592
rect 53190 3572 53280 3592
rect 21571 3508 21580 3548
rect 21620 3508 24308 3548
rect 24547 3508 24556 3548
rect 24596 3508 25612 3548
rect 25652 3508 25661 3548
rect 24268 3464 24308 3508
rect 21641 3424 21772 3464
rect 21812 3424 21821 3464
rect 21955 3424 21964 3464
rect 22004 3424 23116 3464
rect 23156 3424 23165 3464
rect 24259 3424 24268 3464
rect 24308 3424 24317 3464
rect 24713 3424 24844 3464
rect 24884 3424 24893 3464
rect 25219 3424 25228 3464
rect 25268 3424 25277 3464
rect 28169 3424 28300 3464
rect 28340 3424 28349 3464
rect 47299 3424 47308 3464
rect 47348 3424 51436 3464
rect 51476 3424 51485 3464
rect 51689 3424 51820 3464
rect 51860 3424 51869 3464
rect 25228 3380 25268 3424
rect 7843 3340 7852 3380
rect 7892 3340 22292 3380
rect 22339 3340 22348 3380
rect 22388 3340 25268 3380
rect 0 3296 90 3316
rect 22252 3296 22292 3340
rect 53190 3296 53280 3316
rect 0 3256 22196 3296
rect 22252 3256 24652 3296
rect 24692 3256 24701 3296
rect 51667 3256 51676 3296
rect 51716 3256 53280 3296
rect 0 3236 90 3256
rect 22156 3212 22196 3256
rect 53190 3236 53280 3256
rect 22156 3172 23212 3212
rect 23252 3172 23261 3212
rect 25075 3172 25084 3212
rect 25124 3172 25324 3212
rect 25364 3172 25373 3212
rect 18307 3088 18316 3128
rect 18356 3088 23308 3128
rect 23348 3088 23357 3128
rect 4919 3004 4928 3044
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 5296 3004 5305 3044
rect 20039 3004 20048 3044
rect 20088 3004 20130 3044
rect 20170 3004 20212 3044
rect 20252 3004 20294 3044
rect 20334 3004 20376 3044
rect 20416 3004 20425 3044
rect 35159 3004 35168 3044
rect 35208 3004 35250 3044
rect 35290 3004 35332 3044
rect 35372 3004 35414 3044
rect 35454 3004 35496 3044
rect 35536 3004 35545 3044
rect 50279 3004 50288 3044
rect 50328 3004 50370 3044
rect 50410 3004 50452 3044
rect 50492 3004 50534 3044
rect 50574 3004 50616 3044
rect 50656 3004 50665 3044
rect 0 2960 90 2980
rect 53190 2960 53280 2980
rect 0 2920 24076 2960
rect 24116 2920 24125 2960
rect 52684 2920 53280 2960
rect 0 2900 90 2920
rect 52684 2876 52724 2920
rect 53190 2900 53280 2920
rect 25459 2836 25468 2876
rect 25508 2836 25708 2876
rect 25748 2836 25757 2876
rect 52051 2836 52060 2876
rect 52100 2836 52724 2876
rect 172 2752 24844 2792
rect 24884 2752 24893 2792
rect 25315 2752 25324 2792
rect 25364 2752 51476 2792
rect 0 2624 90 2644
rect 0 2564 116 2624
rect 76 2540 116 2564
rect 172 2540 212 2752
rect 24451 2668 24460 2708
rect 24500 2668 51188 2708
rect 76 2500 212 2540
rect 7180 2584 24556 2624
rect 24596 2584 24605 2624
rect 25219 2584 25228 2624
rect 25268 2584 25277 2624
rect 25324 2584 51052 2624
rect 51092 2584 51101 2624
rect 7180 2456 7220 2584
rect 25228 2456 25268 2584
rect 172 2416 7220 2456
rect 17260 2416 25268 2456
rect 0 2288 90 2308
rect 172 2288 212 2416
rect 17260 2372 17300 2416
rect 1027 2332 1036 2372
rect 1076 2332 17300 2372
rect 25324 2288 25364 2584
rect 51148 2540 51188 2668
rect 51436 2624 51476 2752
rect 53190 2624 53280 2644
rect 51427 2584 51436 2624
rect 51476 2584 51485 2624
rect 51532 2584 51820 2624
rect 51860 2584 51869 2624
rect 52588 2584 53280 2624
rect 51532 2540 51572 2584
rect 52588 2540 52628 2584
rect 53190 2564 53280 2584
rect 51148 2500 51572 2540
rect 51667 2500 51676 2540
rect 51716 2500 52628 2540
rect 51283 2416 51292 2456
rect 51332 2416 51956 2456
rect 0 2248 212 2288
rect 3679 2248 3688 2288
rect 3728 2248 3770 2288
rect 3810 2248 3852 2288
rect 3892 2248 3934 2288
rect 3974 2248 4016 2288
rect 4056 2248 4065 2288
rect 18799 2248 18808 2288
rect 18848 2248 18890 2288
rect 18930 2248 18972 2288
rect 19012 2248 19054 2288
rect 19094 2248 19136 2288
rect 19176 2248 19185 2288
rect 21859 2248 21868 2288
rect 21908 2248 25364 2288
rect 25420 2332 50380 2372
rect 50420 2332 50429 2372
rect 0 2228 90 2248
rect 25420 2204 25460 2332
rect 33919 2248 33928 2288
rect 33968 2248 34010 2288
rect 34050 2248 34092 2288
rect 34132 2248 34174 2288
rect 34214 2248 34256 2288
rect 34296 2248 34305 2288
rect 49039 2248 49048 2288
rect 49088 2248 49130 2288
rect 49170 2248 49212 2288
rect 49252 2248 49294 2288
rect 49334 2248 49376 2288
rect 49416 2248 49425 2288
rect 49516 2248 51860 2288
rect 49516 2204 49556 2248
rect 24163 2164 24172 2204
rect 24212 2164 25460 2204
rect 25891 2164 25900 2204
rect 25940 2164 49556 2204
rect 23395 2080 23404 2120
rect 23444 2080 50420 2120
rect 50380 2036 50420 2080
rect 23107 1996 23116 2036
rect 23156 1996 45292 2036
rect 45332 1996 45341 2036
rect 50380 1996 51476 2036
rect 0 1952 90 1972
rect 51436 1952 51476 1996
rect 51820 1952 51860 2248
rect 51916 1952 51956 2416
rect 53190 2288 53280 2308
rect 52492 2248 53280 2288
rect 52492 2120 52532 2248
rect 53190 2228 53280 2248
rect 52051 2080 52060 2120
rect 52100 2080 52532 2120
rect 53190 1952 53280 1972
rect 0 1912 19468 1952
rect 19508 1912 19517 1952
rect 21475 1912 21484 1952
rect 21524 1912 23060 1952
rect 50314 1912 50323 1952
rect 50363 1912 50380 1952
rect 50420 1912 50503 1952
rect 50659 1912 50668 1952
rect 50708 1912 50717 1952
rect 50764 1912 51052 1952
rect 51092 1912 51101 1952
rect 51283 1912 51292 1952
rect 51332 1912 51380 1952
rect 51427 1912 51436 1952
rect 51476 1912 51485 1952
rect 51811 1912 51820 1952
rect 51860 1912 51869 1952
rect 51916 1912 53280 1952
rect 0 1892 90 1912
rect 23020 1868 23060 1912
rect 23020 1828 43084 1868
rect 43124 1828 43133 1868
rect 43267 1828 43276 1868
rect 43316 1828 50572 1868
rect 50612 1828 50621 1868
rect 50668 1784 50708 1912
rect 50764 1868 50804 1912
rect 51340 1868 51380 1912
rect 53190 1892 53280 1912
rect 50755 1828 50764 1868
rect 50804 1828 50813 1868
rect 51340 1828 52300 1868
rect 52340 1828 52349 1868
rect 45283 1744 45292 1784
rect 45332 1744 50708 1784
rect 50899 1744 50908 1784
rect 50948 1744 52972 1784
rect 53012 1744 53021 1784
rect 50515 1660 50524 1700
rect 50564 1660 51572 1700
rect 51667 1660 51676 1700
rect 51716 1660 51725 1700
rect 0 1616 90 1636
rect 0 1576 19852 1616
rect 19892 1576 19901 1616
rect 0 1556 90 1576
rect 51532 1532 51572 1660
rect 51676 1616 51716 1660
rect 53190 1616 53280 1636
rect 51676 1576 53280 1616
rect 53190 1556 53280 1576
rect 4919 1492 4928 1532
rect 4968 1492 5010 1532
rect 5050 1492 5092 1532
rect 5132 1492 5174 1532
rect 5214 1492 5256 1532
rect 5296 1492 5305 1532
rect 20039 1492 20048 1532
rect 20088 1492 20130 1532
rect 20170 1492 20212 1532
rect 20252 1492 20294 1532
rect 20334 1492 20376 1532
rect 20416 1492 20425 1532
rect 35159 1492 35168 1532
rect 35208 1492 35250 1532
rect 35290 1492 35332 1532
rect 35372 1492 35414 1532
rect 35454 1492 35496 1532
rect 35536 1492 35545 1532
rect 50279 1492 50288 1532
rect 50328 1492 50370 1532
rect 50410 1492 50452 1532
rect 50492 1492 50534 1532
rect 50574 1492 50616 1532
rect 50656 1492 50665 1532
rect 51532 1492 52532 1532
rect 52492 1448 52532 1492
rect 52492 1408 53164 1448
rect 53204 1408 53213 1448
rect 0 1280 90 1300
rect 53190 1280 53280 1300
rect 0 1240 18316 1280
rect 18356 1240 18365 1280
rect 53155 1240 53164 1280
rect 53204 1240 53280 1280
rect 0 1220 90 1240
rect 53190 1220 53280 1240
rect 0 944 90 964
rect 53190 944 53280 964
rect 0 904 18124 944
rect 18164 904 18173 944
rect 52963 904 52972 944
rect 53012 904 53280 944
rect 0 884 90 904
rect 53190 884 53280 904
rect 0 608 90 628
rect 53190 608 53280 628
rect 0 568 17932 608
rect 17972 568 17981 608
rect 52291 568 52300 608
rect 52340 568 53280 608
rect 0 548 90 568
rect 53190 548 53280 568
<< via2 >>
rect 17164 11740 17204 11780
rect 31948 11740 31988 11780
rect 17260 11656 17300 11696
rect 31564 11656 31604 11696
rect 19372 11572 19412 11612
rect 32716 11572 32756 11612
rect 19564 11488 19604 11528
rect 31180 11488 31220 11528
rect 19852 11404 19892 11444
rect 30796 11404 30836 11444
rect 16684 11152 16724 11192
rect 25036 11152 25076 11192
rect 748 10984 788 11024
rect 50860 10984 50900 11024
rect 556 10648 596 10688
rect 50764 10648 50804 10688
rect 1228 10312 1268 10352
rect 52300 10312 52340 10352
rect 18028 10228 18068 10268
rect 24652 10228 24692 10268
rect 23116 10144 23156 10184
rect 23308 10060 23348 10100
rect 35788 10060 35828 10100
rect 1420 9976 1460 10016
rect 8620 9976 8660 10016
rect 3688 9808 3728 9848
rect 3770 9808 3810 9848
rect 3852 9808 3892 9848
rect 3934 9808 3974 9848
rect 4016 9808 4056 9848
rect 10636 9724 10676 9764
rect 2764 9640 2804 9680
rect 3148 9640 3188 9680
rect 3532 9640 3572 9680
rect 4108 9640 4148 9680
rect 4300 9640 4340 9680
rect 4684 9640 4724 9680
rect 5068 9640 5108 9680
rect 5452 9640 5492 9680
rect 5836 9640 5876 9680
rect 6220 9640 6260 9680
rect 6604 9640 6644 9680
rect 6988 9640 7028 9680
rect 7372 9640 7412 9680
rect 7756 9640 7796 9680
rect 8140 9640 8180 9680
rect 8524 9640 8564 9680
rect 8908 9640 8948 9680
rect 9292 9640 9332 9680
rect 9676 9640 9716 9680
rect 10060 9640 10100 9680
rect 10444 9640 10484 9680
rect 7180 9556 7220 9596
rect 16012 9976 16052 10016
rect 16300 9976 16340 10016
rect 19468 9976 19508 10016
rect 28588 9976 28628 10016
rect 50956 9976 50996 10016
rect 51148 9976 51188 10016
rect 10828 9640 10868 9680
rect 13228 9892 13268 9932
rect 13804 9892 13844 9932
rect 14188 9892 14228 9932
rect 22828 9892 22868 9932
rect 25516 9892 25556 9932
rect 11212 9640 11252 9680
rect 4108 9472 4148 9512
rect 4588 9472 4628 9512
rect 5356 9472 5396 9512
rect 6892 9472 6932 9512
rect 7084 9472 7124 9512
rect 8044 9472 8084 9512
rect 8428 9472 8468 9512
rect 8812 9472 8852 9512
rect 9196 9472 9236 9512
rect 9580 9472 9620 9512
rect 9964 9472 10004 9512
rect 10348 9472 10388 9512
rect 4300 9388 4340 9428
rect 5644 9388 5684 9428
rect 6028 9388 6068 9428
rect 18412 9808 18452 9848
rect 18808 9808 18848 9848
rect 18890 9808 18930 9848
rect 18972 9808 19012 9848
rect 19054 9808 19094 9848
rect 19136 9808 19176 9848
rect 19468 9808 19508 9848
rect 22444 9808 22484 9848
rect 31180 9808 31220 9848
rect 33928 9808 33968 9848
rect 34010 9808 34050 9848
rect 34092 9808 34132 9848
rect 34174 9808 34214 9848
rect 34256 9808 34296 9848
rect 11596 9640 11636 9680
rect 11980 9640 12020 9680
rect 12364 9640 12404 9680
rect 12748 9640 12788 9680
rect 13132 9640 13172 9680
rect 13324 9556 13364 9596
rect 18316 9724 18356 9764
rect 20140 9724 20180 9764
rect 20332 9724 20372 9764
rect 34636 9724 34676 9764
rect 13516 9640 13556 9680
rect 13900 9640 13940 9680
rect 14284 9640 14324 9680
rect 14668 9640 14708 9680
rect 15052 9640 15092 9680
rect 15436 9640 15476 9680
rect 15820 9640 15860 9680
rect 16204 9640 16244 9680
rect 16588 9640 16628 9680
rect 16972 9640 17012 9680
rect 17356 9640 17396 9680
rect 17740 9640 17780 9680
rect 18124 9640 18164 9680
rect 18508 9640 18548 9680
rect 17932 9556 17972 9596
rect 18700 9556 18740 9596
rect 19276 9640 19316 9680
rect 19660 9640 19700 9680
rect 20044 9640 20084 9680
rect 20428 9640 20468 9680
rect 20812 9640 20852 9680
rect 21196 9640 21236 9680
rect 21580 9640 21620 9680
rect 21964 9640 22004 9680
rect 22348 9640 22388 9680
rect 22636 9640 22676 9680
rect 23884 9640 23924 9680
rect 36172 9640 36212 9680
rect 42700 9640 42740 9680
rect 43084 9640 43124 9680
rect 43468 9640 43508 9680
rect 43852 9640 43892 9680
rect 44236 9640 44276 9680
rect 20620 9556 20660 9596
rect 21772 9556 21812 9596
rect 28780 9556 28820 9596
rect 49048 9808 49088 9848
rect 49130 9808 49170 9848
rect 49212 9808 49252 9848
rect 49294 9808 49334 9848
rect 49376 9808 49416 9848
rect 47116 9724 47156 9764
rect 44620 9640 44660 9680
rect 45004 9640 45044 9680
rect 45388 9640 45428 9680
rect 45772 9640 45812 9680
rect 46156 9640 46196 9680
rect 46540 9640 46580 9680
rect 46924 9640 46964 9680
rect 47308 9640 47348 9680
rect 47692 9640 47732 9680
rect 48076 9640 48116 9680
rect 48460 9640 48500 9680
rect 48844 9640 48884 9680
rect 49516 9640 49556 9680
rect 49996 9640 50036 9680
rect 50380 9640 50420 9680
rect 49612 9556 49652 9596
rect 11116 9472 11156 9512
rect 12652 9472 12692 9512
rect 13228 9472 13268 9512
rect 15148 9472 15188 9512
rect 15916 9472 15956 9512
rect 18604 9472 18644 9512
rect 19948 9472 19988 9512
rect 20524 9472 20564 9512
rect 21292 9472 21332 9512
rect 21676 9472 21716 9512
rect 22348 9472 22388 9512
rect 23020 9472 23060 9512
rect 36940 9472 36980 9512
rect 40300 9472 40340 9512
rect 46060 9472 46100 9512
rect 46444 9472 46484 9512
rect 46828 9472 46868 9512
rect 47212 9472 47252 9512
rect 47404 9472 47444 9512
rect 47980 9472 48020 9512
rect 48364 9472 48404 9512
rect 48748 9472 48788 9512
rect 49036 9472 49076 9512
rect 50092 9472 50132 9512
rect 7756 9388 7796 9428
rect 268 9304 308 9344
rect 10156 9304 10196 9344
rect 16396 9388 16436 9428
rect 16300 9304 16340 9344
rect 17836 9388 17876 9428
rect 19084 9388 19124 9428
rect 19276 9388 19316 9428
rect 22252 9388 22292 9428
rect 24940 9388 24980 9428
rect 32716 9388 32756 9428
rect 40588 9388 40628 9428
rect 43180 9388 43220 9428
rect 44236 9388 44276 9428
rect 18988 9304 19028 9344
rect 22156 9304 22196 9344
rect 22348 9304 22388 9344
rect 24844 9304 24884 9344
rect 35020 9304 35060 9344
rect 40492 9304 40532 9344
rect 20140 9220 20180 9260
rect 22924 9220 22964 9260
rect 35404 9220 35444 9260
rect 41740 9220 41780 9260
rect 8044 9136 8084 9176
rect 12940 9136 12980 9176
rect 18700 9136 18740 9176
rect 19084 9136 19124 9176
rect 19660 9136 19700 9176
rect 19948 9136 19988 9176
rect 22732 9136 22772 9176
rect 27724 9136 27764 9176
rect 31468 9136 31508 9176
rect 41836 9136 41876 9176
rect 49996 9388 50036 9428
rect 46732 9304 46772 9344
rect 51052 9472 51092 9512
rect 4928 9052 4968 9092
rect 5010 9052 5050 9092
rect 5092 9052 5132 9092
rect 5174 9052 5214 9092
rect 5256 9052 5296 9092
rect 6028 9052 6068 9092
rect 11500 9052 11540 9092
rect 15052 9052 15092 9092
rect 17548 9052 17588 9092
rect 20048 9052 20088 9092
rect 20130 9052 20170 9092
rect 20212 9052 20252 9092
rect 20294 9052 20334 9092
rect 20376 9052 20416 9092
rect 20620 9052 20660 9092
rect 24172 9052 24212 9092
rect 30220 9052 30260 9092
rect 31084 9052 31124 9092
rect 35168 9052 35208 9092
rect 35250 9052 35290 9092
rect 35332 9052 35372 9092
rect 35414 9052 35454 9092
rect 35496 9052 35536 9092
rect 37996 9052 38036 9092
rect 42316 9052 42356 9092
rect 42604 9052 42644 9092
rect 11596 8968 11636 9008
rect 11788 8968 11828 9008
rect 17452 8968 17492 9008
rect 18604 8968 18644 9008
rect 19756 8968 19796 9008
rect 21484 8968 21524 9008
rect 23116 8968 23156 9008
rect 29356 8968 29396 9008
rect 30988 8968 31028 9008
rect 31372 8968 31412 9008
rect 50188 9052 50228 9092
rect 50288 9052 50328 9092
rect 50370 9052 50410 9092
rect 50452 9052 50492 9092
rect 50534 9052 50574 9092
rect 50616 9052 50656 9092
rect 5644 8884 5684 8924
rect 13708 8884 13748 8924
rect 13900 8884 13940 8924
rect 20236 8884 20276 8924
rect 20716 8884 20756 8924
rect 22156 8884 22196 8924
rect 22636 8884 22676 8924
rect 22828 8884 22868 8924
rect 31276 8884 31316 8924
rect 31468 8884 31508 8924
rect 50860 8968 50900 9008
rect 52684 9220 52724 9260
rect 50764 8884 50804 8924
rect 51052 8884 51092 8924
rect 5356 8800 5396 8840
rect 13324 8800 13364 8840
rect 17836 8800 17876 8840
rect 13228 8716 13268 8756
rect 20140 8716 20180 8756
rect 24844 8716 24884 8756
rect 25036 8716 25076 8756
rect 28588 8716 28628 8756
rect 47116 8800 47156 8840
rect 47404 8800 47444 8840
rect 1420 8632 1460 8672
rect 12652 8632 12692 8672
rect 20716 8632 20756 8672
rect 21868 8632 21908 8672
rect 22732 8632 22772 8672
rect 23308 8632 23348 8672
rect 23884 8632 23924 8672
rect 26764 8632 26804 8672
rect 27148 8632 27188 8672
rect 27532 8632 27572 8672
rect 27724 8632 27764 8672
rect 28012 8632 28052 8672
rect 29068 8632 29108 8672
rect 29452 8632 29492 8672
rect 31180 8632 31220 8672
rect 37996 8632 38036 8672
rect 38188 8632 38228 8672
rect 50284 8632 50324 8672
rect 50956 8632 50996 8672
rect 51436 8632 51476 8672
rect 52684 8632 52724 8672
rect 6124 8548 6164 8588
rect 18028 8548 18068 8588
rect 18604 8548 18644 8588
rect 25228 8548 25268 8588
rect 30220 8548 30260 8588
rect 35308 8548 35348 8588
rect 40396 8548 40436 8588
rect 15820 8464 15860 8504
rect 17068 8464 17108 8504
rect 18220 8464 18260 8504
rect 19852 8464 19892 8504
rect 20044 8464 20084 8504
rect 20332 8464 20372 8504
rect 21484 8464 21524 8504
rect 22444 8464 22484 8504
rect 22924 8464 22964 8504
rect 31084 8464 31124 8504
rect 32908 8464 32948 8504
rect 37132 8464 37172 8504
rect 37612 8464 37652 8504
rect 40012 8464 40052 8504
rect 52684 8464 52724 8504
rect 10060 8380 10100 8420
rect 15916 8380 15956 8420
rect 16300 8380 16340 8420
rect 16780 8380 16820 8420
rect 23500 8380 23540 8420
rect 24172 8380 24212 8420
rect 32812 8380 32852 8420
rect 37804 8380 37844 8420
rect 39628 8380 39668 8420
rect 3688 8296 3728 8336
rect 3770 8296 3810 8336
rect 3852 8296 3892 8336
rect 3934 8296 3974 8336
rect 4016 8296 4056 8336
rect 4108 8128 4148 8168
rect 4300 8128 4340 8168
rect 10252 8296 10292 8336
rect 18808 8296 18848 8336
rect 18890 8296 18930 8336
rect 18972 8296 19012 8336
rect 19054 8296 19094 8336
rect 19136 8296 19176 8336
rect 20140 8296 20180 8336
rect 20332 8296 20372 8336
rect 31852 8296 31892 8336
rect 33928 8296 33968 8336
rect 34010 8296 34050 8336
rect 34092 8296 34132 8336
rect 34174 8296 34214 8336
rect 34256 8296 34296 8336
rect 37708 8296 37748 8336
rect 39052 8296 39092 8336
rect 39340 8296 39380 8336
rect 41548 8296 41588 8336
rect 49048 8296 49088 8336
rect 49130 8296 49170 8336
rect 49212 8296 49252 8336
rect 49294 8296 49334 8336
rect 49376 8296 49416 8336
rect 6892 8128 6932 8168
rect 7756 8128 7796 8168
rect 7084 8044 7124 8084
rect 10156 8128 10196 8168
rect 12844 8128 12884 8168
rect 13036 8128 13076 8168
rect 15628 8128 15668 8168
rect 16012 8128 16052 8168
rect 16396 8128 16436 8168
rect 16780 8128 16820 8168
rect 17260 8128 17300 8168
rect 17548 8128 17588 8168
rect 17932 8128 17972 8168
rect 18316 8128 18356 8168
rect 18700 8128 18740 8168
rect 10252 8044 10292 8084
rect 11500 8044 11540 8084
rect 12172 8044 12212 8084
rect 1228 7960 1268 8000
rect 5836 7960 5876 8000
rect 6124 7960 6164 8000
rect 10636 7960 10676 8000
rect 15340 7960 15380 8000
rect 10060 7876 10100 7916
rect 15436 7876 15476 7916
rect 7180 7792 7220 7832
rect 17068 8044 17108 8084
rect 18412 8044 18452 8084
rect 25132 8212 25172 8252
rect 25324 8212 25364 8252
rect 35404 8212 35444 8252
rect 47980 8212 48020 8252
rect 16108 7960 16148 8000
rect 17452 7960 17492 8000
rect 17836 7960 17876 8000
rect 18220 7960 18260 8000
rect 18604 7960 18644 8000
rect 19276 7960 19316 8000
rect 20716 8128 20756 8168
rect 25036 8128 25076 8168
rect 30028 8128 30068 8168
rect 32716 8128 32756 8168
rect 36556 8128 36596 8168
rect 36940 8128 36980 8168
rect 37420 8128 37460 8168
rect 37900 8128 37940 8168
rect 38860 8128 38900 8168
rect 52300 8128 52340 8168
rect 20236 8044 20276 8084
rect 28492 8044 28532 8084
rect 33292 8044 33332 8084
rect 33484 8044 33524 8084
rect 37612 8044 37652 8084
rect 37804 8044 37844 8084
rect 39244 8044 39284 8084
rect 39436 8044 39476 8084
rect 39724 8044 39764 8084
rect 41932 8044 41972 8084
rect 47500 8044 47540 8084
rect 21004 7960 21044 8000
rect 21196 7960 21236 8000
rect 22540 7960 22580 8000
rect 22732 7960 22772 8000
rect 28396 7960 28436 8000
rect 28588 7960 28628 8000
rect 28972 7960 29012 8000
rect 33196 7960 33236 8000
rect 33580 7960 33620 8000
rect 34636 7960 34676 8000
rect 34924 7960 34964 8000
rect 35308 7960 35348 8000
rect 36556 7960 36596 8000
rect 36748 7960 36788 8000
rect 37228 7960 37268 8000
rect 38380 7960 38420 8000
rect 39052 7960 39092 8000
rect 51916 7960 51956 8000
rect 52684 7960 52724 8000
rect 25036 7876 25076 7916
rect 28780 7876 28820 7916
rect 39628 7876 39668 7916
rect 23212 7792 23252 7832
rect 28108 7792 28148 7832
rect 33292 7792 33332 7832
rect 38476 7792 38516 7832
rect 39820 7792 39860 7832
rect 48748 7792 48788 7832
rect 17644 7708 17684 7748
rect 17836 7708 17876 7748
rect 19372 7708 19412 7748
rect 19564 7708 19604 7748
rect 20332 7708 20372 7748
rect 22540 7708 22580 7748
rect 22732 7708 22772 7748
rect 23980 7708 24020 7748
rect 27916 7708 27956 7748
rect 29644 7708 29684 7748
rect 29836 7708 29876 7748
rect 33868 7708 33908 7748
rect 37324 7708 37364 7748
rect 38860 7708 38900 7748
rect 39532 7708 39572 7748
rect 12172 7624 12212 7664
rect 48364 7624 48404 7664
rect 1132 7288 1172 7328
rect 4928 7540 4968 7580
rect 5010 7540 5050 7580
rect 5092 7540 5132 7580
rect 5174 7540 5214 7580
rect 5256 7540 5296 7580
rect 17452 7540 17492 7580
rect 19468 7540 19508 7580
rect 20048 7540 20088 7580
rect 20130 7540 20170 7580
rect 20212 7540 20252 7580
rect 20294 7540 20334 7580
rect 20376 7540 20416 7580
rect 22636 7540 22676 7580
rect 23020 7540 23060 7580
rect 24268 7540 24308 7580
rect 24556 7540 24596 7580
rect 32332 7540 32372 7580
rect 35168 7540 35208 7580
rect 35250 7540 35290 7580
rect 35332 7540 35372 7580
rect 35414 7540 35454 7580
rect 35496 7540 35536 7580
rect 36748 7540 36788 7580
rect 39052 7540 39092 7580
rect 50288 7540 50328 7580
rect 50370 7540 50410 7580
rect 50452 7540 50492 7580
rect 50534 7540 50574 7580
rect 50616 7540 50656 7580
rect 5836 7456 5876 7496
rect 25132 7456 25172 7496
rect 30028 7456 30068 7496
rect 34540 7456 34580 7496
rect 37900 7456 37940 7496
rect 41164 7456 41204 7496
rect 15532 7372 15572 7412
rect 20908 7372 20948 7412
rect 26956 7372 26996 7412
rect 27916 7372 27956 7412
rect 30412 7372 30452 7412
rect 33772 7372 33812 7412
rect 34636 7372 34676 7412
rect 38956 7372 38996 7412
rect 40780 7372 40820 7412
rect 52684 7708 52724 7748
rect 16108 7288 16148 7328
rect 23020 7288 23060 7328
rect 33868 7288 33908 7328
rect 52684 7288 52724 7328
rect 19276 7204 19316 7244
rect 23980 7204 24020 7244
rect 30220 7204 30260 7244
rect 39148 7204 39188 7244
rect 10348 7120 10388 7160
rect 11116 7120 11156 7160
rect 11788 7120 11828 7160
rect 12652 7120 12692 7160
rect 13612 7120 13652 7160
rect 14860 7120 14900 7160
rect 15052 7120 15092 7160
rect 16972 7120 17012 7160
rect 17164 7120 17204 7160
rect 27244 7120 27284 7160
rect 28780 7120 28820 7160
rect 37228 7120 37268 7160
rect 37804 7120 37844 7160
rect 38092 7120 38132 7160
rect 39244 7120 39284 7160
rect 51820 7120 51860 7160
rect 9964 7036 10004 7076
rect 26092 7036 26132 7076
rect 26284 7036 26324 7076
rect 37324 7036 37364 7076
rect 38956 7036 38996 7076
rect 39340 7036 39380 7076
rect 40972 7036 41012 7076
rect 652 6952 692 6992
rect 9580 6952 9620 6992
rect 9196 6868 9236 6908
rect 11404 6868 11444 6908
rect 11596 6868 11636 6908
rect 13708 6952 13748 6992
rect 14092 6952 14132 6992
rect 15148 6952 15188 6992
rect 17068 6952 17108 6992
rect 26572 6952 26612 6992
rect 27532 6952 27572 6992
rect 27916 6952 27956 6992
rect 21580 6868 21620 6908
rect 3688 6784 3728 6824
rect 3770 6784 3810 6824
rect 3852 6784 3892 6824
rect 3934 6784 3974 6824
rect 4016 6784 4056 6824
rect 8812 6784 8852 6824
rect 14860 6784 14900 6824
rect 18700 6784 18740 6824
rect 18808 6784 18848 6824
rect 18890 6784 18930 6824
rect 18972 6784 19012 6824
rect 19054 6784 19094 6824
rect 19136 6784 19176 6824
rect 19468 6784 19508 6824
rect 27628 6784 27668 6824
rect 41164 6952 41204 6992
rect 47308 6952 47348 6992
rect 37804 6868 37844 6908
rect 47212 6868 47252 6908
rect 33928 6784 33968 6824
rect 34010 6784 34050 6824
rect 34092 6784 34132 6824
rect 34174 6784 34214 6824
rect 34256 6784 34296 6824
rect 47404 6784 47444 6824
rect 49048 6784 49088 6824
rect 49130 6784 49170 6824
rect 49212 6784 49252 6824
rect 49294 6784 49334 6824
rect 49376 6784 49416 6824
rect 13612 6700 13652 6740
rect 27820 6700 27860 6740
rect 29260 6700 29300 6740
rect 40492 6700 40532 6740
rect 940 6616 980 6656
rect 11788 6616 11828 6656
rect 19180 6616 19220 6656
rect 23308 6616 23348 6656
rect 25516 6616 25556 6656
rect 25708 6616 25748 6656
rect 29068 6616 29108 6656
rect 37324 6616 37364 6656
rect 48940 6616 48980 6656
rect 50092 6616 50132 6656
rect 8428 6532 8468 6572
rect 14092 6532 14132 6572
rect 15244 6532 15284 6572
rect 20524 6532 20564 6572
rect 23404 6532 23444 6572
rect 4108 6448 4148 6488
rect 18700 6448 18740 6488
rect 23212 6448 23252 6488
rect 42604 6532 42644 6572
rect 47308 6532 47348 6572
rect 26380 6448 26420 6488
rect 28204 6448 28244 6488
rect 28396 6448 28436 6488
rect 28876 6448 28916 6488
rect 41548 6448 41588 6488
rect 44044 6448 44084 6488
rect 48940 6448 48980 6488
rect 1420 6280 1460 6320
rect 6604 6280 6644 6320
rect 34732 6364 34772 6404
rect 9100 6196 9140 6236
rect 25708 6196 25748 6236
rect 28972 6196 29012 6236
rect 34732 6196 34772 6236
rect 1132 6112 1172 6152
rect 11596 6112 11636 6152
rect 23212 6112 23252 6152
rect 23788 6112 23828 6152
rect 26380 6112 26420 6152
rect 26572 6112 26612 6152
rect 46828 6280 46868 6320
rect 35116 6196 35156 6236
rect 43084 6196 43124 6236
rect 35020 6112 35060 6152
rect 40588 6112 40628 6152
rect 4928 6028 4968 6068
rect 5010 6028 5050 6068
rect 5092 6028 5132 6068
rect 5174 6028 5214 6068
rect 5256 6028 5296 6068
rect 20048 6028 20088 6068
rect 20130 6028 20170 6068
rect 20212 6028 20252 6068
rect 20294 6028 20334 6068
rect 20376 6028 20416 6068
rect 20524 6028 20564 6068
rect 23116 6028 23156 6068
rect 23308 6028 23348 6068
rect 28396 6028 28436 6068
rect 28588 6028 28628 6068
rect 35168 6028 35208 6068
rect 35250 6028 35290 6068
rect 35332 6028 35372 6068
rect 35414 6028 35454 6068
rect 35496 6028 35536 6068
rect 50288 6028 50328 6068
rect 50370 6028 50410 6068
rect 50452 6028 50492 6068
rect 50534 6028 50574 6068
rect 50616 6028 50656 6068
rect 1036 5944 1076 5984
rect 1228 5944 1268 5984
rect 27244 5944 27284 5984
rect 27532 5944 27572 5984
rect 47500 5944 47540 5984
rect 51916 5944 51956 5984
rect 12652 5860 12692 5900
rect 15244 5860 15284 5900
rect 28780 5860 28820 5900
rect 28972 5860 29012 5900
rect 47308 5860 47348 5900
rect 11116 5776 11156 5816
rect 27436 5776 27476 5816
rect 27916 5776 27956 5816
rect 51820 5776 51860 5816
rect 26380 5692 26420 5732
rect 38092 5692 38132 5732
rect 51532 5692 51572 5732
rect 1612 5608 1652 5648
rect 27628 5608 27668 5648
rect 30028 5608 30068 5648
rect 33292 5608 33332 5648
rect 41740 5608 41780 5648
rect 46540 5608 46580 5648
rect 46732 5608 46772 5648
rect 49996 5608 50036 5648
rect 51820 5608 51860 5648
rect 40300 5524 40340 5564
rect 40492 5524 40532 5564
rect 21964 5440 22004 5480
rect 33100 5440 33140 5480
rect 46444 5440 46484 5480
rect 16588 5356 16628 5396
rect 29836 5356 29876 5396
rect 3688 5272 3728 5312
rect 3770 5272 3810 5312
rect 3852 5272 3892 5312
rect 3934 5272 3974 5312
rect 4016 5272 4056 5312
rect 18808 5272 18848 5312
rect 18890 5272 18930 5312
rect 18972 5272 19012 5312
rect 19054 5272 19094 5312
rect 19136 5272 19176 5312
rect 30124 5272 30164 5312
rect 33292 5272 33332 5312
rect 33928 5272 33968 5312
rect 34010 5272 34050 5312
rect 34092 5272 34132 5312
rect 34174 5272 34214 5312
rect 34256 5272 34296 5312
rect 49048 5272 49088 5312
rect 49130 5272 49170 5312
rect 49212 5272 49252 5312
rect 49294 5272 49334 5312
rect 49376 5272 49416 5312
rect 14092 5188 14132 5228
rect 26380 5188 26420 5228
rect 38092 5188 38132 5228
rect 21772 5104 21812 5144
rect 22060 5104 22100 5144
rect 26764 5104 26804 5144
rect 33196 5104 33236 5144
rect 44236 5104 44276 5144
rect 652 5020 692 5060
rect 27628 5020 27668 5060
rect 41836 5020 41876 5060
rect 21580 4936 21620 4976
rect 32428 4936 32468 4976
rect 32620 4936 32660 4976
rect 25516 4852 25556 4892
rect 19276 4768 19316 4808
rect 26764 4768 26804 4808
rect 40492 4768 40532 4808
rect 51820 4768 51860 4808
rect 23980 4684 24020 4724
rect 30124 4684 30164 4724
rect 46060 4684 46100 4724
rect 22348 4600 22388 4640
rect 4928 4516 4968 4556
rect 5010 4516 5050 4556
rect 5092 4516 5132 4556
rect 5174 4516 5214 4556
rect 5256 4516 5296 4556
rect 20048 4516 20088 4556
rect 20130 4516 20170 4556
rect 20212 4516 20252 4556
rect 20294 4516 20334 4556
rect 20376 4516 20416 4556
rect 21676 4516 21716 4556
rect 32428 4516 32468 4556
rect 35168 4516 35208 4556
rect 35250 4516 35290 4556
rect 35332 4516 35372 4556
rect 35414 4516 35454 4556
rect 35496 4516 35536 4556
rect 50288 4516 50328 4556
rect 50370 4516 50410 4556
rect 50452 4516 50492 4556
rect 50534 4516 50574 4556
rect 50616 4516 50656 4556
rect 23500 4432 23540 4472
rect 24748 4348 24788 4388
rect 32620 4348 32660 4388
rect 19852 4180 19892 4220
rect 31180 4180 31220 4220
rect 17932 4096 17972 4136
rect 23308 4096 23348 4136
rect 24076 4096 24116 4136
rect 24652 4096 24692 4136
rect 19468 4012 19508 4052
rect 7852 3928 7892 3968
rect 21484 3928 21524 3968
rect 21868 3928 21908 3968
rect 3688 3760 3728 3800
rect 3770 3760 3810 3800
rect 3852 3760 3892 3800
rect 3934 3760 3974 3800
rect 4016 3760 4056 3800
rect 18808 3760 18848 3800
rect 18890 3760 18930 3800
rect 18972 3760 19012 3800
rect 19054 3760 19094 3800
rect 19136 3760 19176 3800
rect 31372 4180 31412 4220
rect 51820 4180 51860 4220
rect 25228 4096 25268 4136
rect 25612 4096 25652 4136
rect 25996 4096 26036 4136
rect 26284 4096 26324 4136
rect 47308 4096 47348 4136
rect 22924 3928 22964 3968
rect 23404 3928 23444 3968
rect 24172 3928 24212 3968
rect 24460 3928 24500 3968
rect 25900 3928 25940 3968
rect 33928 3760 33968 3800
rect 34010 3760 34050 3800
rect 34092 3760 34132 3800
rect 34174 3760 34214 3800
rect 34256 3760 34296 3800
rect 49048 3760 49088 3800
rect 49130 3760 49170 3800
rect 49212 3760 49252 3800
rect 49294 3760 49334 3800
rect 49376 3760 49416 3800
rect 18124 3676 18164 3716
rect 23212 3676 23252 3716
rect 25228 3676 25268 3716
rect 22060 3592 22100 3632
rect 23500 3592 23540 3632
rect 24748 3592 24788 3632
rect 25516 3592 25556 3632
rect 28588 3592 28628 3632
rect 21580 3508 21620 3548
rect 24556 3508 24596 3548
rect 25612 3508 25652 3548
rect 21772 3424 21812 3464
rect 21964 3424 22004 3464
rect 24844 3424 24884 3464
rect 28300 3424 28340 3464
rect 47308 3424 47348 3464
rect 51820 3424 51860 3464
rect 7852 3340 7892 3380
rect 22348 3340 22388 3380
rect 24652 3256 24692 3296
rect 23212 3172 23252 3212
rect 25324 3172 25364 3212
rect 18316 3088 18356 3128
rect 23308 3088 23348 3128
rect 4928 3004 4968 3044
rect 5010 3004 5050 3044
rect 5092 3004 5132 3044
rect 5174 3004 5214 3044
rect 5256 3004 5296 3044
rect 20048 3004 20088 3044
rect 20130 3004 20170 3044
rect 20212 3004 20252 3044
rect 20294 3004 20334 3044
rect 20376 3004 20416 3044
rect 35168 3004 35208 3044
rect 35250 3004 35290 3044
rect 35332 3004 35372 3044
rect 35414 3004 35454 3044
rect 35496 3004 35536 3044
rect 50288 3004 50328 3044
rect 50370 3004 50410 3044
rect 50452 3004 50492 3044
rect 50534 3004 50574 3044
rect 50616 3004 50656 3044
rect 24076 2920 24116 2960
rect 25708 2836 25748 2876
rect 24844 2752 24884 2792
rect 25324 2752 25364 2792
rect 24460 2668 24500 2708
rect 24556 2584 24596 2624
rect 1036 2332 1076 2372
rect 3688 2248 3728 2288
rect 3770 2248 3810 2288
rect 3852 2248 3892 2288
rect 3934 2248 3974 2288
rect 4016 2248 4056 2288
rect 18808 2248 18848 2288
rect 18890 2248 18930 2288
rect 18972 2248 19012 2288
rect 19054 2248 19094 2288
rect 19136 2248 19176 2288
rect 21868 2248 21908 2288
rect 50380 2332 50420 2372
rect 33928 2248 33968 2288
rect 34010 2248 34050 2288
rect 34092 2248 34132 2288
rect 34174 2248 34214 2288
rect 34256 2248 34296 2288
rect 49048 2248 49088 2288
rect 49130 2248 49170 2288
rect 49212 2248 49252 2288
rect 49294 2248 49334 2288
rect 49376 2248 49416 2288
rect 24172 2164 24212 2204
rect 25900 2164 25940 2204
rect 23404 2080 23444 2120
rect 23116 1996 23156 2036
rect 45292 1996 45332 2036
rect 19468 1912 19508 1952
rect 21484 1912 21524 1952
rect 50380 1912 50420 1952
rect 43084 1828 43124 1868
rect 43276 1828 43316 1868
rect 50572 1828 50612 1868
rect 50764 1828 50804 1868
rect 52300 1828 52340 1868
rect 45292 1744 45332 1784
rect 52972 1744 53012 1784
rect 19852 1576 19892 1616
rect 4928 1492 4968 1532
rect 5010 1492 5050 1532
rect 5092 1492 5132 1532
rect 5174 1492 5214 1532
rect 5256 1492 5296 1532
rect 20048 1492 20088 1532
rect 20130 1492 20170 1532
rect 20212 1492 20252 1532
rect 20294 1492 20334 1532
rect 20376 1492 20416 1532
rect 35168 1492 35208 1532
rect 35250 1492 35290 1532
rect 35332 1492 35372 1532
rect 35414 1492 35454 1532
rect 35496 1492 35536 1532
rect 50288 1492 50328 1532
rect 50370 1492 50410 1532
rect 50452 1492 50492 1532
rect 50534 1492 50574 1532
rect 50616 1492 50656 1532
rect 53164 1408 53204 1448
rect 18316 1240 18356 1280
rect 53164 1240 53204 1280
rect 18124 904 18164 944
rect 52972 904 53012 944
rect 17932 568 17972 608
rect 52300 568 52340 608
<< metal3 >>
rect 2744 11764 2824 11844
rect 3128 11764 3208 11844
rect 3512 11764 3592 11844
rect 3896 11764 3976 11844
rect 4280 11764 4360 11844
rect 4664 11764 4744 11844
rect 5048 11764 5128 11844
rect 5432 11764 5512 11844
rect 5816 11764 5896 11844
rect 6200 11764 6280 11844
rect 6584 11764 6664 11844
rect 6968 11764 7048 11844
rect 7352 11764 7432 11844
rect 7736 11764 7816 11844
rect 8120 11764 8200 11844
rect 8504 11764 8584 11844
rect 8888 11764 8968 11844
rect 9272 11764 9352 11844
rect 9656 11764 9736 11844
rect 10040 11764 10120 11844
rect 10424 11764 10504 11844
rect 10808 11764 10888 11844
rect 11192 11764 11272 11844
rect 11576 11764 11656 11844
rect 11960 11764 12040 11844
rect 12344 11764 12424 11844
rect 12728 11764 12808 11844
rect 13112 11764 13192 11844
rect 13496 11764 13576 11844
rect 13880 11764 13960 11844
rect 14264 11764 14344 11844
rect 14648 11764 14728 11844
rect 15032 11764 15112 11844
rect 15416 11764 15496 11844
rect 15800 11764 15880 11844
rect 16184 11764 16264 11844
rect 16568 11764 16648 11844
rect 16952 11764 17032 11844
rect 17164 11780 17204 11789
rect 748 11024 788 11033
rect 556 10688 596 10697
rect 268 9344 308 9353
rect 268 8000 308 9304
rect 556 8840 596 10648
rect 556 8791 596 8800
rect 748 8672 788 10984
rect 1228 10352 1268 10361
rect 1228 8924 1268 10312
rect 1420 10016 1460 10025
rect 1420 9881 1460 9976
rect 2764 9680 2804 11764
rect 2764 9631 2804 9640
rect 3148 9680 3188 11764
rect 3148 9631 3188 9640
rect 3532 9680 3572 11764
rect 3916 10352 3956 11764
rect 3916 10312 4148 10352
rect 3688 9848 4056 9857
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 3688 9799 4056 9808
rect 3532 9631 3572 9640
rect 4108 9680 4148 10312
rect 4108 9631 4148 9640
rect 4300 9680 4340 11764
rect 4300 9631 4340 9640
rect 4684 9680 4724 11764
rect 4684 9631 4724 9640
rect 5068 9680 5108 11764
rect 5068 9631 5108 9640
rect 5452 9680 5492 11764
rect 5452 9631 5492 9640
rect 5836 9680 5876 11764
rect 5836 9631 5876 9640
rect 6220 9680 6260 11764
rect 6220 9631 6260 9640
rect 6604 9680 6644 11764
rect 6604 9631 6644 9640
rect 6988 9680 7028 11764
rect 6988 9631 7028 9640
rect 7372 9680 7412 11764
rect 7372 9631 7412 9640
rect 7756 9680 7796 11764
rect 7756 9631 7796 9640
rect 8140 9680 8180 11764
rect 8140 9631 8180 9640
rect 8524 9680 8564 11764
rect 8524 9631 8564 9640
rect 8620 10016 8660 10025
rect 7180 9596 7220 9605
rect 4108 9512 4148 9521
rect 1228 8875 1268 8884
rect 1420 9008 1460 9017
rect 748 8623 788 8632
rect 1420 8672 1460 8968
rect 1420 8623 1460 8632
rect 3688 8336 4056 8345
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 3688 8287 4056 8296
rect 4108 8168 4148 9472
rect 4588 9512 4628 9521
rect 4108 8119 4148 8128
rect 4300 9428 4340 9437
rect 4300 8168 4340 9388
rect 4588 9260 4628 9472
rect 4588 9211 4628 9220
rect 5356 9512 5396 9521
rect 4928 9092 5296 9101
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 4928 9043 5296 9052
rect 5356 8840 5396 9472
rect 6892 9512 6932 9521
rect 5644 9428 5684 9437
rect 5644 8924 5684 9388
rect 6028 9428 6068 9437
rect 6028 9092 6068 9388
rect 6028 9043 6068 9052
rect 5644 8875 5684 8884
rect 5356 8791 5396 8800
rect 4300 8119 4340 8128
rect 6124 8588 6164 8597
rect 268 7951 308 7960
rect 1228 8000 1268 8009
rect 1132 7328 1172 7337
rect 652 6992 692 7001
rect 652 5060 692 6952
rect 652 5011 692 5020
rect 940 6656 980 6665
rect 940 4136 980 6616
rect 1132 6152 1172 7288
rect 1132 6103 1172 6112
rect 940 4087 980 4096
rect 1036 5984 1076 5993
rect 1036 2372 1076 5944
rect 1228 5984 1268 7960
rect 5836 8000 5876 8009
rect 4928 7580 5296 7589
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 4928 7531 5296 7540
rect 5836 7496 5876 7960
rect 6124 8000 6164 8548
rect 6892 8168 6932 9472
rect 6892 8119 6932 8128
rect 7084 9512 7124 9521
rect 7084 8084 7124 9472
rect 7084 8035 7124 8044
rect 6124 7951 6164 7960
rect 7180 7832 7220 9556
rect 8044 9512 8084 9521
rect 7756 9428 7796 9437
rect 7756 8168 7796 9388
rect 8044 9176 8084 9472
rect 8044 9127 8084 9136
rect 8428 9512 8468 9521
rect 7756 8119 7796 8128
rect 7180 7783 7220 7792
rect 5836 7447 5876 7456
rect 3688 6824 4056 6833
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 3688 6775 4056 6784
rect 8428 6572 8468 9472
rect 8620 9344 8660 9976
rect 8908 9680 8948 11764
rect 8908 9631 8948 9640
rect 9292 9680 9332 11764
rect 9292 9631 9332 9640
rect 9676 9680 9716 11764
rect 9676 9631 9716 9640
rect 10060 9680 10100 11764
rect 10060 9631 10100 9640
rect 10444 9680 10484 11764
rect 10444 9631 10484 9640
rect 10636 9764 10676 9773
rect 8620 9295 8660 9304
rect 8812 9512 8852 9521
rect 8812 6824 8852 9472
rect 9196 9512 9236 9521
rect 9196 6908 9236 9472
rect 9580 9512 9620 9521
rect 9580 6992 9620 9472
rect 9964 9512 10004 9521
rect 9964 7076 10004 9472
rect 10348 9512 10388 9521
rect 10156 9344 10196 9353
rect 10060 8420 10100 8429
rect 10060 8285 10100 8380
rect 10156 8168 10196 9304
rect 10156 8119 10196 8128
rect 10252 8336 10292 8345
rect 10252 8084 10292 8296
rect 10252 8035 10292 8044
rect 10060 7916 10100 7925
rect 10060 7781 10100 7876
rect 10348 7160 10388 9472
rect 10636 8000 10676 9724
rect 10828 9680 10868 11764
rect 10828 9631 10868 9640
rect 11212 9680 11252 11764
rect 11212 9631 11252 9640
rect 11596 9680 11636 11764
rect 11596 9631 11636 9640
rect 11980 9680 12020 11764
rect 11980 9631 12020 9640
rect 12364 9680 12404 11764
rect 12364 9631 12404 9640
rect 12748 9680 12788 11764
rect 12748 9631 12788 9640
rect 13132 9680 13172 11764
rect 13228 9932 13268 9941
rect 13228 9797 13268 9892
rect 13132 9631 13172 9640
rect 13516 9680 13556 11764
rect 13516 9631 13556 9640
rect 13804 9932 13844 9941
rect 13324 9596 13364 9605
rect 11116 9512 11156 9521
rect 11116 9377 11156 9472
rect 12652 9512 12692 9521
rect 11500 9092 11540 9101
rect 11500 8084 11540 9052
rect 11596 9008 11636 9017
rect 11788 9008 11828 9017
rect 11636 8968 11788 9008
rect 11596 8959 11636 8968
rect 11788 8959 11828 8968
rect 12652 8672 12692 9472
rect 13228 9512 13268 9521
rect 12940 9176 12980 9185
rect 12980 9136 13076 9176
rect 12940 9108 12980 9136
rect 12652 8623 12692 8632
rect 12844 8420 12884 8429
rect 12844 8168 12884 8380
rect 12844 8119 12884 8128
rect 13036 8168 13076 9136
rect 13228 8756 13268 9472
rect 13324 8840 13364 9556
rect 13324 8791 13364 8800
rect 13708 8924 13748 8933
rect 13804 8924 13844 9892
rect 13900 9680 13940 11764
rect 13900 9631 13940 9640
rect 14188 9932 14228 9941
rect 14188 9512 14228 9892
rect 14284 9680 14324 11764
rect 14284 9631 14324 9640
rect 14668 9680 14708 11764
rect 14668 9631 14708 9640
rect 15052 9680 15092 11764
rect 15052 9631 15092 9640
rect 15436 9680 15476 11764
rect 15436 9631 15476 9640
rect 15820 9680 15860 11764
rect 15820 9631 15860 9640
rect 16012 10016 16052 10025
rect 14188 9463 14228 9472
rect 14380 9512 14420 9521
rect 13900 8924 13940 8933
rect 13804 8884 13900 8924
rect 13228 8707 13268 8716
rect 13036 8119 13076 8128
rect 11500 8035 11540 8044
rect 12172 8084 12212 8093
rect 10636 7951 10676 7960
rect 12172 7664 12212 8044
rect 12172 7615 12212 7624
rect 10348 7111 10388 7120
rect 11116 7160 11156 7169
rect 9964 7027 10004 7036
rect 9580 6943 9620 6952
rect 9196 6859 9236 6868
rect 8812 6775 8852 6784
rect 8428 6523 8468 6532
rect 4108 6488 4148 6497
rect 1228 5935 1268 5944
rect 1420 6320 1460 6329
rect 1420 3464 1460 6280
rect 1420 3415 1460 3424
rect 1612 5648 1652 5657
rect 1036 2323 1076 2332
rect 1612 80 1652 5608
rect 3688 5312 4056 5321
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 3688 5263 4056 5272
rect 3688 3800 4056 3809
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 3688 3751 4056 3760
rect 3688 2288 4056 2297
rect 3728 2248 3770 2288
rect 3810 2248 3852 2288
rect 3892 2248 3934 2288
rect 3974 2248 4016 2288
rect 3688 2239 4056 2248
rect 4108 80 4148 6448
rect 6604 6320 6644 6329
rect 4928 6068 5296 6077
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 4928 6019 5296 6028
rect 4928 4556 5296 4565
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 4928 4507 5296 4516
rect 4928 3044 5296 3053
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 4928 2995 5296 3004
rect 4928 1532 5296 1541
rect 4968 1492 5010 1532
rect 5050 1492 5092 1532
rect 5132 1492 5174 1532
rect 5214 1492 5256 1532
rect 4928 1483 5296 1492
rect 6604 80 6644 6280
rect 9100 6236 9140 6245
rect 7852 3968 7892 3977
rect 7852 3380 7892 3928
rect 7852 3331 7892 3340
rect 9100 80 9140 6196
rect 11116 5816 11156 7120
rect 11788 7160 11828 7169
rect 11404 6908 11444 6917
rect 11596 6908 11636 6917
rect 11444 6868 11596 6908
rect 11404 6859 11444 6868
rect 11596 6859 11636 6868
rect 11788 6656 11828 7120
rect 11788 6607 11828 6616
rect 12652 7160 12692 7169
rect 11116 5767 11156 5776
rect 11596 6152 11636 6161
rect 11596 80 11636 6112
rect 12652 5900 12692 7120
rect 13612 7160 13652 7169
rect 13612 6740 13652 7120
rect 13708 6992 13748 8884
rect 13900 8875 13940 8884
rect 14380 8420 14420 9472
rect 15148 9512 15188 9521
rect 14380 8371 14420 8380
rect 15052 9092 15092 9101
rect 14860 7160 14900 7169
rect 13708 6943 13748 6952
rect 14092 6992 14132 7001
rect 13612 6691 13652 6700
rect 14092 6572 14132 6952
rect 14860 6824 14900 7120
rect 15052 7160 15092 9052
rect 15052 7111 15092 7120
rect 15148 6992 15188 9472
rect 15916 9512 15956 9521
rect 15628 9260 15668 9269
rect 15340 8504 15380 8513
rect 15340 8000 15380 8464
rect 15628 8168 15668 9220
rect 15820 8588 15860 8597
rect 15820 8504 15860 8548
rect 15820 8453 15860 8464
rect 15916 8420 15956 9472
rect 15916 8371 15956 8380
rect 15628 8119 15668 8128
rect 16012 8168 16052 9976
rect 16204 9680 16244 11764
rect 16300 10016 16340 10027
rect 16300 9932 16340 9976
rect 16300 9883 16340 9892
rect 16204 9631 16244 9640
rect 16588 9680 16628 11764
rect 16588 9631 16628 9640
rect 16684 11192 16724 11201
rect 16396 9428 16436 9437
rect 16300 9344 16340 9353
rect 16300 8420 16340 9304
rect 16300 8371 16340 8380
rect 16012 8119 16052 8128
rect 16396 8168 16436 9388
rect 16396 8119 16436 8128
rect 15340 7951 15380 7960
rect 16108 8000 16148 8009
rect 15436 7916 15476 7925
rect 15436 7412 15476 7876
rect 15532 7412 15572 7421
rect 15436 7372 15532 7412
rect 15532 7363 15572 7372
rect 16108 7328 16148 7960
rect 16684 7916 16724 11152
rect 16972 9680 17012 11764
rect 16972 9631 17012 9640
rect 17336 11764 17416 11844
rect 17720 11764 17800 11844
rect 18104 11764 18184 11844
rect 18488 11764 18568 11844
rect 18872 11764 18952 11844
rect 19256 11764 19336 11844
rect 19640 11764 19720 11844
rect 20024 11764 20104 11844
rect 20408 11764 20488 11844
rect 20792 11764 20872 11844
rect 21176 11764 21256 11844
rect 21560 11764 21640 11844
rect 21944 11764 22024 11844
rect 22328 11764 22408 11844
rect 22712 11764 22792 11844
rect 23096 11764 23176 11844
rect 23480 11764 23560 11844
rect 23864 11764 23944 11844
rect 24248 11764 24328 11844
rect 24632 11764 24712 11844
rect 25016 11764 25096 11844
rect 25400 11764 25480 11844
rect 25784 11764 25864 11844
rect 26168 11764 26248 11844
rect 26552 11764 26632 11844
rect 26936 11764 27016 11844
rect 27320 11764 27400 11844
rect 27704 11764 27784 11844
rect 28088 11764 28168 11844
rect 28472 11764 28552 11844
rect 28856 11764 28936 11844
rect 29240 11764 29320 11844
rect 29624 11764 29704 11844
rect 30008 11764 30088 11844
rect 30392 11764 30472 11844
rect 30776 11764 30856 11844
rect 31160 11764 31240 11844
rect 31544 11764 31624 11844
rect 31928 11780 32008 11844
rect 31928 11764 31948 11780
rect 17068 8504 17108 8513
rect 16780 8420 16820 8429
rect 16780 8168 16820 8380
rect 16780 8119 16820 8128
rect 17068 8084 17108 8464
rect 17068 8035 17108 8044
rect 16684 7867 16724 7876
rect 16108 7279 16148 7288
rect 16972 7160 17012 7169
rect 16972 6992 17012 7120
rect 17164 7160 17204 11740
rect 17260 11696 17300 11705
rect 17260 8168 17300 11656
rect 17356 9680 17396 11764
rect 17356 9631 17396 9640
rect 17740 9680 17780 11764
rect 17740 9631 17780 9640
rect 18028 10268 18068 10277
rect 17932 9596 17972 9605
rect 17836 9428 17876 9437
rect 17836 9293 17876 9388
rect 17548 9092 17588 9101
rect 17452 9008 17492 9017
rect 17452 8756 17492 8968
rect 17452 8707 17492 8716
rect 17260 8119 17300 8128
rect 17548 8168 17588 9052
rect 17836 8840 17876 8849
rect 17836 8756 17876 8800
rect 17836 8705 17876 8716
rect 17548 8119 17588 8128
rect 17932 8168 17972 9556
rect 18028 8588 18068 10228
rect 18124 9680 18164 11764
rect 18412 9848 18452 9857
rect 18124 9631 18164 9640
rect 18316 9764 18356 9773
rect 18028 8539 18068 8548
rect 17932 8119 17972 8128
rect 18220 8504 18260 8513
rect 17452 8000 17492 8009
rect 17452 7580 17492 7960
rect 17836 8000 17876 8009
rect 17644 7748 17684 7757
rect 17644 7613 17684 7708
rect 17836 7748 17876 7960
rect 18220 8000 18260 8464
rect 18316 8168 18356 9724
rect 18316 8119 18356 8128
rect 18412 8084 18452 9808
rect 18508 9680 18548 11764
rect 18892 10016 18932 11764
rect 18508 9631 18548 9640
rect 18700 9976 18932 10016
rect 18700 9596 18740 9976
rect 18808 9848 19176 9857
rect 18848 9808 18890 9848
rect 18930 9808 18972 9848
rect 19012 9808 19054 9848
rect 19094 9808 19136 9848
rect 18808 9799 19176 9808
rect 19276 9680 19316 11764
rect 19276 9631 19316 9640
rect 19372 11612 19412 11621
rect 18700 9547 18740 9556
rect 18604 9512 18644 9521
rect 18604 9008 18644 9472
rect 19084 9428 19124 9437
rect 18988 9344 19028 9353
rect 18604 8959 18644 8968
rect 18700 9176 18740 9185
rect 18412 8035 18452 8044
rect 18604 8588 18644 8597
rect 18220 7951 18260 7960
rect 18604 8000 18644 8548
rect 18700 8168 18740 9136
rect 18988 8756 19028 9304
rect 19084 9176 19124 9388
rect 19276 9428 19316 9437
rect 19276 9293 19316 9388
rect 19084 9127 19124 9136
rect 18988 8707 19028 8716
rect 18808 8336 19176 8345
rect 18848 8296 18890 8336
rect 18930 8296 18972 8336
rect 19012 8296 19054 8336
rect 19094 8296 19136 8336
rect 18808 8287 19176 8296
rect 18700 8119 18740 8128
rect 18604 7951 18644 7960
rect 19276 8000 19316 8009
rect 17836 7699 17876 7708
rect 17452 7531 17492 7540
rect 19276 7244 19316 7960
rect 19372 7748 19412 11572
rect 19564 11528 19604 11537
rect 19468 10016 19508 10025
rect 19468 9848 19508 9976
rect 19468 9799 19508 9808
rect 19564 9680 19604 11488
rect 19372 7699 19412 7708
rect 19468 9640 19604 9680
rect 19660 9680 19700 11764
rect 19468 7580 19508 9640
rect 19660 9631 19700 9640
rect 19852 11444 19892 11453
rect 19660 9176 19700 9185
rect 19564 8252 19604 8261
rect 19564 7748 19604 8212
rect 19564 7699 19604 7708
rect 19468 7531 19508 7540
rect 19660 7496 19700 9136
rect 19756 9008 19796 9017
rect 19756 7748 19796 8968
rect 19852 8504 19892 11404
rect 20044 9680 20084 11764
rect 20044 9631 20084 9640
rect 20140 9764 20180 9773
rect 20140 9629 20180 9724
rect 20332 9764 20372 9773
rect 19948 9512 19988 9521
rect 19948 9176 19988 9472
rect 20140 9260 20180 9269
rect 20332 9260 20372 9724
rect 20428 9680 20468 11764
rect 20428 9631 20468 9640
rect 20812 9680 20852 11764
rect 20812 9631 20852 9640
rect 20908 9848 20948 9857
rect 20620 9596 20660 9605
rect 20180 9220 20372 9260
rect 20524 9512 20564 9521
rect 20140 9211 20180 9220
rect 19948 9127 19988 9136
rect 20524 9176 20564 9472
rect 20524 9127 20564 9136
rect 20048 9092 20416 9101
rect 20088 9052 20130 9092
rect 20170 9052 20212 9092
rect 20252 9052 20294 9092
rect 20334 9052 20376 9092
rect 20048 9043 20416 9052
rect 20620 9092 20660 9556
rect 20620 9043 20660 9052
rect 20236 8924 20276 8933
rect 20716 8924 20756 8933
rect 20276 8884 20716 8924
rect 20236 8875 20276 8884
rect 20716 8875 20756 8884
rect 19852 8455 19892 8464
rect 20044 8756 20084 8765
rect 20044 8504 20084 8716
rect 20140 8756 20180 8765
rect 20140 8672 20180 8716
rect 20716 8672 20756 8681
rect 20140 8632 20276 8672
rect 20044 8455 20084 8464
rect 20140 8336 20180 8431
rect 20140 8287 20180 8296
rect 20236 8084 20276 8632
rect 20332 8504 20372 8513
rect 20372 8464 20468 8504
rect 20332 8455 20372 8464
rect 20428 8420 20468 8464
rect 20428 8371 20468 8380
rect 20332 8336 20372 8345
rect 20332 8201 20372 8296
rect 20716 8168 20756 8632
rect 20716 8119 20756 8128
rect 20236 8035 20276 8044
rect 20332 7748 20372 7757
rect 19756 7708 20332 7748
rect 20332 7699 20372 7708
rect 20048 7580 20416 7589
rect 20088 7540 20130 7580
rect 20170 7540 20212 7580
rect 20252 7540 20294 7580
rect 20334 7540 20376 7580
rect 20048 7531 20416 7540
rect 19660 7447 19700 7456
rect 20908 7412 20948 9808
rect 21196 9680 21236 11764
rect 21196 9631 21236 9640
rect 21580 9680 21620 11764
rect 21580 9631 21620 9640
rect 21964 9680 22004 11764
rect 21964 9631 22004 9640
rect 22348 9680 22388 11764
rect 22732 9932 22772 11764
rect 23116 10352 23156 11764
rect 23116 10312 23252 10352
rect 23116 10184 23156 10193
rect 22540 9892 22772 9932
rect 22828 9932 22868 9941
rect 22348 9631 22388 9640
rect 22444 9848 22484 9857
rect 21772 9596 21812 9605
rect 21292 9512 21332 9521
rect 21676 9512 21716 9521
rect 21332 9472 21620 9512
rect 21292 9463 21332 9472
rect 21004 9428 21044 9437
rect 21004 8000 21044 9388
rect 21484 9008 21524 9017
rect 21484 8504 21524 8968
rect 21484 8455 21524 8464
rect 21004 7951 21044 7960
rect 21196 8000 21236 8009
rect 21196 7748 21236 7960
rect 21196 7699 21236 7708
rect 20908 7363 20948 7372
rect 19276 7195 19316 7204
rect 17164 7111 17204 7120
rect 17068 6992 17108 7001
rect 16972 6952 17068 6992
rect 15148 6943 15188 6952
rect 17068 6943 17108 6952
rect 21580 6908 21620 9472
rect 21676 7832 21716 9472
rect 21676 7783 21716 7792
rect 21772 7748 21812 9556
rect 22252 9596 22292 9605
rect 22252 9428 22292 9556
rect 22252 9379 22292 9388
rect 22348 9512 22388 9521
rect 22156 9344 22196 9353
rect 22156 9260 22196 9304
rect 22348 9344 22388 9472
rect 22348 9295 22388 9304
rect 22156 9209 22196 9220
rect 22156 8924 22196 8933
rect 21868 8672 21908 8681
rect 22156 8672 22196 8884
rect 21908 8632 22196 8672
rect 21868 8623 21908 8632
rect 22444 8504 22484 9808
rect 22444 8455 22484 8464
rect 22540 8000 22580 9892
rect 22636 9680 22676 9689
rect 22636 8924 22676 9640
rect 22636 8875 22676 8884
rect 22732 9176 22772 9185
rect 22732 8672 22772 9136
rect 22828 8924 22868 9892
rect 23020 9512 23060 9521
rect 22828 8875 22868 8884
rect 22924 9260 22964 9269
rect 22732 8623 22772 8632
rect 22924 8504 22964 9220
rect 23020 9092 23060 9472
rect 23020 9043 23060 9052
rect 23116 9008 23156 10144
rect 23116 8959 23156 8968
rect 22924 8455 22964 8464
rect 22540 7951 22580 7960
rect 22732 8000 22772 8009
rect 21772 7699 21812 7708
rect 22540 7748 22580 7757
rect 22540 7328 22580 7708
rect 22732 7748 22772 7960
rect 23212 7832 23252 10312
rect 23308 10100 23348 10109
rect 23308 8672 23348 10060
rect 23308 8623 23348 8632
rect 23500 8420 23540 11764
rect 23884 9848 23924 11764
rect 23884 9799 23924 9808
rect 23884 9680 23924 9689
rect 23884 8672 23924 9640
rect 23884 8623 23924 8632
rect 24172 9092 24212 9101
rect 23500 8371 23540 8380
rect 24172 8420 24212 9052
rect 24172 8371 24212 8380
rect 23212 7783 23252 7792
rect 22732 7699 22772 7708
rect 23980 7748 24020 7757
rect 22636 7580 22676 7589
rect 22636 7496 22676 7540
rect 23020 7580 23060 7589
rect 23020 7496 23060 7540
rect 22636 7456 23060 7496
rect 23020 7328 23060 7337
rect 22540 7288 23020 7328
rect 23020 7279 23060 7288
rect 23980 7244 24020 7708
rect 24268 7580 24308 11764
rect 24652 10268 24692 11764
rect 25036 11192 25076 11764
rect 25036 11143 25076 11152
rect 24652 10219 24692 10228
rect 24940 9596 24980 9605
rect 24940 9428 24980 9556
rect 25420 9512 25460 11764
rect 25420 9463 25460 9472
rect 25516 9932 25556 9941
rect 24940 9379 24980 9388
rect 24844 9344 24884 9353
rect 24268 7531 24308 7540
rect 24556 9260 24596 9269
rect 24556 7580 24596 9220
rect 24844 8756 24884 9304
rect 24844 8707 24884 8716
rect 25036 9344 25076 9353
rect 25036 8756 25076 9304
rect 25036 8707 25076 8716
rect 25228 9344 25268 9353
rect 25228 8588 25268 9304
rect 25228 8539 25268 8548
rect 25324 9176 25364 9185
rect 25132 8252 25172 8261
rect 25036 8168 25076 8177
rect 25036 7916 25076 8128
rect 25036 7867 25076 7876
rect 24556 7531 24596 7540
rect 25132 7496 25172 8212
rect 25324 8252 25364 9136
rect 25324 8203 25364 8212
rect 25132 7447 25172 7456
rect 23980 7195 24020 7204
rect 21580 6859 21620 6868
rect 14860 6775 14900 6784
rect 18700 6824 18740 6833
rect 14092 6523 14132 6532
rect 15244 6572 15284 6581
rect 12652 5851 12692 5860
rect 15244 5900 15284 6532
rect 18700 6488 18740 6784
rect 18808 6824 19176 6833
rect 18848 6784 18890 6824
rect 18930 6784 18972 6824
rect 19012 6784 19054 6824
rect 19094 6784 19136 6824
rect 18808 6775 19176 6784
rect 19468 6824 19508 6833
rect 19180 6656 19220 6665
rect 19468 6656 19508 6784
rect 19220 6616 19508 6656
rect 23308 6656 23348 6665
rect 19180 6607 19220 6616
rect 18700 6439 18740 6448
rect 20524 6572 20564 6581
rect 20048 6068 20416 6077
rect 20088 6028 20130 6068
rect 20170 6028 20212 6068
rect 20252 6028 20294 6068
rect 20334 6028 20376 6068
rect 20048 6019 20416 6028
rect 20524 6068 20564 6532
rect 23212 6488 23252 6497
rect 23212 6152 23252 6448
rect 23212 6103 23252 6112
rect 20524 6019 20564 6028
rect 23116 6068 23156 6077
rect 23116 5933 23156 6028
rect 23308 6068 23348 6616
rect 25516 6656 25556 9892
rect 25804 8504 25844 11764
rect 25804 8455 25844 8464
rect 26092 7076 26132 7085
rect 26188 7076 26228 11764
rect 26132 7036 26228 7076
rect 26284 7076 26324 7085
rect 26092 7027 26132 7036
rect 25516 6607 25556 6616
rect 25708 6656 25748 6667
rect 23404 6572 23444 6581
rect 23404 6437 23444 6532
rect 25708 6572 25748 6616
rect 25708 6523 25748 6532
rect 25708 6236 25748 6245
rect 23308 6019 23348 6028
rect 23788 6152 23828 6163
rect 23788 6068 23828 6112
rect 23788 6019 23828 6028
rect 15244 5851 15284 5860
rect 21964 5480 22004 5489
rect 16588 5396 16628 5405
rect 14092 5228 14132 5237
rect 14092 80 14132 5188
rect 16588 80 16628 5356
rect 18808 5312 19176 5321
rect 18848 5272 18890 5312
rect 18930 5272 18972 5312
rect 19012 5272 19054 5312
rect 19094 5272 19136 5312
rect 18808 5263 19176 5272
rect 21772 5144 21812 5153
rect 21580 4976 21620 4985
rect 19276 4808 19316 4817
rect 17932 4136 17972 4145
rect 17932 608 17972 4096
rect 18808 3800 19176 3809
rect 18848 3760 18890 3800
rect 18930 3760 18972 3800
rect 19012 3760 19054 3800
rect 19094 3760 19136 3800
rect 18808 3751 19176 3760
rect 18124 3716 18164 3725
rect 18124 944 18164 3676
rect 18316 3128 18356 3137
rect 18316 1280 18356 3088
rect 18808 2288 19176 2297
rect 18848 2248 18890 2288
rect 18930 2248 18972 2288
rect 19012 2248 19054 2288
rect 19094 2248 19136 2288
rect 18808 2239 19176 2248
rect 18316 1231 18356 1240
rect 18124 895 18164 904
rect 17932 559 17972 568
rect 19276 188 19316 4768
rect 20048 4556 20416 4565
rect 20088 4516 20130 4556
rect 20170 4516 20212 4556
rect 20252 4516 20294 4556
rect 20334 4516 20376 4556
rect 20048 4507 20416 4516
rect 19852 4220 19892 4229
rect 19468 4052 19508 4061
rect 19468 1952 19508 4012
rect 19468 1903 19508 1912
rect 19852 1616 19892 4180
rect 21484 3968 21524 3977
rect 20048 3044 20416 3053
rect 20088 3004 20130 3044
rect 20170 3004 20212 3044
rect 20252 3004 20294 3044
rect 20334 3004 20376 3044
rect 20048 2995 20416 3004
rect 21484 1952 21524 3928
rect 21580 3548 21620 4936
rect 21580 3499 21620 3508
rect 21676 4556 21716 4565
rect 21484 1903 21524 1912
rect 21676 1868 21716 4516
rect 21772 3464 21812 5104
rect 21772 3415 21812 3424
rect 21868 3968 21908 3977
rect 21868 2288 21908 3928
rect 21964 3464 22004 5440
rect 22060 5144 22100 5153
rect 22060 3632 22100 5104
rect 25516 4892 25556 4901
rect 23980 4724 24020 4733
rect 22060 3583 22100 3592
rect 22348 4640 22388 4649
rect 21964 3415 22004 3424
rect 22348 3380 22388 4600
rect 23500 4472 23540 4481
rect 23308 4136 23348 4145
rect 22348 3331 22388 3340
rect 22924 3968 22964 3977
rect 22924 2900 22964 3928
rect 23212 3716 23252 3725
rect 23212 3212 23252 3676
rect 23212 3163 23252 3172
rect 23308 3128 23348 4096
rect 23308 3079 23348 3088
rect 23404 3968 23444 3977
rect 22924 2860 23156 2900
rect 21868 2239 21908 2248
rect 23116 2036 23156 2860
rect 23404 2120 23444 3928
rect 23500 3632 23540 4432
rect 23500 3583 23540 3592
rect 23404 2071 23444 2080
rect 23116 1987 23156 1996
rect 19852 1567 19892 1576
rect 21580 1828 21716 1868
rect 20048 1532 20416 1541
rect 20088 1492 20130 1532
rect 20170 1492 20212 1532
rect 20252 1492 20294 1532
rect 20334 1492 20376 1532
rect 20048 1483 20416 1492
rect 19084 148 19316 188
rect 19084 80 19124 148
rect 21580 80 21620 1828
rect 23980 1448 24020 4684
rect 24748 4388 24788 4397
rect 24076 4136 24116 4145
rect 24076 2960 24116 4096
rect 24652 4136 24692 4145
rect 24076 2911 24116 2920
rect 24172 3968 24212 3977
rect 24172 2204 24212 3928
rect 24460 3968 24500 3977
rect 24460 2708 24500 3928
rect 24460 2659 24500 2668
rect 24556 3548 24596 3557
rect 24556 2624 24596 3508
rect 24652 3296 24692 4096
rect 24748 3632 24788 4348
rect 25228 4136 25268 4145
rect 25228 3716 25268 4096
rect 25228 3667 25268 3676
rect 24748 3583 24788 3592
rect 25516 3632 25556 4852
rect 25516 3583 25556 3592
rect 25612 4136 25652 4145
rect 25612 3548 25652 4096
rect 25612 3499 25652 3508
rect 24652 3247 24692 3256
rect 24844 3464 24884 3473
rect 24844 2792 24884 3424
rect 24844 2743 24884 2752
rect 25324 3212 25364 3221
rect 25324 2792 25364 3172
rect 25708 2876 25748 6196
rect 25996 4136 26036 4145
rect 25996 4001 26036 4096
rect 26284 4136 26324 7036
rect 26572 6992 26612 11764
rect 26764 8672 26804 8681
rect 26764 8588 26804 8632
rect 26764 8537 26804 8548
rect 26956 7412 26996 11764
rect 27340 9512 27380 11764
rect 27340 9472 27476 9512
rect 27148 8924 27188 8933
rect 27148 8672 27188 8884
rect 27148 8623 27188 8632
rect 26956 7363 26996 7372
rect 26572 6943 26612 6952
rect 27244 7160 27284 7169
rect 26380 6488 26420 6497
rect 26380 6152 26420 6448
rect 26380 6103 26420 6112
rect 26572 6152 26612 6161
rect 26380 5732 26420 5741
rect 26380 5228 26420 5692
rect 26380 5179 26420 5188
rect 26284 4087 26324 4096
rect 25708 2827 25748 2836
rect 25900 3968 25940 3977
rect 25324 2743 25364 2752
rect 24556 2575 24596 2584
rect 24172 2155 24212 2164
rect 25900 2204 25940 3928
rect 25900 2155 25940 2164
rect 23980 1408 24116 1448
rect 24076 80 24116 1408
rect 26572 80 26612 6112
rect 27244 5984 27284 7120
rect 27244 5935 27284 5944
rect 27436 5816 27476 9472
rect 27724 9344 27764 11764
rect 28108 11696 28148 11764
rect 27628 9304 27764 9344
rect 27820 11656 28148 11696
rect 27532 8840 27572 8849
rect 27532 8672 27572 8800
rect 27532 8623 27572 8632
rect 27532 6992 27572 7001
rect 27532 5984 27572 6952
rect 27628 6824 27668 9304
rect 27724 9176 27764 9185
rect 27724 8672 27764 9136
rect 27724 8623 27764 8632
rect 27628 6775 27668 6784
rect 27820 6740 27860 11656
rect 28012 10016 28052 10025
rect 28012 8672 28052 9976
rect 28492 8924 28532 11764
rect 28012 8623 28052 8632
rect 28300 8884 28532 8924
rect 28588 10016 28628 10025
rect 28108 8420 28148 8429
rect 28108 7832 28148 8380
rect 28108 7783 28148 7792
rect 27916 7748 27956 7757
rect 27916 7412 27956 7708
rect 27916 7363 27956 7372
rect 27820 6691 27860 6700
rect 27916 6992 27956 7001
rect 27532 5935 27572 5944
rect 27436 5767 27476 5776
rect 27916 5816 27956 6952
rect 28204 6488 28244 6497
rect 28300 6488 28340 8884
rect 28588 8756 28628 9976
rect 28780 9596 28820 9605
rect 28588 8707 28628 8716
rect 28684 8840 28724 8849
rect 28492 8084 28532 8093
rect 28396 8000 28436 8009
rect 28396 7865 28436 7960
rect 28492 7496 28532 8044
rect 28588 8000 28628 8009
rect 28684 8000 28724 8800
rect 28628 7960 28724 8000
rect 28588 7951 28628 7960
rect 28780 7916 28820 9556
rect 28780 7867 28820 7876
rect 28492 7447 28532 7456
rect 28780 7160 28820 7169
rect 28244 6448 28340 6488
rect 28396 6488 28436 6497
rect 28204 6439 28244 6448
rect 28396 6068 28436 6448
rect 28396 6019 28436 6028
rect 28588 6068 28628 6077
rect 27916 5767 27956 5776
rect 27628 5648 27668 5657
rect 26764 5144 26804 5153
rect 26764 4808 26804 5104
rect 27628 5060 27668 5608
rect 27628 5011 27668 5020
rect 26764 4759 26804 4768
rect 28588 3632 28628 6028
rect 28780 5900 28820 7120
rect 28876 6488 28916 11764
rect 28972 9764 29012 9773
rect 28972 8000 29012 9724
rect 29068 9008 29108 9017
rect 29068 8672 29108 8968
rect 29068 8623 29108 8632
rect 28972 7951 29012 7960
rect 29260 6740 29300 11764
rect 29356 9008 29396 9017
rect 29356 8756 29396 8968
rect 29356 8707 29396 8716
rect 29452 8672 29492 8681
rect 29452 8537 29492 8632
rect 29644 7748 29684 11764
rect 30028 8168 30068 11764
rect 30220 9092 30260 9101
rect 30220 8957 30260 9052
rect 30028 8119 30068 8128
rect 30220 8588 30260 8597
rect 29644 7699 29684 7708
rect 29836 7748 29876 7757
rect 29836 7580 29876 7708
rect 29836 7531 29876 7540
rect 30028 7496 30068 7505
rect 30028 7361 30068 7456
rect 30220 7244 30260 8548
rect 30412 7412 30452 11764
rect 30796 11444 30836 11764
rect 31180 11528 31220 11764
rect 31564 11696 31604 11764
rect 31988 11764 32008 11780
rect 32312 11764 32392 11844
rect 32696 11764 32776 11844
rect 33080 11764 33160 11844
rect 33464 11764 33544 11844
rect 33848 11764 33928 11844
rect 34232 11764 34312 11844
rect 34616 11764 34696 11844
rect 35000 11764 35080 11844
rect 35384 11764 35464 11844
rect 35768 11764 35848 11844
rect 36152 11764 36232 11844
rect 36536 11764 36616 11844
rect 36920 11764 37000 11844
rect 37304 11764 37384 11844
rect 37688 11764 37768 11844
rect 38072 11780 38152 11844
rect 38072 11764 38092 11780
rect 31948 11731 31988 11740
rect 31564 11647 31604 11656
rect 31180 11479 31220 11488
rect 30796 11395 30836 11404
rect 31180 9848 31220 9857
rect 31084 9092 31124 9101
rect 30988 9008 31028 9017
rect 30988 8873 31028 8968
rect 31084 8504 31124 9052
rect 31180 8672 31220 9808
rect 31468 9176 31508 9185
rect 31372 9008 31412 9017
rect 31276 8924 31316 8933
rect 31276 8789 31316 8884
rect 31372 8873 31412 8968
rect 31468 8924 31508 9136
rect 31468 8875 31508 8884
rect 31180 8623 31220 8632
rect 31084 8455 31124 8464
rect 31852 8336 31892 8345
rect 31852 8201 31892 8296
rect 32332 7580 32372 11764
rect 32716 11612 32756 11764
rect 32716 11563 32756 11572
rect 33100 11444 33140 11764
rect 33100 11404 33236 11444
rect 32716 9428 32756 9437
rect 32716 8168 32756 9388
rect 33196 9344 33236 11404
rect 33196 9295 33236 9304
rect 32908 8504 32948 8513
rect 32716 8119 32756 8128
rect 32812 8420 32852 8429
rect 32812 8168 32852 8380
rect 32812 8119 32852 8128
rect 32908 7580 32948 8464
rect 33484 8336 33524 11764
rect 33868 10268 33908 11764
rect 34252 10604 34292 11764
rect 34252 10564 34388 10604
rect 33484 8287 33524 8296
rect 33772 10228 33908 10268
rect 33580 8252 33620 8261
rect 33292 8084 33332 8093
rect 33484 8084 33524 8093
rect 33332 8044 33484 8084
rect 33292 8035 33332 8044
rect 33484 8035 33524 8044
rect 33196 8000 33236 8009
rect 33196 7865 33236 7960
rect 33580 8000 33620 8212
rect 33580 7951 33620 7960
rect 33292 7832 33332 7841
rect 33292 7580 33332 7792
rect 32908 7540 33332 7580
rect 32332 7531 32372 7540
rect 30412 7363 30452 7372
rect 33772 7412 33812 10228
rect 33928 9848 34296 9857
rect 33968 9808 34010 9848
rect 34050 9808 34092 9848
rect 34132 9808 34174 9848
rect 34214 9808 34256 9848
rect 33928 9799 34296 9808
rect 34348 9428 34388 10564
rect 34636 9764 34676 11764
rect 34636 9715 34676 9724
rect 34348 9379 34388 9388
rect 35020 9344 35060 11764
rect 35020 9295 35060 9304
rect 35404 9260 35444 11764
rect 35788 10100 35828 11764
rect 35788 10051 35828 10060
rect 36172 9680 36212 11764
rect 36172 9631 36212 9640
rect 35404 9211 35444 9220
rect 35168 9092 35536 9101
rect 35208 9052 35250 9092
rect 35290 9052 35332 9092
rect 35372 9052 35414 9092
rect 35454 9052 35496 9092
rect 35168 9043 35536 9052
rect 35308 8588 35348 8597
rect 33928 8336 34296 8345
rect 33968 8296 34010 8336
rect 34050 8296 34092 8336
rect 34132 8296 34174 8336
rect 34214 8296 34256 8336
rect 33928 8287 34296 8296
rect 34636 8000 34676 8009
rect 33772 7363 33812 7372
rect 33868 7748 33908 7757
rect 33868 7328 33908 7708
rect 33868 7279 33908 7288
rect 34540 7496 34580 7505
rect 30220 7195 30260 7204
rect 33928 6824 34296 6833
rect 33968 6784 34010 6824
rect 34050 6784 34092 6824
rect 34132 6784 34174 6824
rect 34214 6784 34256 6824
rect 33928 6775 34296 6784
rect 29260 6691 29300 6700
rect 28876 6439 28916 6448
rect 29068 6656 29108 6665
rect 28780 5851 28820 5860
rect 28972 6236 29012 6245
rect 28972 5900 29012 6196
rect 28972 5851 29012 5860
rect 28588 3583 28628 3592
rect 28300 3464 28340 3473
rect 28300 3329 28340 3424
rect 29068 80 29108 6616
rect 31564 5900 31604 5909
rect 30028 5648 30068 5657
rect 29836 5396 29876 5405
rect 30028 5396 30068 5608
rect 29876 5356 30068 5396
rect 29836 5347 29876 5356
rect 30124 5312 30164 5321
rect 30124 4724 30164 5272
rect 30124 4675 30164 4684
rect 31180 4220 31220 4229
rect 31372 4220 31412 4229
rect 31220 4180 31372 4220
rect 31180 4171 31220 4180
rect 31372 4171 31412 4180
rect 31564 80 31604 5860
rect 33292 5648 33332 5657
rect 33100 5480 33140 5489
rect 33140 5440 33236 5480
rect 33100 5412 33140 5440
rect 33196 5144 33236 5440
rect 33292 5312 33332 5608
rect 33292 5263 33332 5272
rect 33928 5312 34296 5321
rect 33968 5272 34010 5312
rect 34050 5272 34092 5312
rect 34132 5272 34174 5312
rect 34214 5272 34256 5312
rect 33928 5263 34296 5272
rect 33196 5095 33236 5104
rect 32428 4976 32468 4985
rect 32428 4556 32468 4936
rect 32428 4507 32468 4516
rect 32620 4976 32660 4985
rect 32620 4388 32660 4936
rect 32620 4339 32660 4348
rect 33928 3800 34296 3809
rect 33968 3760 34010 3800
rect 34050 3760 34092 3800
rect 34132 3760 34174 3800
rect 34214 3760 34256 3800
rect 33928 3751 34296 3760
rect 33928 2288 34296 2297
rect 33968 2248 34010 2288
rect 34050 2248 34092 2288
rect 34132 2248 34174 2288
rect 34214 2248 34256 2288
rect 33928 2239 34296 2248
rect 34060 104 34100 113
rect 1592 0 1672 80
rect 4088 0 4168 80
rect 6584 0 6664 80
rect 9080 0 9160 80
rect 11576 0 11656 80
rect 14072 0 14152 80
rect 16568 0 16648 80
rect 19064 0 19144 80
rect 21560 0 21640 80
rect 24056 0 24136 80
rect 26552 0 26632 80
rect 29048 0 29128 80
rect 31544 0 31624 80
rect 34040 64 34060 80
rect 34348 104 34388 113
rect 34100 64 34120 80
rect 34040 0 34120 64
rect 34348 60 34388 64
rect 34540 60 34580 7456
rect 34636 7412 34676 7960
rect 34636 7363 34676 7372
rect 34924 8000 34964 8009
rect 34924 7412 34964 7960
rect 35308 8000 35348 8548
rect 35404 8252 35444 8261
rect 35404 8084 35444 8212
rect 36556 8168 36596 11764
rect 36940 9932 36980 11764
rect 36940 9892 37268 9932
rect 36556 8119 36596 8128
rect 36940 9512 36980 9521
rect 36940 8168 36980 9472
rect 36940 8119 36980 8128
rect 37132 8504 37172 8513
rect 35404 8035 35444 8044
rect 35308 7951 35348 7960
rect 36556 8000 36596 8009
rect 35168 7580 35536 7589
rect 35208 7540 35250 7580
rect 35290 7540 35332 7580
rect 35372 7540 35414 7580
rect 35454 7540 35496 7580
rect 35168 7531 35536 7540
rect 34924 7363 34964 7372
rect 34732 6404 34772 6413
rect 34772 6364 35060 6404
rect 34732 6355 34772 6364
rect 34732 6236 34772 6245
rect 34732 6101 34772 6196
rect 35020 6152 35060 6364
rect 35116 6236 35156 6331
rect 35116 6187 35156 6196
rect 35020 6103 35060 6112
rect 35168 6068 35536 6077
rect 35208 6028 35250 6068
rect 35290 6028 35332 6068
rect 35372 6028 35414 6068
rect 35454 6028 35496 6068
rect 35168 6019 35536 6028
rect 35168 4556 35536 4565
rect 35208 4516 35250 4556
rect 35290 4516 35332 4556
rect 35372 4516 35414 4556
rect 35454 4516 35496 4556
rect 35168 4507 35536 4516
rect 35168 3044 35536 3053
rect 35208 3004 35250 3044
rect 35290 3004 35332 3044
rect 35372 3004 35414 3044
rect 35454 3004 35496 3044
rect 35168 2995 35536 3004
rect 35168 1532 35536 1541
rect 35208 1492 35250 1532
rect 35290 1492 35332 1532
rect 35372 1492 35414 1532
rect 35454 1492 35496 1532
rect 35168 1483 35536 1492
rect 36556 80 36596 7960
rect 36748 8000 36788 8009
rect 36748 7580 36788 7960
rect 37132 7748 37172 8464
rect 37228 8000 37268 9892
rect 37324 9092 37364 11764
rect 37324 9043 37364 9052
rect 37612 8504 37652 8513
rect 37420 8168 37460 8177
rect 37420 8033 37460 8128
rect 37612 8084 37652 8464
rect 37708 8336 37748 11764
rect 38132 11764 38152 11780
rect 38284 11780 38324 11789
rect 38092 11731 38132 11740
rect 38456 11764 38536 11844
rect 38840 11764 38920 11844
rect 39224 11764 39304 11844
rect 39608 11764 39688 11844
rect 39992 11764 40072 11844
rect 40376 11764 40456 11844
rect 40760 11764 40840 11844
rect 41144 11764 41224 11844
rect 41528 11764 41608 11844
rect 41912 11764 41992 11844
rect 42296 11764 42376 11844
rect 42680 11764 42760 11844
rect 43064 11764 43144 11844
rect 43448 11764 43528 11844
rect 43832 11764 43912 11844
rect 44216 11764 44296 11844
rect 44600 11764 44680 11844
rect 44984 11764 45064 11844
rect 45368 11764 45448 11844
rect 45752 11764 45832 11844
rect 46136 11764 46216 11844
rect 46520 11764 46600 11844
rect 46904 11764 46984 11844
rect 47288 11764 47368 11844
rect 47672 11764 47752 11844
rect 48056 11764 48136 11844
rect 48440 11764 48520 11844
rect 48824 11764 48904 11844
rect 49208 11764 49288 11844
rect 49592 11764 49672 11844
rect 49976 11764 50056 11844
rect 50360 11764 50440 11844
rect 37996 9092 38036 9101
rect 37996 8672 38036 9052
rect 37996 8623 38036 8632
rect 38188 8924 38228 8933
rect 38188 8672 38228 8884
rect 38188 8623 38228 8632
rect 37708 8287 37748 8296
rect 37804 8420 37844 8429
rect 37612 8035 37652 8044
rect 37804 8084 37844 8380
rect 37804 8035 37844 8044
rect 37900 8168 37940 8177
rect 37228 7951 37268 7960
rect 37324 7748 37364 7757
rect 37132 7708 37324 7748
rect 37324 7699 37364 7708
rect 36748 7531 36788 7540
rect 37900 7496 37940 8128
rect 37900 7447 37940 7456
rect 38284 7244 38324 11740
rect 38380 9092 38420 9101
rect 38380 8000 38420 9052
rect 38380 7951 38420 7960
rect 38476 7832 38516 11764
rect 38860 8168 38900 11764
rect 38860 8119 38900 8128
rect 39052 8336 39092 8345
rect 39052 8000 39092 8296
rect 39244 8084 39284 11764
rect 39628 8420 39668 11764
rect 40012 8504 40052 11764
rect 40012 8455 40052 8464
rect 40300 9512 40340 9521
rect 39628 8371 39668 8380
rect 39340 8336 39380 8347
rect 39340 8252 39380 8296
rect 39340 8203 39380 8212
rect 39244 8035 39284 8044
rect 39436 8084 39476 8093
rect 39052 7951 39092 7960
rect 39436 7949 39476 8044
rect 39724 8084 39764 8095
rect 39724 8000 39764 8044
rect 39724 7951 39764 7960
rect 39628 7916 39668 7925
rect 38476 7783 38516 7792
rect 38860 7832 38900 7843
rect 39628 7832 39668 7876
rect 39820 7832 39860 7841
rect 39628 7792 39820 7832
rect 38860 7748 38900 7792
rect 39820 7783 39860 7792
rect 38860 7699 38900 7708
rect 39532 7748 39572 7757
rect 39532 7613 39572 7708
rect 39052 7580 39092 7589
rect 38956 7412 38996 7421
rect 38956 7277 38996 7372
rect 38284 7195 38324 7204
rect 37228 7160 37268 7169
rect 37228 7025 37268 7120
rect 37804 7160 37844 7169
rect 37324 7076 37364 7085
rect 37324 6656 37364 7036
rect 37804 6908 37844 7120
rect 37804 6859 37844 6868
rect 38092 7160 38132 7169
rect 37324 6607 37364 6616
rect 38092 5900 38132 7120
rect 38956 7076 38996 7085
rect 38956 6941 38996 7036
rect 38092 5851 38132 5860
rect 38092 5732 38132 5741
rect 38092 5228 38132 5692
rect 38092 5179 38132 5188
rect 39052 80 39092 7540
rect 39148 7244 39188 7253
rect 39148 7109 39188 7204
rect 39244 7160 39284 7169
rect 39244 7025 39284 7120
rect 39340 7076 39380 7085
rect 39340 6941 39380 7036
rect 40300 5564 40340 9472
rect 40396 8588 40436 11764
rect 40588 9428 40628 9437
rect 40396 8539 40436 8548
rect 40492 9344 40532 9353
rect 40492 6740 40532 9304
rect 40492 6691 40532 6700
rect 40588 6152 40628 9388
rect 40780 7412 40820 11764
rect 41164 7496 41204 11764
rect 41548 8336 41588 11764
rect 41548 8287 41588 8296
rect 41740 9260 41780 9269
rect 41164 7447 41204 7456
rect 40780 7363 40820 7372
rect 40972 7076 41012 7085
rect 41012 7036 41204 7076
rect 40972 7027 41012 7036
rect 41164 6992 41204 7036
rect 41164 6943 41204 6952
rect 40588 6103 40628 6112
rect 41548 6488 41588 6497
rect 40300 5515 40340 5524
rect 40492 5564 40532 5573
rect 40492 4808 40532 5524
rect 40492 4759 40532 4768
rect 41548 80 41588 6448
rect 41740 5648 41780 9220
rect 41740 5599 41780 5608
rect 41836 9176 41876 9185
rect 41836 5060 41876 9136
rect 41932 8084 41972 11764
rect 42316 9092 42356 11764
rect 42700 9680 42740 11764
rect 42700 9631 42740 9640
rect 43084 9680 43124 11764
rect 43084 9631 43124 9640
rect 43468 9680 43508 11764
rect 43468 9631 43508 9640
rect 43852 9680 43892 11764
rect 43852 9631 43892 9640
rect 44236 9680 44276 11764
rect 44236 9631 44276 9640
rect 44620 9680 44660 11764
rect 44620 9631 44660 9640
rect 45004 9680 45044 11764
rect 45004 9631 45044 9640
rect 45388 9680 45428 11764
rect 45388 9631 45428 9640
rect 45772 9680 45812 11764
rect 45772 9631 45812 9640
rect 46156 9680 46196 11764
rect 46156 9631 46196 9640
rect 46540 9680 46580 11764
rect 46540 9631 46580 9640
rect 46924 9680 46964 11764
rect 46924 9631 46964 9640
rect 47116 9764 47156 9773
rect 46060 9512 46100 9521
rect 43180 9428 43220 9437
rect 43084 9388 43180 9428
rect 42316 9043 42356 9052
rect 42604 9092 42644 9101
rect 41932 8035 41972 8044
rect 42604 6572 42644 9052
rect 42604 6523 42644 6532
rect 43084 6236 43124 9388
rect 43180 9360 43220 9388
rect 44236 9428 44276 9437
rect 43084 6187 43124 6196
rect 44044 6488 44084 6497
rect 41836 5011 41876 5020
rect 43084 1868 43124 1877
rect 43276 1868 43316 1877
rect 43124 1828 43276 1868
rect 43084 1819 43124 1828
rect 43276 1819 43316 1828
rect 44044 80 44084 6448
rect 44236 5144 44276 9388
rect 44236 5095 44276 5104
rect 46060 4724 46100 9472
rect 46444 9512 46484 9521
rect 46444 5480 46484 9472
rect 46828 9512 46868 9521
rect 46732 9344 46772 9353
rect 46444 5431 46484 5440
rect 46540 5648 46580 5657
rect 46060 4675 46100 4684
rect 45292 2036 45332 2045
rect 45292 1784 45332 1996
rect 45292 1735 45332 1744
rect 46540 80 46580 5608
rect 46732 5648 46772 9304
rect 46828 6320 46868 9472
rect 47116 8840 47156 9724
rect 47308 9680 47348 11764
rect 47308 9631 47348 9640
rect 47692 9680 47732 11764
rect 47692 9631 47732 9640
rect 48076 9680 48116 11764
rect 48076 9631 48116 9640
rect 48460 9680 48500 11764
rect 48460 9631 48500 9640
rect 48844 9680 48884 11764
rect 49228 10016 49268 11764
rect 49228 9976 49556 10016
rect 49048 9848 49416 9857
rect 49088 9808 49130 9848
rect 49170 9808 49212 9848
rect 49252 9808 49294 9848
rect 49334 9808 49376 9848
rect 49048 9799 49416 9808
rect 48844 9631 48884 9640
rect 49516 9680 49556 9976
rect 49516 9631 49556 9640
rect 49612 9596 49652 11764
rect 49996 9680 50036 11764
rect 49996 9631 50036 9640
rect 50380 9680 50420 11764
rect 50860 11024 50900 11033
rect 50380 9631 50420 9640
rect 50764 10688 50804 10697
rect 49612 9547 49652 9556
rect 47116 8791 47156 8800
rect 47212 9512 47252 9521
rect 47404 9512 47444 9521
rect 47212 6908 47252 9472
rect 47308 9472 47404 9512
rect 47308 6992 47348 9472
rect 47404 9463 47444 9472
rect 47980 9512 48020 9521
rect 47308 6943 47348 6952
rect 47404 8840 47444 8849
rect 47212 6859 47252 6868
rect 47404 6824 47444 8800
rect 47980 8252 48020 9472
rect 47980 8203 48020 8212
rect 48364 9512 48404 9521
rect 47404 6775 47444 6784
rect 47500 8084 47540 8093
rect 46828 6271 46868 6280
rect 47308 6572 47348 6581
rect 47308 5900 47348 6532
rect 47500 5984 47540 8044
rect 48364 7664 48404 9472
rect 48748 9512 48788 9521
rect 48748 7832 48788 9472
rect 48940 9512 48980 9521
rect 48940 8756 48980 9472
rect 48940 8707 48980 8716
rect 49036 9512 49076 9521
rect 49036 8504 49076 9472
rect 50092 9512 50132 9521
rect 48748 7783 48788 7792
rect 48940 8464 49076 8504
rect 49996 9428 50036 9437
rect 48364 7615 48404 7624
rect 48940 6656 48980 8464
rect 49048 8336 49416 8345
rect 49088 8296 49130 8336
rect 49170 8296 49212 8336
rect 49252 8296 49294 8336
rect 49334 8296 49376 8336
rect 49048 8287 49416 8296
rect 49048 6824 49416 6833
rect 49088 6784 49130 6824
rect 49170 6784 49212 6824
rect 49252 6784 49294 6824
rect 49334 6784 49376 6824
rect 49048 6775 49416 6784
rect 48940 6607 48980 6616
rect 47500 5935 47540 5944
rect 48940 6488 48980 6497
rect 47308 5851 47348 5860
rect 46732 5599 46772 5608
rect 47308 4136 47348 4145
rect 47308 3464 47348 4096
rect 47308 3415 47348 3424
rect 48940 1448 48980 6448
rect 49996 5648 50036 9388
rect 50092 6656 50132 9472
rect 50188 9092 50228 9101
rect 50188 8672 50228 9052
rect 50288 9092 50656 9101
rect 50328 9052 50370 9092
rect 50410 9052 50452 9092
rect 50492 9052 50534 9092
rect 50574 9052 50616 9092
rect 50288 9043 50656 9052
rect 50764 8924 50804 10648
rect 50860 9008 50900 10984
rect 52300 10352 52340 10361
rect 50860 8959 50900 8968
rect 50956 10016 50996 10025
rect 50764 8875 50804 8884
rect 50284 8672 50324 8681
rect 50188 8632 50284 8672
rect 50284 8623 50324 8632
rect 50956 8672 50996 9976
rect 51148 10016 51188 10025
rect 51052 9512 51092 9521
rect 51052 9377 51092 9472
rect 51052 8924 51092 8933
rect 51148 8924 51188 9976
rect 51092 8884 51188 8924
rect 51052 8875 51092 8884
rect 50956 8623 50996 8632
rect 51436 8672 51476 8681
rect 51436 8537 51476 8632
rect 52300 8168 52340 10312
rect 52684 9260 52724 9269
rect 52684 8672 52724 9220
rect 52684 8623 52724 8632
rect 52300 8119 52340 8128
rect 52684 8504 52724 8513
rect 51916 8000 51956 8009
rect 50288 7580 50656 7589
rect 50328 7540 50370 7580
rect 50410 7540 50452 7580
rect 50492 7540 50534 7580
rect 50574 7540 50616 7580
rect 50288 7531 50656 7540
rect 50092 6607 50132 6616
rect 51820 7160 51860 7169
rect 50288 6068 50656 6077
rect 50328 6028 50370 6068
rect 50410 6028 50452 6068
rect 50492 6028 50534 6068
rect 50574 6028 50616 6068
rect 50288 6019 50656 6028
rect 51820 5816 51860 7120
rect 51916 5984 51956 7960
rect 52684 8000 52724 8464
rect 52684 7951 52724 7960
rect 52684 7748 52724 7757
rect 52684 7328 52724 7708
rect 52684 7279 52724 7288
rect 51916 5935 51956 5944
rect 51820 5767 51860 5776
rect 49996 5599 50036 5608
rect 51532 5732 51572 5741
rect 49048 5312 49416 5321
rect 49088 5272 49130 5312
rect 49170 5272 49212 5312
rect 49252 5272 49294 5312
rect 49334 5272 49376 5312
rect 49048 5263 49416 5272
rect 50288 4556 50656 4565
rect 50328 4516 50370 4556
rect 50410 4516 50452 4556
rect 50492 4516 50534 4556
rect 50574 4516 50616 4556
rect 50288 4507 50656 4516
rect 49048 3800 49416 3809
rect 49088 3760 49130 3800
rect 49170 3760 49212 3800
rect 49252 3760 49294 3800
rect 49334 3760 49376 3800
rect 49048 3751 49416 3760
rect 50288 3044 50656 3053
rect 50328 3004 50370 3044
rect 50410 3004 50452 3044
rect 50492 3004 50534 3044
rect 50574 3004 50616 3044
rect 50288 2995 50656 3004
rect 50380 2372 50420 2381
rect 49048 2288 49416 2297
rect 49088 2248 49130 2288
rect 49170 2248 49212 2288
rect 49252 2248 49294 2288
rect 49334 2248 49376 2288
rect 49048 2239 49416 2248
rect 50380 1952 50420 2332
rect 50380 1903 50420 1912
rect 50572 1868 50612 1877
rect 50764 1868 50804 1877
rect 50612 1828 50764 1868
rect 50572 1819 50612 1828
rect 50764 1819 50804 1828
rect 50288 1532 50656 1541
rect 50328 1492 50370 1532
rect 50410 1492 50452 1532
rect 50492 1492 50534 1532
rect 50574 1492 50616 1532
rect 50288 1483 50656 1492
rect 48940 1408 49076 1448
rect 49036 80 49076 1408
rect 51532 80 51572 5692
rect 51820 5648 51860 5657
rect 51820 4808 51860 5608
rect 51820 4759 51860 4768
rect 51820 4220 51860 4229
rect 51820 3464 51860 4180
rect 51820 3415 51860 3424
rect 52300 1868 52340 1877
rect 52300 608 52340 1828
rect 52972 1784 53012 1793
rect 52972 944 53012 1744
rect 53164 1448 53204 1457
rect 53164 1280 53204 1408
rect 53164 1231 53204 1240
rect 52972 895 53012 904
rect 52300 559 52340 568
rect 34348 20 34580 60
rect 36536 0 36616 80
rect 39032 0 39112 80
rect 41528 0 41608 80
rect 44024 0 44104 80
rect 46520 0 46600 80
rect 49016 0 49096 80
rect 51512 0 51592 80
<< via3 >>
rect 556 8800 596 8840
rect 1420 9976 1460 10016
rect 3688 9808 3728 9848
rect 3770 9808 3810 9848
rect 3852 9808 3892 9848
rect 3934 9808 3974 9848
rect 4016 9808 4056 9848
rect 1228 8884 1268 8924
rect 1420 8968 1460 9008
rect 748 8632 788 8672
rect 3688 8296 3728 8336
rect 3770 8296 3810 8336
rect 3852 8296 3892 8336
rect 3934 8296 3974 8336
rect 4016 8296 4056 8336
rect 4588 9220 4628 9260
rect 4928 9052 4968 9092
rect 5010 9052 5050 9092
rect 5092 9052 5132 9092
rect 5174 9052 5214 9092
rect 5256 9052 5296 9092
rect 268 7960 308 8000
rect 940 4096 980 4136
rect 4928 7540 4968 7580
rect 5010 7540 5050 7580
rect 5092 7540 5132 7580
rect 5174 7540 5214 7580
rect 5256 7540 5296 7580
rect 3688 6784 3728 6824
rect 3770 6784 3810 6824
rect 3852 6784 3892 6824
rect 3934 6784 3974 6824
rect 4016 6784 4056 6824
rect 8620 9304 8660 9344
rect 10060 8380 10100 8420
rect 10060 7876 10100 7916
rect 13228 9892 13268 9932
rect 11116 9472 11156 9512
rect 12844 8380 12884 8420
rect 14188 9472 14228 9512
rect 14380 9472 14420 9512
rect 1420 3424 1460 3464
rect 3688 5272 3728 5312
rect 3770 5272 3810 5312
rect 3852 5272 3892 5312
rect 3934 5272 3974 5312
rect 4016 5272 4056 5312
rect 3688 3760 3728 3800
rect 3770 3760 3810 3800
rect 3852 3760 3892 3800
rect 3934 3760 3974 3800
rect 4016 3760 4056 3800
rect 3688 2248 3728 2288
rect 3770 2248 3810 2288
rect 3852 2248 3892 2288
rect 3934 2248 3974 2288
rect 4016 2248 4056 2288
rect 4928 6028 4968 6068
rect 5010 6028 5050 6068
rect 5092 6028 5132 6068
rect 5174 6028 5214 6068
rect 5256 6028 5296 6068
rect 4928 4516 4968 4556
rect 5010 4516 5050 4556
rect 5092 4516 5132 4556
rect 5174 4516 5214 4556
rect 5256 4516 5296 4556
rect 4928 3004 4968 3044
rect 5010 3004 5050 3044
rect 5092 3004 5132 3044
rect 5174 3004 5214 3044
rect 5256 3004 5296 3044
rect 4928 1492 4968 1532
rect 5010 1492 5050 1532
rect 5092 1492 5132 1532
rect 5174 1492 5214 1532
rect 5256 1492 5296 1532
rect 14380 8380 14420 8420
rect 15628 9220 15668 9260
rect 15340 8464 15380 8504
rect 15820 8548 15860 8588
rect 16300 9892 16340 9932
rect 16684 7876 16724 7916
rect 17836 9388 17876 9428
rect 17452 8716 17492 8756
rect 17836 8716 17876 8756
rect 17644 7708 17684 7748
rect 18808 9808 18848 9848
rect 18890 9808 18930 9848
rect 18972 9808 19012 9848
rect 19054 9808 19094 9848
rect 19136 9808 19176 9848
rect 19276 9388 19316 9428
rect 18988 8716 19028 8756
rect 18808 8296 18848 8336
rect 18890 8296 18930 8336
rect 18972 8296 19012 8336
rect 19054 8296 19094 8336
rect 19136 8296 19176 8336
rect 19564 8212 19604 8252
rect 20140 9724 20180 9764
rect 20908 9808 20948 9848
rect 20524 9136 20564 9176
rect 20048 9052 20088 9092
rect 20130 9052 20170 9092
rect 20212 9052 20252 9092
rect 20294 9052 20334 9092
rect 20376 9052 20416 9092
rect 20044 8716 20084 8756
rect 20140 8296 20180 8336
rect 20428 8380 20468 8420
rect 20332 8296 20372 8336
rect 20048 7540 20088 7580
rect 20130 7540 20170 7580
rect 20212 7540 20252 7580
rect 20294 7540 20334 7580
rect 20376 7540 20416 7580
rect 19660 7456 19700 7496
rect 21004 9388 21044 9428
rect 21196 7708 21236 7748
rect 21676 7792 21716 7832
rect 22252 9556 22292 9596
rect 22156 9220 22196 9260
rect 23020 9052 23060 9092
rect 21772 7708 21812 7748
rect 23884 9808 23924 9848
rect 24940 9556 24980 9596
rect 25420 9472 25460 9512
rect 24556 9220 24596 9260
rect 25036 9304 25076 9344
rect 25228 9304 25268 9344
rect 25324 9136 25364 9176
rect 18808 6784 18848 6824
rect 18890 6784 18930 6824
rect 18972 6784 19012 6824
rect 19054 6784 19094 6824
rect 19136 6784 19176 6824
rect 20048 6028 20088 6068
rect 20130 6028 20170 6068
rect 20212 6028 20252 6068
rect 20294 6028 20334 6068
rect 20376 6028 20416 6068
rect 23116 6028 23156 6068
rect 25804 8464 25844 8504
rect 23404 6532 23444 6572
rect 25708 6532 25748 6572
rect 23788 6028 23828 6068
rect 18808 5272 18848 5312
rect 18890 5272 18930 5312
rect 18972 5272 19012 5312
rect 19054 5272 19094 5312
rect 19136 5272 19176 5312
rect 18808 3760 18848 3800
rect 18890 3760 18930 3800
rect 18972 3760 19012 3800
rect 19054 3760 19094 3800
rect 19136 3760 19176 3800
rect 18808 2248 18848 2288
rect 18890 2248 18930 2288
rect 18972 2248 19012 2288
rect 19054 2248 19094 2288
rect 19136 2248 19176 2288
rect 20048 4516 20088 4556
rect 20130 4516 20170 4556
rect 20212 4516 20252 4556
rect 20294 4516 20334 4556
rect 20376 4516 20416 4556
rect 20048 3004 20088 3044
rect 20130 3004 20170 3044
rect 20212 3004 20252 3044
rect 20294 3004 20334 3044
rect 20376 3004 20416 3044
rect 20048 1492 20088 1532
rect 20130 1492 20170 1532
rect 20212 1492 20252 1532
rect 20294 1492 20334 1532
rect 20376 1492 20416 1532
rect 25996 4096 26036 4136
rect 26764 8548 26804 8588
rect 27148 8884 27188 8924
rect 27532 8800 27572 8840
rect 28012 9976 28052 10016
rect 28108 8380 28148 8420
rect 28684 8800 28724 8840
rect 28396 7960 28436 8000
rect 28492 7456 28532 7496
rect 28972 9724 29012 9764
rect 29068 8968 29108 9008
rect 29356 8716 29396 8756
rect 29452 8632 29492 8672
rect 30220 9052 30260 9092
rect 29836 7540 29876 7580
rect 30028 7456 30068 7496
rect 30988 8968 31028 9008
rect 31372 8968 31412 9008
rect 31276 8884 31316 8924
rect 31852 8296 31892 8336
rect 33196 9304 33236 9344
rect 32812 8128 32852 8168
rect 33484 8296 33524 8336
rect 33580 8212 33620 8252
rect 33196 7960 33236 8000
rect 33928 9808 33968 9848
rect 34010 9808 34050 9848
rect 34092 9808 34132 9848
rect 34174 9808 34214 9848
rect 34256 9808 34296 9848
rect 34348 9388 34388 9428
rect 35168 9052 35208 9092
rect 35250 9052 35290 9092
rect 35332 9052 35372 9092
rect 35414 9052 35454 9092
rect 35496 9052 35536 9092
rect 33928 8296 33968 8336
rect 34010 8296 34050 8336
rect 34092 8296 34132 8336
rect 34174 8296 34214 8336
rect 34256 8296 34296 8336
rect 33928 6784 33968 6824
rect 34010 6784 34050 6824
rect 34092 6784 34132 6824
rect 34174 6784 34214 6824
rect 34256 6784 34296 6824
rect 28300 3424 28340 3464
rect 31564 5860 31604 5900
rect 33928 5272 33968 5312
rect 34010 5272 34050 5312
rect 34092 5272 34132 5312
rect 34174 5272 34214 5312
rect 34256 5272 34296 5312
rect 33928 3760 33968 3800
rect 34010 3760 34050 3800
rect 34092 3760 34132 3800
rect 34174 3760 34214 3800
rect 34256 3760 34296 3800
rect 33928 2248 33968 2288
rect 34010 2248 34050 2288
rect 34092 2248 34132 2288
rect 34174 2248 34214 2288
rect 34256 2248 34296 2288
rect 34060 64 34100 104
rect 34348 64 34388 104
rect 35404 8044 35444 8084
rect 35168 7540 35208 7580
rect 35250 7540 35290 7580
rect 35332 7540 35372 7580
rect 35414 7540 35454 7580
rect 35496 7540 35536 7580
rect 34924 7372 34964 7412
rect 34732 6196 34772 6236
rect 35116 6196 35156 6236
rect 35168 6028 35208 6068
rect 35250 6028 35290 6068
rect 35332 6028 35372 6068
rect 35414 6028 35454 6068
rect 35496 6028 35536 6068
rect 35168 4516 35208 4556
rect 35250 4516 35290 4556
rect 35332 4516 35372 4556
rect 35414 4516 35454 4556
rect 35496 4516 35536 4556
rect 35168 3004 35208 3044
rect 35250 3004 35290 3044
rect 35332 3004 35372 3044
rect 35414 3004 35454 3044
rect 35496 3004 35536 3044
rect 35168 1492 35208 1532
rect 35250 1492 35290 1532
rect 35332 1492 35372 1532
rect 35414 1492 35454 1532
rect 35496 1492 35536 1532
rect 37324 9052 37364 9092
rect 37420 8128 37460 8168
rect 38092 11740 38132 11780
rect 38284 11740 38324 11780
rect 38188 8884 38228 8924
rect 38380 9052 38420 9092
rect 39340 8212 39380 8252
rect 39436 8044 39476 8084
rect 39724 7960 39764 8000
rect 38860 7792 38900 7832
rect 39532 7708 39572 7748
rect 38956 7372 38996 7412
rect 38284 7204 38324 7244
rect 37228 7120 37268 7160
rect 38956 7036 38996 7076
rect 38092 5860 38132 5900
rect 39148 7204 39188 7244
rect 39244 7120 39284 7160
rect 39340 7036 39380 7076
rect 49048 9808 49088 9848
rect 49130 9808 49170 9848
rect 49212 9808 49252 9848
rect 49294 9808 49334 9848
rect 49376 9808 49416 9848
rect 48940 9472 48980 9512
rect 48940 8716 48980 8756
rect 49048 8296 49088 8336
rect 49130 8296 49170 8336
rect 49212 8296 49252 8336
rect 49294 8296 49334 8336
rect 49376 8296 49416 8336
rect 49048 6784 49088 6824
rect 49130 6784 49170 6824
rect 49212 6784 49252 6824
rect 49294 6784 49334 6824
rect 49376 6784 49416 6824
rect 50288 9052 50328 9092
rect 50370 9052 50410 9092
rect 50452 9052 50492 9092
rect 50534 9052 50574 9092
rect 50616 9052 50656 9092
rect 51052 9472 51092 9512
rect 51436 8632 51476 8672
rect 50288 7540 50328 7580
rect 50370 7540 50410 7580
rect 50452 7540 50492 7580
rect 50534 7540 50574 7580
rect 50616 7540 50656 7580
rect 50288 6028 50328 6068
rect 50370 6028 50410 6068
rect 50452 6028 50492 6068
rect 50534 6028 50574 6068
rect 50616 6028 50656 6068
rect 49048 5272 49088 5312
rect 49130 5272 49170 5312
rect 49212 5272 49252 5312
rect 49294 5272 49334 5312
rect 49376 5272 49416 5312
rect 50288 4516 50328 4556
rect 50370 4516 50410 4556
rect 50452 4516 50492 4556
rect 50534 4516 50574 4556
rect 50616 4516 50656 4556
rect 49048 3760 49088 3800
rect 49130 3760 49170 3800
rect 49212 3760 49252 3800
rect 49294 3760 49334 3800
rect 49376 3760 49416 3800
rect 50288 3004 50328 3044
rect 50370 3004 50410 3044
rect 50452 3004 50492 3044
rect 50534 3004 50574 3044
rect 50616 3004 50656 3044
rect 49048 2248 49088 2288
rect 49130 2248 49170 2288
rect 49212 2248 49252 2288
rect 49294 2248 49334 2288
rect 49376 2248 49416 2288
rect 50288 1492 50328 1532
rect 50370 1492 50410 1532
rect 50452 1492 50492 1532
rect 50534 1492 50574 1532
rect 50616 1492 50656 1532
<< metal4 >>
rect 38083 11740 38092 11780
rect 38132 11740 38284 11780
rect 38324 11740 38333 11780
rect 1411 9976 1420 10016
rect 1460 9976 28012 10016
rect 28052 9976 28061 10016
rect 13219 9892 13228 9932
rect 13268 9892 16300 9932
rect 16340 9892 16349 9932
rect 3679 9808 3688 9848
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 4056 9808 4065 9848
rect 18799 9808 18808 9848
rect 18848 9808 18890 9848
rect 18930 9808 18972 9848
rect 19012 9808 19054 9848
rect 19094 9808 19136 9848
rect 19176 9808 19185 9848
rect 20899 9808 20908 9848
rect 20948 9808 23884 9848
rect 23924 9808 23933 9848
rect 33919 9808 33928 9848
rect 33968 9808 34010 9848
rect 34050 9808 34092 9848
rect 34132 9808 34174 9848
rect 34214 9808 34256 9848
rect 34296 9808 34305 9848
rect 49039 9808 49048 9848
rect 49088 9808 49130 9848
rect 49170 9808 49212 9848
rect 49252 9808 49294 9848
rect 49334 9808 49376 9848
rect 49416 9808 49425 9848
rect 20131 9724 20140 9764
rect 20180 9724 28972 9764
rect 29012 9724 29021 9764
rect 22243 9556 22252 9596
rect 22292 9556 24940 9596
rect 24980 9556 24989 9596
rect 11107 9472 11116 9512
rect 11156 9472 14188 9512
rect 14228 9472 14237 9512
rect 14371 9472 14380 9512
rect 14420 9472 25420 9512
rect 25460 9472 25469 9512
rect 48931 9472 48940 9512
rect 48980 9472 51052 9512
rect 51092 9472 51101 9512
rect 17827 9388 17836 9428
rect 17876 9388 19276 9428
rect 19316 9388 19325 9428
rect 20995 9388 21004 9428
rect 21044 9388 34348 9428
rect 34388 9388 34397 9428
rect 8611 9304 8620 9344
rect 8660 9304 25036 9344
rect 25076 9304 25085 9344
rect 25219 9304 25228 9344
rect 25268 9304 33196 9344
rect 33236 9304 33245 9344
rect 4579 9220 4588 9260
rect 4628 9220 15628 9260
rect 15668 9220 15677 9260
rect 22147 9220 22156 9260
rect 22196 9220 24556 9260
rect 24596 9220 24605 9260
rect 20515 9136 20524 9176
rect 20564 9136 25324 9176
rect 25364 9136 25373 9176
rect 4919 9052 4928 9092
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 5296 9052 5305 9092
rect 20039 9052 20048 9092
rect 20088 9052 20130 9092
rect 20170 9052 20212 9092
rect 20252 9052 20294 9092
rect 20334 9052 20376 9092
rect 20416 9052 20425 9092
rect 23011 9052 23020 9092
rect 23060 9052 30220 9092
rect 30260 9052 30269 9092
rect 35159 9052 35168 9092
rect 35208 9052 35250 9092
rect 35290 9052 35332 9092
rect 35372 9052 35414 9092
rect 35454 9052 35496 9092
rect 35536 9052 35545 9092
rect 37315 9052 37324 9092
rect 37364 9052 38380 9092
rect 38420 9052 38429 9092
rect 50279 9052 50288 9092
rect 50328 9052 50370 9092
rect 50410 9052 50452 9092
rect 50492 9052 50534 9092
rect 50574 9052 50616 9092
rect 50656 9052 50665 9092
rect 1411 8968 1420 9008
rect 1460 8968 29068 9008
rect 29108 8968 29117 9008
rect 30979 8968 30988 9008
rect 31028 8968 31372 9008
rect 31412 8968 31421 9008
rect 1219 8884 1228 8924
rect 1268 8884 27148 8924
rect 27188 8884 27197 8924
rect 31267 8884 31276 8924
rect 31316 8884 38188 8924
rect 38228 8884 38237 8924
rect 547 8800 556 8840
rect 596 8800 27532 8840
rect 27572 8800 27581 8840
rect 28675 8800 28684 8840
rect 28724 8800 33140 8840
rect 33100 8756 33140 8800
rect 17443 8716 17452 8756
rect 17492 8716 17836 8756
rect 17876 8716 17885 8756
rect 18979 8716 18988 8756
rect 19028 8716 20044 8756
rect 20084 8716 20093 8756
rect 29347 8716 29356 8756
rect 29396 8716 30068 8756
rect 33100 8716 48940 8756
rect 48980 8716 48989 8756
rect 30028 8672 30068 8716
rect 739 8632 748 8672
rect 788 8632 29452 8672
rect 29492 8632 29501 8672
rect 30028 8632 51436 8672
rect 51476 8632 51485 8672
rect 15811 8548 15820 8588
rect 15860 8548 26764 8588
rect 26804 8548 26813 8588
rect 15331 8464 15340 8504
rect 15380 8464 25804 8504
rect 25844 8464 25853 8504
rect 10051 8380 10060 8420
rect 10100 8380 10109 8420
rect 12835 8380 12844 8420
rect 12884 8380 14380 8420
rect 14420 8380 14429 8420
rect 20419 8380 20428 8420
rect 20468 8380 28108 8420
rect 28148 8380 28157 8420
rect 3679 8296 3688 8336
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 4056 8296 4065 8336
rect 10060 8252 10100 8380
rect 18799 8296 18808 8336
rect 18848 8296 18890 8336
rect 18930 8296 18972 8336
rect 19012 8296 19054 8336
rect 19094 8296 19136 8336
rect 19176 8296 19185 8336
rect 20131 8296 20140 8336
rect 20180 8296 20332 8336
rect 20372 8296 20381 8336
rect 31843 8296 31852 8336
rect 31892 8296 33484 8336
rect 33524 8296 33533 8336
rect 33919 8296 33928 8336
rect 33968 8296 34010 8336
rect 34050 8296 34092 8336
rect 34132 8296 34174 8336
rect 34214 8296 34256 8336
rect 34296 8296 34305 8336
rect 49039 8296 49048 8336
rect 49088 8296 49130 8336
rect 49170 8296 49212 8336
rect 49252 8296 49294 8336
rect 49334 8296 49376 8336
rect 49416 8296 49425 8336
rect 10060 8212 19564 8252
rect 19604 8212 19613 8252
rect 33571 8212 33580 8252
rect 33620 8212 39340 8252
rect 39380 8212 39389 8252
rect 32803 8128 32812 8168
rect 32852 8128 37420 8168
rect 37460 8128 37469 8168
rect 35395 8044 35404 8084
rect 35444 8044 39436 8084
rect 39476 8044 39485 8084
rect 259 7960 268 8000
rect 308 7960 28396 8000
rect 28436 7960 28445 8000
rect 33187 7960 33196 8000
rect 33236 7960 39724 8000
rect 39764 7960 39773 8000
rect 10051 7876 10060 7916
rect 10100 7876 16684 7916
rect 16724 7876 16733 7916
rect 21667 7792 21676 7832
rect 21716 7792 38860 7832
rect 38900 7792 38909 7832
rect 17635 7708 17644 7748
rect 17684 7708 21196 7748
rect 21236 7708 21245 7748
rect 21763 7708 21772 7748
rect 21812 7708 39532 7748
rect 39572 7708 39581 7748
rect 4919 7540 4928 7580
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 5296 7540 5305 7580
rect 20039 7540 20048 7580
rect 20088 7540 20130 7580
rect 20170 7540 20212 7580
rect 20252 7540 20294 7580
rect 20334 7540 20376 7580
rect 20416 7540 20425 7580
rect 25132 7540 29836 7580
rect 29876 7540 29885 7580
rect 35159 7540 35168 7580
rect 35208 7540 35250 7580
rect 35290 7540 35332 7580
rect 35372 7540 35414 7580
rect 35454 7540 35496 7580
rect 35536 7540 35545 7580
rect 50279 7540 50288 7580
rect 50328 7540 50370 7580
rect 50410 7540 50452 7580
rect 50492 7540 50534 7580
rect 50574 7540 50616 7580
rect 50656 7540 50665 7580
rect 25132 7496 25172 7540
rect 19651 7456 19660 7496
rect 19700 7456 25172 7496
rect 28483 7456 28492 7496
rect 28532 7456 30028 7496
rect 30068 7456 30077 7496
rect 34915 7372 34924 7412
rect 34964 7372 38956 7412
rect 38996 7372 39005 7412
rect 38275 7204 38284 7244
rect 38324 7204 39148 7244
rect 39188 7204 39197 7244
rect 37219 7120 37228 7160
rect 37268 7120 39244 7160
rect 39284 7120 39293 7160
rect 38947 7036 38956 7076
rect 38996 7036 39340 7076
rect 39380 7036 39389 7076
rect 3679 6784 3688 6824
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 4056 6784 4065 6824
rect 18799 6784 18808 6824
rect 18848 6784 18890 6824
rect 18930 6784 18972 6824
rect 19012 6784 19054 6824
rect 19094 6784 19136 6824
rect 19176 6784 19185 6824
rect 33919 6784 33928 6824
rect 33968 6784 34010 6824
rect 34050 6784 34092 6824
rect 34132 6784 34174 6824
rect 34214 6784 34256 6824
rect 34296 6784 34305 6824
rect 49039 6784 49048 6824
rect 49088 6784 49130 6824
rect 49170 6784 49212 6824
rect 49252 6784 49294 6824
rect 49334 6784 49376 6824
rect 49416 6784 49425 6824
rect 23395 6532 23404 6572
rect 23444 6532 25708 6572
rect 25748 6532 25757 6572
rect 34723 6196 34732 6236
rect 34772 6196 35116 6236
rect 35156 6196 35165 6236
rect 4919 6028 4928 6068
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 5296 6028 5305 6068
rect 20039 6028 20048 6068
rect 20088 6028 20130 6068
rect 20170 6028 20212 6068
rect 20252 6028 20294 6068
rect 20334 6028 20376 6068
rect 20416 6028 20425 6068
rect 23107 6028 23116 6068
rect 23156 6028 23788 6068
rect 23828 6028 23837 6068
rect 35159 6028 35168 6068
rect 35208 6028 35250 6068
rect 35290 6028 35332 6068
rect 35372 6028 35414 6068
rect 35454 6028 35496 6068
rect 35536 6028 35545 6068
rect 50279 6028 50288 6068
rect 50328 6028 50370 6068
rect 50410 6028 50452 6068
rect 50492 6028 50534 6068
rect 50574 6028 50616 6068
rect 50656 6028 50665 6068
rect 31555 5860 31564 5900
rect 31604 5860 38092 5900
rect 38132 5860 38141 5900
rect 3679 5272 3688 5312
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 4056 5272 4065 5312
rect 18799 5272 18808 5312
rect 18848 5272 18890 5312
rect 18930 5272 18972 5312
rect 19012 5272 19054 5312
rect 19094 5272 19136 5312
rect 19176 5272 19185 5312
rect 33919 5272 33928 5312
rect 33968 5272 34010 5312
rect 34050 5272 34092 5312
rect 34132 5272 34174 5312
rect 34214 5272 34256 5312
rect 34296 5272 34305 5312
rect 49039 5272 49048 5312
rect 49088 5272 49130 5312
rect 49170 5272 49212 5312
rect 49252 5272 49294 5312
rect 49334 5272 49376 5312
rect 49416 5272 49425 5312
rect 4919 4516 4928 4556
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 5296 4516 5305 4556
rect 20039 4516 20048 4556
rect 20088 4516 20130 4556
rect 20170 4516 20212 4556
rect 20252 4516 20294 4556
rect 20334 4516 20376 4556
rect 20416 4516 20425 4556
rect 35159 4516 35168 4556
rect 35208 4516 35250 4556
rect 35290 4516 35332 4556
rect 35372 4516 35414 4556
rect 35454 4516 35496 4556
rect 35536 4516 35545 4556
rect 50279 4516 50288 4556
rect 50328 4516 50370 4556
rect 50410 4516 50452 4556
rect 50492 4516 50534 4556
rect 50574 4516 50616 4556
rect 50656 4516 50665 4556
rect 931 4096 940 4136
rect 980 4096 25996 4136
rect 26036 4096 26045 4136
rect 3679 3760 3688 3800
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 4056 3760 4065 3800
rect 18799 3760 18808 3800
rect 18848 3760 18890 3800
rect 18930 3760 18972 3800
rect 19012 3760 19054 3800
rect 19094 3760 19136 3800
rect 19176 3760 19185 3800
rect 33919 3760 33928 3800
rect 33968 3760 34010 3800
rect 34050 3760 34092 3800
rect 34132 3760 34174 3800
rect 34214 3760 34256 3800
rect 34296 3760 34305 3800
rect 49039 3760 49048 3800
rect 49088 3760 49130 3800
rect 49170 3760 49212 3800
rect 49252 3760 49294 3800
rect 49334 3760 49376 3800
rect 49416 3760 49425 3800
rect 1411 3424 1420 3464
rect 1460 3424 28300 3464
rect 28340 3424 28349 3464
rect 4919 3004 4928 3044
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 5296 3004 5305 3044
rect 20039 3004 20048 3044
rect 20088 3004 20130 3044
rect 20170 3004 20212 3044
rect 20252 3004 20294 3044
rect 20334 3004 20376 3044
rect 20416 3004 20425 3044
rect 35159 3004 35168 3044
rect 35208 3004 35250 3044
rect 35290 3004 35332 3044
rect 35372 3004 35414 3044
rect 35454 3004 35496 3044
rect 35536 3004 35545 3044
rect 50279 3004 50288 3044
rect 50328 3004 50370 3044
rect 50410 3004 50452 3044
rect 50492 3004 50534 3044
rect 50574 3004 50616 3044
rect 50656 3004 50665 3044
rect 3679 2248 3688 2288
rect 3728 2248 3770 2288
rect 3810 2248 3852 2288
rect 3892 2248 3934 2288
rect 3974 2248 4016 2288
rect 4056 2248 4065 2288
rect 18799 2248 18808 2288
rect 18848 2248 18890 2288
rect 18930 2248 18972 2288
rect 19012 2248 19054 2288
rect 19094 2248 19136 2288
rect 19176 2248 19185 2288
rect 33919 2248 33928 2288
rect 33968 2248 34010 2288
rect 34050 2248 34092 2288
rect 34132 2248 34174 2288
rect 34214 2248 34256 2288
rect 34296 2248 34305 2288
rect 49039 2248 49048 2288
rect 49088 2248 49130 2288
rect 49170 2248 49212 2288
rect 49252 2248 49294 2288
rect 49334 2248 49376 2288
rect 49416 2248 49425 2288
rect 4919 1492 4928 1532
rect 4968 1492 5010 1532
rect 5050 1492 5092 1532
rect 5132 1492 5174 1532
rect 5214 1492 5256 1532
rect 5296 1492 5305 1532
rect 20039 1492 20048 1532
rect 20088 1492 20130 1532
rect 20170 1492 20212 1532
rect 20252 1492 20294 1532
rect 20334 1492 20376 1532
rect 20416 1492 20425 1532
rect 35159 1492 35168 1532
rect 35208 1492 35250 1532
rect 35290 1492 35332 1532
rect 35372 1492 35414 1532
rect 35454 1492 35496 1532
rect 35536 1492 35545 1532
rect 50279 1492 50288 1532
rect 50328 1492 50370 1532
rect 50410 1492 50452 1532
rect 50492 1492 50534 1532
rect 50574 1492 50616 1532
rect 50656 1492 50665 1532
rect 34051 64 34060 104
rect 34100 64 34348 104
rect 34388 64 34397 104
<< via4 >>
rect 3688 9808 3728 9848
rect 3770 9808 3810 9848
rect 3852 9808 3892 9848
rect 3934 9808 3974 9848
rect 4016 9808 4056 9848
rect 18808 9808 18848 9848
rect 18890 9808 18930 9848
rect 18972 9808 19012 9848
rect 19054 9808 19094 9848
rect 19136 9808 19176 9848
rect 33928 9808 33968 9848
rect 34010 9808 34050 9848
rect 34092 9808 34132 9848
rect 34174 9808 34214 9848
rect 34256 9808 34296 9848
rect 49048 9808 49088 9848
rect 49130 9808 49170 9848
rect 49212 9808 49252 9848
rect 49294 9808 49334 9848
rect 49376 9808 49416 9848
rect 4928 9052 4968 9092
rect 5010 9052 5050 9092
rect 5092 9052 5132 9092
rect 5174 9052 5214 9092
rect 5256 9052 5296 9092
rect 20048 9052 20088 9092
rect 20130 9052 20170 9092
rect 20212 9052 20252 9092
rect 20294 9052 20334 9092
rect 20376 9052 20416 9092
rect 35168 9052 35208 9092
rect 35250 9052 35290 9092
rect 35332 9052 35372 9092
rect 35414 9052 35454 9092
rect 35496 9052 35536 9092
rect 50288 9052 50328 9092
rect 50370 9052 50410 9092
rect 50452 9052 50492 9092
rect 50534 9052 50574 9092
rect 50616 9052 50656 9092
rect 3688 8296 3728 8336
rect 3770 8296 3810 8336
rect 3852 8296 3892 8336
rect 3934 8296 3974 8336
rect 4016 8296 4056 8336
rect 18808 8296 18848 8336
rect 18890 8296 18930 8336
rect 18972 8296 19012 8336
rect 19054 8296 19094 8336
rect 19136 8296 19176 8336
rect 33928 8296 33968 8336
rect 34010 8296 34050 8336
rect 34092 8296 34132 8336
rect 34174 8296 34214 8336
rect 34256 8296 34296 8336
rect 49048 8296 49088 8336
rect 49130 8296 49170 8336
rect 49212 8296 49252 8336
rect 49294 8296 49334 8336
rect 49376 8296 49416 8336
rect 4928 7540 4968 7580
rect 5010 7540 5050 7580
rect 5092 7540 5132 7580
rect 5174 7540 5214 7580
rect 5256 7540 5296 7580
rect 20048 7540 20088 7580
rect 20130 7540 20170 7580
rect 20212 7540 20252 7580
rect 20294 7540 20334 7580
rect 20376 7540 20416 7580
rect 35168 7540 35208 7580
rect 35250 7540 35290 7580
rect 35332 7540 35372 7580
rect 35414 7540 35454 7580
rect 35496 7540 35536 7580
rect 50288 7540 50328 7580
rect 50370 7540 50410 7580
rect 50452 7540 50492 7580
rect 50534 7540 50574 7580
rect 50616 7540 50656 7580
rect 3688 6784 3728 6824
rect 3770 6784 3810 6824
rect 3852 6784 3892 6824
rect 3934 6784 3974 6824
rect 4016 6784 4056 6824
rect 18808 6784 18848 6824
rect 18890 6784 18930 6824
rect 18972 6784 19012 6824
rect 19054 6784 19094 6824
rect 19136 6784 19176 6824
rect 33928 6784 33968 6824
rect 34010 6784 34050 6824
rect 34092 6784 34132 6824
rect 34174 6784 34214 6824
rect 34256 6784 34296 6824
rect 49048 6784 49088 6824
rect 49130 6784 49170 6824
rect 49212 6784 49252 6824
rect 49294 6784 49334 6824
rect 49376 6784 49416 6824
rect 4928 6028 4968 6068
rect 5010 6028 5050 6068
rect 5092 6028 5132 6068
rect 5174 6028 5214 6068
rect 5256 6028 5296 6068
rect 20048 6028 20088 6068
rect 20130 6028 20170 6068
rect 20212 6028 20252 6068
rect 20294 6028 20334 6068
rect 20376 6028 20416 6068
rect 35168 6028 35208 6068
rect 35250 6028 35290 6068
rect 35332 6028 35372 6068
rect 35414 6028 35454 6068
rect 35496 6028 35536 6068
rect 50288 6028 50328 6068
rect 50370 6028 50410 6068
rect 50452 6028 50492 6068
rect 50534 6028 50574 6068
rect 50616 6028 50656 6068
rect 3688 5272 3728 5312
rect 3770 5272 3810 5312
rect 3852 5272 3892 5312
rect 3934 5272 3974 5312
rect 4016 5272 4056 5312
rect 18808 5272 18848 5312
rect 18890 5272 18930 5312
rect 18972 5272 19012 5312
rect 19054 5272 19094 5312
rect 19136 5272 19176 5312
rect 33928 5272 33968 5312
rect 34010 5272 34050 5312
rect 34092 5272 34132 5312
rect 34174 5272 34214 5312
rect 34256 5272 34296 5312
rect 49048 5272 49088 5312
rect 49130 5272 49170 5312
rect 49212 5272 49252 5312
rect 49294 5272 49334 5312
rect 49376 5272 49416 5312
rect 4928 4516 4968 4556
rect 5010 4516 5050 4556
rect 5092 4516 5132 4556
rect 5174 4516 5214 4556
rect 5256 4516 5296 4556
rect 20048 4516 20088 4556
rect 20130 4516 20170 4556
rect 20212 4516 20252 4556
rect 20294 4516 20334 4556
rect 20376 4516 20416 4556
rect 35168 4516 35208 4556
rect 35250 4516 35290 4556
rect 35332 4516 35372 4556
rect 35414 4516 35454 4556
rect 35496 4516 35536 4556
rect 50288 4516 50328 4556
rect 50370 4516 50410 4556
rect 50452 4516 50492 4556
rect 50534 4516 50574 4556
rect 50616 4516 50656 4556
rect 3688 3760 3728 3800
rect 3770 3760 3810 3800
rect 3852 3760 3892 3800
rect 3934 3760 3974 3800
rect 4016 3760 4056 3800
rect 18808 3760 18848 3800
rect 18890 3760 18930 3800
rect 18972 3760 19012 3800
rect 19054 3760 19094 3800
rect 19136 3760 19176 3800
rect 33928 3760 33968 3800
rect 34010 3760 34050 3800
rect 34092 3760 34132 3800
rect 34174 3760 34214 3800
rect 34256 3760 34296 3800
rect 49048 3760 49088 3800
rect 49130 3760 49170 3800
rect 49212 3760 49252 3800
rect 49294 3760 49334 3800
rect 49376 3760 49416 3800
rect 4928 3004 4968 3044
rect 5010 3004 5050 3044
rect 5092 3004 5132 3044
rect 5174 3004 5214 3044
rect 5256 3004 5296 3044
rect 20048 3004 20088 3044
rect 20130 3004 20170 3044
rect 20212 3004 20252 3044
rect 20294 3004 20334 3044
rect 20376 3004 20416 3044
rect 35168 3004 35208 3044
rect 35250 3004 35290 3044
rect 35332 3004 35372 3044
rect 35414 3004 35454 3044
rect 35496 3004 35536 3044
rect 50288 3004 50328 3044
rect 50370 3004 50410 3044
rect 50452 3004 50492 3044
rect 50534 3004 50574 3044
rect 50616 3004 50656 3044
rect 3688 2248 3728 2288
rect 3770 2248 3810 2288
rect 3852 2248 3892 2288
rect 3934 2248 3974 2288
rect 4016 2248 4056 2288
rect 18808 2248 18848 2288
rect 18890 2248 18930 2288
rect 18972 2248 19012 2288
rect 19054 2248 19094 2288
rect 19136 2248 19176 2288
rect 33928 2248 33968 2288
rect 34010 2248 34050 2288
rect 34092 2248 34132 2288
rect 34174 2248 34214 2288
rect 34256 2248 34296 2288
rect 49048 2248 49088 2288
rect 49130 2248 49170 2288
rect 49212 2248 49252 2288
rect 49294 2248 49334 2288
rect 49376 2248 49416 2288
rect 4928 1492 4968 1532
rect 5010 1492 5050 1532
rect 5092 1492 5132 1532
rect 5174 1492 5214 1532
rect 5256 1492 5296 1532
rect 20048 1492 20088 1532
rect 20130 1492 20170 1532
rect 20212 1492 20252 1532
rect 20294 1492 20334 1532
rect 20376 1492 20416 1532
rect 35168 1492 35208 1532
rect 35250 1492 35290 1532
rect 35332 1492 35372 1532
rect 35414 1492 35454 1532
rect 35496 1492 35536 1532
rect 50288 1492 50328 1532
rect 50370 1492 50410 1532
rect 50452 1492 50492 1532
rect 50534 1492 50574 1532
rect 50616 1492 50656 1532
<< metal5 >>
rect 3652 9848 4092 11844
rect 3652 9808 3688 9848
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 4056 9808 4092 9848
rect 3652 8336 4092 9808
rect 3652 8296 3688 8336
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 4056 8296 4092 8336
rect 3652 6824 4092 8296
rect 3652 6784 3688 6824
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 4056 6784 4092 6824
rect 3652 5312 4092 6784
rect 3652 5272 3688 5312
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 4056 5272 4092 5312
rect 3652 3800 4092 5272
rect 3652 3760 3688 3800
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 4056 3760 4092 3800
rect 3652 2288 4092 3760
rect 3652 2248 3688 2288
rect 3728 2248 3770 2288
rect 3810 2248 3852 2288
rect 3892 2248 3934 2288
rect 3974 2248 4016 2288
rect 4056 2248 4092 2288
rect 3652 0 4092 2248
rect 4892 9092 5332 11844
rect 4892 9052 4928 9092
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 5296 9052 5332 9092
rect 4892 7580 5332 9052
rect 4892 7540 4928 7580
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 5296 7540 5332 7580
rect 4892 6068 5332 7540
rect 4892 6028 4928 6068
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 5296 6028 5332 6068
rect 4892 4556 5332 6028
rect 4892 4516 4928 4556
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 5296 4516 5332 4556
rect 4892 3044 5332 4516
rect 4892 3004 4928 3044
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 5296 3004 5332 3044
rect 4892 1532 5332 3004
rect 4892 1492 4928 1532
rect 4968 1492 5010 1532
rect 5050 1492 5092 1532
rect 5132 1492 5174 1532
rect 5214 1492 5256 1532
rect 5296 1492 5332 1532
rect 4892 0 5332 1492
rect 18772 9848 19212 11844
rect 18772 9808 18808 9848
rect 18848 9808 18890 9848
rect 18930 9808 18972 9848
rect 19012 9808 19054 9848
rect 19094 9808 19136 9848
rect 19176 9808 19212 9848
rect 18772 8336 19212 9808
rect 18772 8296 18808 8336
rect 18848 8296 18890 8336
rect 18930 8296 18972 8336
rect 19012 8296 19054 8336
rect 19094 8296 19136 8336
rect 19176 8296 19212 8336
rect 18772 6824 19212 8296
rect 18772 6784 18808 6824
rect 18848 6784 18890 6824
rect 18930 6784 18972 6824
rect 19012 6784 19054 6824
rect 19094 6784 19136 6824
rect 19176 6784 19212 6824
rect 18772 5312 19212 6784
rect 18772 5272 18808 5312
rect 18848 5272 18890 5312
rect 18930 5272 18972 5312
rect 19012 5272 19054 5312
rect 19094 5272 19136 5312
rect 19176 5272 19212 5312
rect 18772 3800 19212 5272
rect 18772 3760 18808 3800
rect 18848 3760 18890 3800
rect 18930 3760 18972 3800
rect 19012 3760 19054 3800
rect 19094 3760 19136 3800
rect 19176 3760 19212 3800
rect 18772 2288 19212 3760
rect 18772 2248 18808 2288
rect 18848 2248 18890 2288
rect 18930 2248 18972 2288
rect 19012 2248 19054 2288
rect 19094 2248 19136 2288
rect 19176 2248 19212 2288
rect 18772 0 19212 2248
rect 20012 9092 20452 11844
rect 20012 9052 20048 9092
rect 20088 9052 20130 9092
rect 20170 9052 20212 9092
rect 20252 9052 20294 9092
rect 20334 9052 20376 9092
rect 20416 9052 20452 9092
rect 20012 7580 20452 9052
rect 20012 7540 20048 7580
rect 20088 7540 20130 7580
rect 20170 7540 20212 7580
rect 20252 7540 20294 7580
rect 20334 7540 20376 7580
rect 20416 7540 20452 7580
rect 20012 6068 20452 7540
rect 20012 6028 20048 6068
rect 20088 6028 20130 6068
rect 20170 6028 20212 6068
rect 20252 6028 20294 6068
rect 20334 6028 20376 6068
rect 20416 6028 20452 6068
rect 20012 4556 20452 6028
rect 20012 4516 20048 4556
rect 20088 4516 20130 4556
rect 20170 4516 20212 4556
rect 20252 4516 20294 4556
rect 20334 4516 20376 4556
rect 20416 4516 20452 4556
rect 20012 3044 20452 4516
rect 20012 3004 20048 3044
rect 20088 3004 20130 3044
rect 20170 3004 20212 3044
rect 20252 3004 20294 3044
rect 20334 3004 20376 3044
rect 20416 3004 20452 3044
rect 20012 1532 20452 3004
rect 20012 1492 20048 1532
rect 20088 1492 20130 1532
rect 20170 1492 20212 1532
rect 20252 1492 20294 1532
rect 20334 1492 20376 1532
rect 20416 1492 20452 1532
rect 20012 0 20452 1492
rect 33892 9848 34332 11844
rect 33892 9808 33928 9848
rect 33968 9808 34010 9848
rect 34050 9808 34092 9848
rect 34132 9808 34174 9848
rect 34214 9808 34256 9848
rect 34296 9808 34332 9848
rect 33892 8336 34332 9808
rect 33892 8296 33928 8336
rect 33968 8296 34010 8336
rect 34050 8296 34092 8336
rect 34132 8296 34174 8336
rect 34214 8296 34256 8336
rect 34296 8296 34332 8336
rect 33892 6824 34332 8296
rect 33892 6784 33928 6824
rect 33968 6784 34010 6824
rect 34050 6784 34092 6824
rect 34132 6784 34174 6824
rect 34214 6784 34256 6824
rect 34296 6784 34332 6824
rect 33892 5312 34332 6784
rect 33892 5272 33928 5312
rect 33968 5272 34010 5312
rect 34050 5272 34092 5312
rect 34132 5272 34174 5312
rect 34214 5272 34256 5312
rect 34296 5272 34332 5312
rect 33892 3800 34332 5272
rect 33892 3760 33928 3800
rect 33968 3760 34010 3800
rect 34050 3760 34092 3800
rect 34132 3760 34174 3800
rect 34214 3760 34256 3800
rect 34296 3760 34332 3800
rect 33892 2288 34332 3760
rect 33892 2248 33928 2288
rect 33968 2248 34010 2288
rect 34050 2248 34092 2288
rect 34132 2248 34174 2288
rect 34214 2248 34256 2288
rect 34296 2248 34332 2288
rect 33892 0 34332 2248
rect 35132 9092 35572 11844
rect 35132 9052 35168 9092
rect 35208 9052 35250 9092
rect 35290 9052 35332 9092
rect 35372 9052 35414 9092
rect 35454 9052 35496 9092
rect 35536 9052 35572 9092
rect 35132 7580 35572 9052
rect 35132 7540 35168 7580
rect 35208 7540 35250 7580
rect 35290 7540 35332 7580
rect 35372 7540 35414 7580
rect 35454 7540 35496 7580
rect 35536 7540 35572 7580
rect 35132 6068 35572 7540
rect 35132 6028 35168 6068
rect 35208 6028 35250 6068
rect 35290 6028 35332 6068
rect 35372 6028 35414 6068
rect 35454 6028 35496 6068
rect 35536 6028 35572 6068
rect 35132 4556 35572 6028
rect 35132 4516 35168 4556
rect 35208 4516 35250 4556
rect 35290 4516 35332 4556
rect 35372 4516 35414 4556
rect 35454 4516 35496 4556
rect 35536 4516 35572 4556
rect 35132 3044 35572 4516
rect 35132 3004 35168 3044
rect 35208 3004 35250 3044
rect 35290 3004 35332 3044
rect 35372 3004 35414 3044
rect 35454 3004 35496 3044
rect 35536 3004 35572 3044
rect 35132 1532 35572 3004
rect 35132 1492 35168 1532
rect 35208 1492 35250 1532
rect 35290 1492 35332 1532
rect 35372 1492 35414 1532
rect 35454 1492 35496 1532
rect 35536 1492 35572 1532
rect 35132 0 35572 1492
rect 49012 9848 49452 11844
rect 49012 9808 49048 9848
rect 49088 9808 49130 9848
rect 49170 9808 49212 9848
rect 49252 9808 49294 9848
rect 49334 9808 49376 9848
rect 49416 9808 49452 9848
rect 49012 8336 49452 9808
rect 49012 8296 49048 8336
rect 49088 8296 49130 8336
rect 49170 8296 49212 8336
rect 49252 8296 49294 8336
rect 49334 8296 49376 8336
rect 49416 8296 49452 8336
rect 49012 6824 49452 8296
rect 49012 6784 49048 6824
rect 49088 6784 49130 6824
rect 49170 6784 49212 6824
rect 49252 6784 49294 6824
rect 49334 6784 49376 6824
rect 49416 6784 49452 6824
rect 49012 5312 49452 6784
rect 49012 5272 49048 5312
rect 49088 5272 49130 5312
rect 49170 5272 49212 5312
rect 49252 5272 49294 5312
rect 49334 5272 49376 5312
rect 49416 5272 49452 5312
rect 49012 3800 49452 5272
rect 49012 3760 49048 3800
rect 49088 3760 49130 3800
rect 49170 3760 49212 3800
rect 49252 3760 49294 3800
rect 49334 3760 49376 3800
rect 49416 3760 49452 3800
rect 49012 2288 49452 3760
rect 49012 2248 49048 2288
rect 49088 2248 49130 2288
rect 49170 2248 49212 2288
rect 49252 2248 49294 2288
rect 49334 2248 49376 2288
rect 49416 2248 49452 2288
rect 49012 0 49452 2248
rect 50252 9092 50692 11844
rect 50252 9052 50288 9092
rect 50328 9052 50370 9092
rect 50410 9052 50452 9092
rect 50492 9052 50534 9092
rect 50574 9052 50616 9092
rect 50656 9052 50692 9092
rect 50252 7580 50692 9052
rect 50252 7540 50288 7580
rect 50328 7540 50370 7580
rect 50410 7540 50452 7580
rect 50492 7540 50534 7580
rect 50574 7540 50616 7580
rect 50656 7540 50692 7580
rect 50252 6068 50692 7540
rect 50252 6028 50288 6068
rect 50328 6028 50370 6068
rect 50410 6028 50452 6068
rect 50492 6028 50534 6068
rect 50574 6028 50616 6068
rect 50656 6028 50692 6068
rect 50252 4556 50692 6028
rect 50252 4516 50288 4556
rect 50328 4516 50370 4556
rect 50410 4516 50452 4556
rect 50492 4516 50534 4556
rect 50574 4516 50616 4556
rect 50656 4516 50692 4556
rect 50252 3044 50692 4516
rect 50252 3004 50288 3044
rect 50328 3004 50370 3044
rect 50410 3004 50452 3044
rect 50492 3004 50534 3044
rect 50574 3004 50616 3044
rect 50656 3004 50692 3044
rect 50252 1532 50692 3004
rect 50252 1492 50288 1532
rect 50328 1492 50370 1532
rect 50410 1492 50452 1532
rect 50492 1492 50534 1532
rect 50574 1492 50616 1532
rect 50656 1492 50692 1532
rect 50252 0 50692 1492
use sg13g2_buf_1  _000_
timestamp 1676381911
transform 1 0 20544 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _001_
timestamp 1676381911
transform 1 0 22464 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _002_
timestamp 1676381911
transform 1 0 23232 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _003_
timestamp 1676381911
transform 1 0 22848 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _004_
timestamp 1676381911
transform 1 0 21600 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _005_
timestamp 1676381911
transform 1 0 25536 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _006_
timestamp 1676381911
transform 1 0 24768 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _007_
timestamp 1676381911
transform 1 0 24000 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _008_
timestamp 1676381911
transform 1 0 25152 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _009_
timestamp 1676381911
transform 1 0 21984 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _010_
timestamp 1676381911
transform 1 0 24768 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _011_
timestamp 1676381911
transform 1 0 24384 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _012_
timestamp 1676381911
transform 1 0 25152 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _013_
timestamp 1676381911
transform 1 0 24192 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _014_
timestamp 1676381911
transform 1 0 21696 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _015_
timestamp 1676381911
transform 1 0 23040 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _016_
timestamp 1676381911
transform 1 0 25152 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _017_
timestamp 1676381911
transform 1 0 28224 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _018_
timestamp 1676381911
transform 1 0 25920 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _019_
timestamp 1676381911
transform 1 0 27552 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _020_
timestamp 1676381911
transform 1 0 27360 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _021_
timestamp 1676381911
transform 1 0 26976 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _022_
timestamp 1676381911
transform 1 0 28704 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _023_
timestamp 1676381911
transform 1 0 26688 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _024_
timestamp 1676381911
transform 1 0 28992 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _025_
timestamp 1676381911
transform 1 0 28608 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _026_
timestamp 1676381911
transform 1 0 28320 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _027_
timestamp 1676381911
transform 1 0 28224 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _028_
timestamp 1676381911
transform 1 0 27840 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _029_
timestamp 1676381911
transform 1 0 27072 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _030_
timestamp 1676381911
transform 1 0 27456 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _031_
timestamp 1676381911
transform 1 0 29376 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _032_
timestamp 1676381911
transform 1 0 24960 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _033_
timestamp 1676381911
transform 1 0 23520 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _034_
timestamp 1676381911
transform 1 0 25536 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _035_
timestamp 1676381911
transform 1 0 23136 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _036_
timestamp 1676381911
transform 1 0 29760 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _037_
timestamp 1676381911
transform 1 0 31584 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _038_
timestamp 1676381911
transform 1 0 31680 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _039_
timestamp 1676381911
transform 1 0 32352 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _040_
timestamp 1676381911
transform 1 0 33024 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _041_
timestamp 1676381911
transform 1 0 34752 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _042_
timestamp 1676381911
transform 1 0 37344 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _043_
timestamp 1676381911
transform 1 0 38016 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _044_
timestamp 1676381911
transform 1 0 37824 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _045_
timestamp 1676381911
transform 1 0 36288 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _046_
timestamp 1676381911
transform 1 0 36672 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _047_
timestamp 1676381911
transform 1 0 39552 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _048_
timestamp 1676381911
transform 1 0 42240 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _049_
timestamp 1676381911
transform 1 0 46368 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _050_
timestamp 1676381911
transform 1 0 49248 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _051_
timestamp 1676381911
transform 1 0 49152 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _052_
timestamp 1676381911
transform -1 0 10944 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _053_
timestamp 1676381911
transform -1 0 8544 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _054_
timestamp 1676381911
transform -1 0 4704 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _055_
timestamp 1676381911
transform 1 0 3168 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _056_
timestamp 1676381911
transform -1 0 16032 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _057_
timestamp 1676381911
transform -1 0 15360 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _058_
timestamp 1676381911
transform -1 0 14112 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _059_
timestamp 1676381911
transform -1 0 12288 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _060_
timestamp 1676381911
transform -1 0 10560 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _061_
timestamp 1676381911
transform -1 0 8160 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _062_
timestamp 1676381911
transform 1 0 6048 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _063_
timestamp 1676381911
transform 1 0 5184 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _064_
timestamp 1676381911
transform -1 0 16416 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _065_
timestamp 1676381911
transform -1 0 15648 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _066_
timestamp 1676381911
transform -1 0 14976 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _067_
timestamp 1676381911
transform -1 0 13728 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _068_
timestamp 1676381911
transform -1 0 12768 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _069_
timestamp 1676381911
transform -1 0 12096 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _070_
timestamp 1676381911
transform -1 0 11616 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _071_
timestamp 1676381911
transform -1 0 11232 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _072_
timestamp 1676381911
transform -1 0 24000 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _073_
timestamp 1676381911
transform -1 0 23424 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _074_
timestamp 1676381911
transform -1 0 22848 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _075_
timestamp 1676381911
transform -1 0 22464 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _076_
timestamp 1676381911
transform -1 0 21984 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _077_
timestamp 1676381911
transform -1 0 21120 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _078_
timestamp 1676381911
transform -1 0 20640 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _079_
timestamp 1676381911
transform -1 0 19776 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _080_
timestamp 1676381911
transform -1 0 18720 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _081_
timestamp 1676381911
transform -1 0 17952 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _082_
timestamp 1676381911
transform -1 0 17184 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _083_
timestamp 1676381911
transform -1 0 17280 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _084_
timestamp 1676381911
transform -1 0 16800 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _085_
timestamp 1676381911
transform -1 0 17568 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _086_
timestamp 1676381911
transform -1 0 18336 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _087_
timestamp 1676381911
transform -1 0 19392 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _088_
timestamp 1676381911
transform -1 0 31584 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _089_
timestamp 1676381911
transform -1 0 33120 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _090_
timestamp 1676381911
transform -1 0 33504 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _091_
timestamp 1676381911
transform -1 0 33888 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _092_
timestamp 1676381911
transform -1 0 35040 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _093_
timestamp 1676381911
transform -1 0 35424 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _094_
timestamp 1676381911
transform -1 0 36192 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _095_
timestamp 1676381911
transform -1 0 37824 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _096_
timestamp 1676381911
transform -1 0 38976 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _097_
timestamp 1676381911
transform -1 0 39744 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _098_
timestamp 1676381911
transform -1 0 40128 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _099_
timestamp 1676381911
transform -1 0 39264 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _100_
timestamp 1676381911
transform -1 0 39360 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _101_
timestamp 1676381911
transform -1 0 38592 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _102_
timestamp 1676381911
transform -1 0 37440 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _103_
timestamp 1676381911
transform -1 0 35808 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _104_
timestamp 1676381911
transform 1 0 26688 0 -1 6048
box -48 -56 432 834
use sg13g2_decap_8  FILLER_0_0
timestamp 1679581782
transform 1 0 1152 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_7
timestamp 1679581782
transform 1 0 1824 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_14
timestamp 1679581782
transform 1 0 2496 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_21
timestamp 1679581782
transform 1 0 3168 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_28
timestamp 1679581782
transform 1 0 3840 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_35
timestamp 1679581782
transform 1 0 4512 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_42
timestamp 1679581782
transform 1 0 5184 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_49
timestamp 1679581782
transform 1 0 5856 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_56
timestamp 1679581782
transform 1 0 6528 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_63
timestamp 1679581782
transform 1 0 7200 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_70
timestamp 1679581782
transform 1 0 7872 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_77
timestamp 1679581782
transform 1 0 8544 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_84
timestamp 1679581782
transform 1 0 9216 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_91
timestamp 1679581782
transform 1 0 9888 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_98
timestamp 1679581782
transform 1 0 10560 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_105
timestamp 1679581782
transform 1 0 11232 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_112
timestamp 1679581782
transform 1 0 11904 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_119
timestamp 1679581782
transform 1 0 12576 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_126
timestamp 1679581782
transform 1 0 13248 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_133
timestamp 1679581782
transform 1 0 13920 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_140
timestamp 1679581782
transform 1 0 14592 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_147
timestamp 1679581782
transform 1 0 15264 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_154
timestamp 1679581782
transform 1 0 15936 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_161
timestamp 1679581782
transform 1 0 16608 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_168
timestamp 1679581782
transform 1 0 17280 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_175
timestamp 1679581782
transform 1 0 17952 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_182
timestamp 1679581782
transform 1 0 18624 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_189
timestamp 1679581782
transform 1 0 19296 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_196
timestamp 1679581782
transform 1 0 19968 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_203
timestamp 1679581782
transform 1 0 20640 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_210
timestamp 1679581782
transform 1 0 21312 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_217
timestamp 1679581782
transform 1 0 21984 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_224
timestamp 1679581782
transform 1 0 22656 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_231
timestamp 1679581782
transform 1 0 23328 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_238
timestamp 1679581782
transform 1 0 24000 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_245
timestamp 1679581782
transform 1 0 24672 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_252
timestamp 1679581782
transform 1 0 25344 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_259
timestamp 1679581782
transform 1 0 26016 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_266
timestamp 1679581782
transform 1 0 26688 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_273
timestamp 1679581782
transform 1 0 27360 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_280
timestamp 1679581782
transform 1 0 28032 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_287
timestamp 1679581782
transform 1 0 28704 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_294
timestamp 1679581782
transform 1 0 29376 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_301
timestamp 1679581782
transform 1 0 30048 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_308
timestamp 1679581782
transform 1 0 30720 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_315
timestamp 1679581782
transform 1 0 31392 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_322
timestamp 1679581782
transform 1 0 32064 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_329
timestamp 1679581782
transform 1 0 32736 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_336
timestamp 1679581782
transform 1 0 33408 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_343
timestamp 1679581782
transform 1 0 34080 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_350
timestamp 1679581782
transform 1 0 34752 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_357
timestamp 1679581782
transform 1 0 35424 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_364
timestamp 1679581782
transform 1 0 36096 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_371
timestamp 1679581782
transform 1 0 36768 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_378
timestamp 1679581782
transform 1 0 37440 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_385
timestamp 1679581782
transform 1 0 38112 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_392
timestamp 1679581782
transform 1 0 38784 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_399
timestamp 1679581782
transform 1 0 39456 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_406
timestamp 1679581782
transform 1 0 40128 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_413
timestamp 1679581782
transform 1 0 40800 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_420
timestamp 1679581782
transform 1 0 41472 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_427
timestamp 1679581782
transform 1 0 42144 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_434
timestamp 1679581782
transform 1 0 42816 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_441
timestamp 1679581782
transform 1 0 43488 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_448
timestamp 1679581782
transform 1 0 44160 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_455
timestamp 1679581782
transform 1 0 44832 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_462
timestamp 1679581782
transform 1 0 45504 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_469
timestamp 1679581782
transform 1 0 46176 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_476
timestamp 1679581782
transform 1 0 46848 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_483
timestamp 1679581782
transform 1 0 47520 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_490
timestamp 1679581782
transform 1 0 48192 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_497
timestamp 1679581782
transform 1 0 48864 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_504
timestamp 1679581782
transform 1 0 49536 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_0
timestamp 1679581782
transform 1 0 1152 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_7
timestamp 1679581782
transform 1 0 1824 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_14
timestamp 1679581782
transform 1 0 2496 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_21
timestamp 1679581782
transform 1 0 3168 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_28
timestamp 1679581782
transform 1 0 3840 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_35
timestamp 1679581782
transform 1 0 4512 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_42
timestamp 1679581782
transform 1 0 5184 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_49
timestamp 1679581782
transform 1 0 5856 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_56
timestamp 1679581782
transform 1 0 6528 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_63
timestamp 1679581782
transform 1 0 7200 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_70
timestamp 1679581782
transform 1 0 7872 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_77
timestamp 1679581782
transform 1 0 8544 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_84
timestamp 1679581782
transform 1 0 9216 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_91
timestamp 1679581782
transform 1 0 9888 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_98
timestamp 1679581782
transform 1 0 10560 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_105
timestamp 1679581782
transform 1 0 11232 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_112
timestamp 1679581782
transform 1 0 11904 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_119
timestamp 1679581782
transform 1 0 12576 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_126
timestamp 1679581782
transform 1 0 13248 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_133
timestamp 1679581782
transform 1 0 13920 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_140
timestamp 1679581782
transform 1 0 14592 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_147
timestamp 1679581782
transform 1 0 15264 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_154
timestamp 1679581782
transform 1 0 15936 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_161
timestamp 1679581782
transform 1 0 16608 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_168
timestamp 1679581782
transform 1 0 17280 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_175
timestamp 1679581782
transform 1 0 17952 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_182
timestamp 1679581782
transform 1 0 18624 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_189
timestamp 1679581782
transform 1 0 19296 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_196
timestamp 1679581782
transform 1 0 19968 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_203
timestamp 1679581782
transform 1 0 20640 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_210
timestamp 1679581782
transform 1 0 21312 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_217
timestamp 1679581782
transform 1 0 21984 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_224
timestamp 1679581782
transform 1 0 22656 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_231
timestamp 1679581782
transform 1 0 23328 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_238
timestamp 1679581782
transform 1 0 24000 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_4  FILLER_1_245
timestamp 1679577901
transform 1 0 24672 0 -1 3024
box -48 -56 432 834
use sg13g2_fill_1  FILLER_1_249
timestamp 1677579658
transform 1 0 25056 0 -1 3024
box -48 -56 144 834
use sg13g2_decap_8  FILLER_1_254
timestamp 1679581782
transform 1 0 25536 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_261
timestamp 1679581782
transform 1 0 26208 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_268
timestamp 1679581782
transform 1 0 26880 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_275
timestamp 1679581782
transform 1 0 27552 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_282
timestamp 1679581782
transform 1 0 28224 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_289
timestamp 1679581782
transform 1 0 28896 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_296
timestamp 1679581782
transform 1 0 29568 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_303
timestamp 1679581782
transform 1 0 30240 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_310
timestamp 1679581782
transform 1 0 30912 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_317
timestamp 1679581782
transform 1 0 31584 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_324
timestamp 1679581782
transform 1 0 32256 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_331
timestamp 1679581782
transform 1 0 32928 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_338
timestamp 1679581782
transform 1 0 33600 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_345
timestamp 1679581782
transform 1 0 34272 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_352
timestamp 1679581782
transform 1 0 34944 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_359
timestamp 1679581782
transform 1 0 35616 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_366
timestamp 1679581782
transform 1 0 36288 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_373
timestamp 1679581782
transform 1 0 36960 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_380
timestamp 1679581782
transform 1 0 37632 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_387
timestamp 1679581782
transform 1 0 38304 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_394
timestamp 1679581782
transform 1 0 38976 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_401
timestamp 1679581782
transform 1 0 39648 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_408
timestamp 1679581782
transform 1 0 40320 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_415
timestamp 1679581782
transform 1 0 40992 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_422
timestamp 1679581782
transform 1 0 41664 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_429
timestamp 1679581782
transform 1 0 42336 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_436
timestamp 1679581782
transform 1 0 43008 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_443
timestamp 1679581782
transform 1 0 43680 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_450
timestamp 1679581782
transform 1 0 44352 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_457
timestamp 1679581782
transform 1 0 45024 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_464
timestamp 1679581782
transform 1 0 45696 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_471
timestamp 1679581782
transform 1 0 46368 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_478
timestamp 1679581782
transform 1 0 47040 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_485
timestamp 1679581782
transform 1 0 47712 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_492
timestamp 1679581782
transform 1 0 48384 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_499
timestamp 1679581782
transform 1 0 49056 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_506
timestamp 1679581782
transform 1 0 49728 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_4  FILLER_1_513
timestamp 1679577901
transform 1 0 50400 0 -1 3024
box -48 -56 432 834
use sg13g2_fill_2  FILLER_1_517
timestamp 1677580104
transform 1 0 50784 0 -1 3024
box -48 -56 240 834
use sg13g2_decap_8  FILLER_2_0
timestamp 1679581782
transform 1 0 1152 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_7
timestamp 1679581782
transform 1 0 1824 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_14
timestamp 1679581782
transform 1 0 2496 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_21
timestamp 1679581782
transform 1 0 3168 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_28
timestamp 1679581782
transform 1 0 3840 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_35
timestamp 1679581782
transform 1 0 4512 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_42
timestamp 1679581782
transform 1 0 5184 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_49
timestamp 1679581782
transform 1 0 5856 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_56
timestamp 1679581782
transform 1 0 6528 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_63
timestamp 1679581782
transform 1 0 7200 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_70
timestamp 1679581782
transform 1 0 7872 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_77
timestamp 1679581782
transform 1 0 8544 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_84
timestamp 1679581782
transform 1 0 9216 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_91
timestamp 1679581782
transform 1 0 9888 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_98
timestamp 1679581782
transform 1 0 10560 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_105
timestamp 1679581782
transform 1 0 11232 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_112
timestamp 1679581782
transform 1 0 11904 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_119
timestamp 1679581782
transform 1 0 12576 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_126
timestamp 1679581782
transform 1 0 13248 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_133
timestamp 1679581782
transform 1 0 13920 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_140
timestamp 1679581782
transform 1 0 14592 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_147
timestamp 1679581782
transform 1 0 15264 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_154
timestamp 1679581782
transform 1 0 15936 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_161
timestamp 1679581782
transform 1 0 16608 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_168
timestamp 1679581782
transform 1 0 17280 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_175
timestamp 1679581782
transform 1 0 17952 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_182
timestamp 1679581782
transform 1 0 18624 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_189
timestamp 1679581782
transform 1 0 19296 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_196
timestamp 1679581782
transform 1 0 19968 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_203
timestamp 1679581782
transform 1 0 20640 0 1 3024
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_210
timestamp 1679577901
transform 1 0 21312 0 1 3024
box -48 -56 432 834
use sg13g2_decap_8  FILLER_2_218
timestamp 1679581782
transform 1 0 22080 0 1 3024
box -48 -56 720 834
use sg13g2_fill_2  FILLER_2_225
timestamp 1677580104
transform 1 0 22752 0 1 3024
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_227
timestamp 1677579658
transform 1 0 22944 0 1 3024
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_232
timestamp 1679581782
transform 1 0 23424 0 1 3024
box -48 -56 720 834
use sg13g2_fill_1  FILLER_2_239
timestamp 1677579658
transform 1 0 24096 0 1 3024
box -48 -56 144 834
use sg13g2_fill_2  FILLER_2_244
timestamp 1677580104
transform 1 0 24576 0 1 3024
box -48 -56 240 834
use sg13g2_decap_8  FILLER_2_254
timestamp 1679581782
transform 1 0 25536 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_261
timestamp 1679581782
transform 1 0 26208 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_268
timestamp 1679581782
transform 1 0 26880 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_275
timestamp 1679581782
transform 1 0 27552 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_286
timestamp 1679581782
transform 1 0 28608 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_293
timestamp 1679581782
transform 1 0 29280 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_300
timestamp 1679581782
transform 1 0 29952 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_307
timestamp 1679581782
transform 1 0 30624 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_314
timestamp 1679581782
transform 1 0 31296 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_321
timestamp 1679581782
transform 1 0 31968 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_328
timestamp 1679581782
transform 1 0 32640 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_335
timestamp 1679581782
transform 1 0 33312 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_342
timestamp 1679581782
transform 1 0 33984 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_349
timestamp 1679581782
transform 1 0 34656 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_356
timestamp 1679581782
transform 1 0 35328 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_363
timestamp 1679581782
transform 1 0 36000 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_370
timestamp 1679581782
transform 1 0 36672 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_377
timestamp 1679581782
transform 1 0 37344 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_384
timestamp 1679581782
transform 1 0 38016 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_391
timestamp 1679581782
transform 1 0 38688 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_398
timestamp 1679581782
transform 1 0 39360 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_405
timestamp 1679581782
transform 1 0 40032 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_412
timestamp 1679581782
transform 1 0 40704 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_419
timestamp 1679581782
transform 1 0 41376 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_426
timestamp 1679581782
transform 1 0 42048 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_433
timestamp 1679581782
transform 1 0 42720 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_440
timestamp 1679581782
transform 1 0 43392 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_447
timestamp 1679581782
transform 1 0 44064 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_454
timestamp 1679581782
transform 1 0 44736 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_461
timestamp 1679581782
transform 1 0 45408 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_468
timestamp 1679581782
transform 1 0 46080 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_475
timestamp 1679581782
transform 1 0 46752 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_482
timestamp 1679581782
transform 1 0 47424 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_489
timestamp 1679581782
transform 1 0 48096 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_496
timestamp 1679581782
transform 1 0 48768 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_503
timestamp 1679581782
transform 1 0 49440 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_510
timestamp 1679581782
transform 1 0 50112 0 1 3024
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_517
timestamp 1679577901
transform 1 0 50784 0 1 3024
box -48 -56 432 834
use sg13g2_fill_2  FILLER_2_521
timestamp 1677580104
transform 1 0 51168 0 1 3024
box -48 -56 240 834
use sg13g2_decap_8  FILLER_3_0
timestamp 1679581782
transform 1 0 1152 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_7
timestamp 1679581782
transform 1 0 1824 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_14
timestamp 1679581782
transform 1 0 2496 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_21
timestamp 1679581782
transform 1 0 3168 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_28
timestamp 1679581782
transform 1 0 3840 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_35
timestamp 1679581782
transform 1 0 4512 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_42
timestamp 1679581782
transform 1 0 5184 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_49
timestamp 1679581782
transform 1 0 5856 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_56
timestamp 1679581782
transform 1 0 6528 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_63
timestamp 1679581782
transform 1 0 7200 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_70
timestamp 1679581782
transform 1 0 7872 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_77
timestamp 1679581782
transform 1 0 8544 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_84
timestamp 1679581782
transform 1 0 9216 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_91
timestamp 1679581782
transform 1 0 9888 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_98
timestamp 1679581782
transform 1 0 10560 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_105
timestamp 1679581782
transform 1 0 11232 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_112
timestamp 1679581782
transform 1 0 11904 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_119
timestamp 1679581782
transform 1 0 12576 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_126
timestamp 1679581782
transform 1 0 13248 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_133
timestamp 1679581782
transform 1 0 13920 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_140
timestamp 1679581782
transform 1 0 14592 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_147
timestamp 1679581782
transform 1 0 15264 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_154
timestamp 1679581782
transform 1 0 15936 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_161
timestamp 1679581782
transform 1 0 16608 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_168
timestamp 1679581782
transform 1 0 17280 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_175
timestamp 1679581782
transform 1 0 17952 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_182
timestamp 1679581782
transform 1 0 18624 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_189
timestamp 1679581782
transform 1 0 19296 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_196
timestamp 1679577901
transform 1 0 19968 0 -1 4536
box -48 -56 432 834
use sg13g2_fill_2  FILLER_3_200
timestamp 1677580104
transform 1 0 20352 0 -1 4536
box -48 -56 240 834
use sg13g2_decap_8  FILLER_3_206
timestamp 1679581782
transform 1 0 20928 0 -1 4536
box -48 -56 720 834
use sg13g2_fill_1  FILLER_3_221
timestamp 1677579658
transform 1 0 22368 0 -1 4536
box -48 -56 144 834
use sg13g2_decap_4  FILLER_3_234
timestamp 1679577901
transform 1 0 23616 0 -1 4536
box -48 -56 432 834
use sg13g2_decap_8  FILLER_3_262
timestamp 1679581782
transform 1 0 26304 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_269
timestamp 1679581782
transform 1 0 26976 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_276
timestamp 1679581782
transform 1 0 27648 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_283
timestamp 1679581782
transform 1 0 28320 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_290
timestamp 1679581782
transform 1 0 28992 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_297
timestamp 1679581782
transform 1 0 29664 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_304
timestamp 1679581782
transform 1 0 30336 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_311
timestamp 1679581782
transform 1 0 31008 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_318
timestamp 1679581782
transform 1 0 31680 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_325
timestamp 1679581782
transform 1 0 32352 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_332
timestamp 1679581782
transform 1 0 33024 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_339
timestamp 1679581782
transform 1 0 33696 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_346
timestamp 1679581782
transform 1 0 34368 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_353
timestamp 1679581782
transform 1 0 35040 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_360
timestamp 1679581782
transform 1 0 35712 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_367
timestamp 1679581782
transform 1 0 36384 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_374
timestamp 1679581782
transform 1 0 37056 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_381
timestamp 1679581782
transform 1 0 37728 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_388
timestamp 1679581782
transform 1 0 38400 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_395
timestamp 1679581782
transform 1 0 39072 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_402
timestamp 1679581782
transform 1 0 39744 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_409
timestamp 1679581782
transform 1 0 40416 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_416
timestamp 1679581782
transform 1 0 41088 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_423
timestamp 1679581782
transform 1 0 41760 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_430
timestamp 1679581782
transform 1 0 42432 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_437
timestamp 1679581782
transform 1 0 43104 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_444
timestamp 1679581782
transform 1 0 43776 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_451
timestamp 1679581782
transform 1 0 44448 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_458
timestamp 1679581782
transform 1 0 45120 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_465
timestamp 1679581782
transform 1 0 45792 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_472
timestamp 1679581782
transform 1 0 46464 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_479
timestamp 1679581782
transform 1 0 47136 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_486
timestamp 1679581782
transform 1 0 47808 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_493
timestamp 1679581782
transform 1 0 48480 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_500
timestamp 1679581782
transform 1 0 49152 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_507
timestamp 1679581782
transform 1 0 49824 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_514
timestamp 1679581782
transform 1 0 50496 0 -1 4536
box -48 -56 720 834
use sg13g2_fill_2  FILLER_3_521
timestamp 1677580104
transform 1 0 51168 0 -1 4536
box -48 -56 240 834
use sg13g2_decap_8  FILLER_4_0
timestamp 1679581782
transform 1 0 1152 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_7
timestamp 1679581782
transform 1 0 1824 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_14
timestamp 1679581782
transform 1 0 2496 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_21
timestamp 1679581782
transform 1 0 3168 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_28
timestamp 1679581782
transform 1 0 3840 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_35
timestamp 1679581782
transform 1 0 4512 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_42
timestamp 1679581782
transform 1 0 5184 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_49
timestamp 1679581782
transform 1 0 5856 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_56
timestamp 1679581782
transform 1 0 6528 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_63
timestamp 1679581782
transform 1 0 7200 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_70
timestamp 1679581782
transform 1 0 7872 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_77
timestamp 1679581782
transform 1 0 8544 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_84
timestamp 1679581782
transform 1 0 9216 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_91
timestamp 1679581782
transform 1 0 9888 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_98
timestamp 1679581782
transform 1 0 10560 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_105
timestamp 1679581782
transform 1 0 11232 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_112
timestamp 1679581782
transform 1 0 11904 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_119
timestamp 1679581782
transform 1 0 12576 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_126
timestamp 1679581782
transform 1 0 13248 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_133
timestamp 1679581782
transform 1 0 13920 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_140
timestamp 1679581782
transform 1 0 14592 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_147
timestamp 1679581782
transform 1 0 15264 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_154
timestamp 1679581782
transform 1 0 15936 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_161
timestamp 1679581782
transform 1 0 16608 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_168
timestamp 1679581782
transform 1 0 17280 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_175
timestamp 1679581782
transform 1 0 17952 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_182
timestamp 1679581782
transform 1 0 18624 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_189
timestamp 1679581782
transform 1 0 19296 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_196
timestamp 1679581782
transform 1 0 19968 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_203
timestamp 1679581782
transform 1 0 20640 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_210
timestamp 1679581782
transform 1 0 21312 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_217
timestamp 1679581782
transform 1 0 21984 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_224
timestamp 1679581782
transform 1 0 22656 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_231
timestamp 1679581782
transform 1 0 23328 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_238
timestamp 1679581782
transform 1 0 24000 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_245
timestamp 1679581782
transform 1 0 24672 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_252
timestamp 1679581782
transform 1 0 25344 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_259
timestamp 1679581782
transform 1 0 26016 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_266
timestamp 1679581782
transform 1 0 26688 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_273
timestamp 1679581782
transform 1 0 27360 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_280
timestamp 1679581782
transform 1 0 28032 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_287
timestamp 1679581782
transform 1 0 28704 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_294
timestamp 1679581782
transform 1 0 29376 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_301
timestamp 1679581782
transform 1 0 30048 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_308
timestamp 1679581782
transform 1 0 30720 0 1 4536
box -48 -56 720 834
use sg13g2_fill_2  FILLER_4_315
timestamp 1677580104
transform 1 0 31392 0 1 4536
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_317
timestamp 1677579658
transform 1 0 31584 0 1 4536
box -48 -56 144 834
use sg13g2_fill_2  FILLER_4_322
timestamp 1677580104
transform 1 0 32064 0 1 4536
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_324
timestamp 1677579658
transform 1 0 32256 0 1 4536
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_329
timestamp 1679581782
transform 1 0 32736 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_336
timestamp 1679581782
transform 1 0 33408 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_343
timestamp 1679581782
transform 1 0 34080 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_350
timestamp 1679581782
transform 1 0 34752 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_357
timestamp 1679581782
transform 1 0 35424 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_364
timestamp 1679581782
transform 1 0 36096 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_371
timestamp 1679581782
transform 1 0 36768 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_378
timestamp 1679581782
transform 1 0 37440 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_385
timestamp 1679581782
transform 1 0 38112 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_392
timestamp 1679581782
transform 1 0 38784 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_399
timestamp 1679581782
transform 1 0 39456 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_406
timestamp 1679581782
transform 1 0 40128 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_413
timestamp 1679581782
transform 1 0 40800 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_420
timestamp 1679581782
transform 1 0 41472 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_427
timestamp 1679581782
transform 1 0 42144 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_434
timestamp 1679581782
transform 1 0 42816 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_441
timestamp 1679581782
transform 1 0 43488 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_448
timestamp 1679581782
transform 1 0 44160 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_455
timestamp 1679581782
transform 1 0 44832 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_462
timestamp 1679581782
transform 1 0 45504 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_469
timestamp 1679581782
transform 1 0 46176 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_476
timestamp 1679581782
transform 1 0 46848 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_483
timestamp 1679581782
transform 1 0 47520 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_490
timestamp 1679581782
transform 1 0 48192 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_497
timestamp 1679581782
transform 1 0 48864 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_504
timestamp 1679581782
transform 1 0 49536 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_511
timestamp 1679581782
transform 1 0 50208 0 1 4536
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_518
timestamp 1679577901
transform 1 0 50880 0 1 4536
box -48 -56 432 834
use sg13g2_fill_1  FILLER_4_522
timestamp 1677579658
transform 1 0 51264 0 1 4536
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_0
timestamp 1679581782
transform 1 0 1152 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_7
timestamp 1679581782
transform 1 0 1824 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_14
timestamp 1679581782
transform 1 0 2496 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_21
timestamp 1679581782
transform 1 0 3168 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_28
timestamp 1679581782
transform 1 0 3840 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_35
timestamp 1679581782
transform 1 0 4512 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_42
timestamp 1679581782
transform 1 0 5184 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_49
timestamp 1679581782
transform 1 0 5856 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_56
timestamp 1679581782
transform 1 0 6528 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_63
timestamp 1679581782
transform 1 0 7200 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_70
timestamp 1679581782
transform 1 0 7872 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_77
timestamp 1679581782
transform 1 0 8544 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_84
timestamp 1679581782
transform 1 0 9216 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_91
timestamp 1679581782
transform 1 0 9888 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_98
timestamp 1679581782
transform 1 0 10560 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_105
timestamp 1679581782
transform 1 0 11232 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_112
timestamp 1679581782
transform 1 0 11904 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_119
timestamp 1679581782
transform 1 0 12576 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_126
timestamp 1679581782
transform 1 0 13248 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_133
timestamp 1679581782
transform 1 0 13920 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_140
timestamp 1679581782
transform 1 0 14592 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_147
timestamp 1679581782
transform 1 0 15264 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_154
timestamp 1679581782
transform 1 0 15936 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_161
timestamp 1679581782
transform 1 0 16608 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_168
timestamp 1679581782
transform 1 0 17280 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_175
timestamp 1679581782
transform 1 0 17952 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_182
timestamp 1679581782
transform 1 0 18624 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_189
timestamp 1679581782
transform 1 0 19296 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_196
timestamp 1679581782
transform 1 0 19968 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_203
timestamp 1679581782
transform 1 0 20640 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_210
timestamp 1679581782
transform 1 0 21312 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_217
timestamp 1679581782
transform 1 0 21984 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_224
timestamp 1679581782
transform 1 0 22656 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_231
timestamp 1679581782
transform 1 0 23328 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_238
timestamp 1679581782
transform 1 0 24000 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_245
timestamp 1679581782
transform 1 0 24672 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_252
timestamp 1679581782
transform 1 0 25344 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_259
timestamp 1679581782
transform 1 0 26016 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_270
timestamp 1679577901
transform 1 0 27072 0 -1 6048
box -48 -56 432 834
use sg13g2_fill_1  FILLER_5_274
timestamp 1677579658
transform 1 0 27456 0 -1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_279
timestamp 1679581782
transform 1 0 27936 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_286
timestamp 1679581782
transform 1 0 28608 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_293
timestamp 1679577901
transform 1 0 29280 0 -1 6048
box -48 -56 432 834
use sg13g2_fill_1  FILLER_5_297
timestamp 1677579658
transform 1 0 29664 0 -1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_302
timestamp 1679581782
transform 1 0 30144 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_309
timestamp 1679581782
transform 1 0 30816 0 -1 6048
box -48 -56 720 834
use sg13g2_fill_1  FILLER_5_316
timestamp 1677579658
transform 1 0 31488 0 -1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_321
timestamp 1679581782
transform 1 0 31968 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_328
timestamp 1679577901
transform 1 0 32640 0 -1 6048
box -48 -56 432 834
use sg13g2_decap_8  FILLER_5_336
timestamp 1679581782
transform 1 0 33408 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_343
timestamp 1679581782
transform 1 0 34080 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_350
timestamp 1679581782
transform 1 0 34752 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_357
timestamp 1679581782
transform 1 0 35424 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_364
timestamp 1679581782
transform 1 0 36096 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_371
timestamp 1679581782
transform 1 0 36768 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_378
timestamp 1679581782
transform 1 0 37440 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_385
timestamp 1679581782
transform 1 0 38112 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_392
timestamp 1679581782
transform 1 0 38784 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_399
timestamp 1679581782
transform 1 0 39456 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_406
timestamp 1679581782
transform 1 0 40128 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_413
timestamp 1679581782
transform 1 0 40800 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_420
timestamp 1679581782
transform 1 0 41472 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_427
timestamp 1679581782
transform 1 0 42144 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_434
timestamp 1679581782
transform 1 0 42816 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_441
timestamp 1679581782
transform 1 0 43488 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_448
timestamp 1679581782
transform 1 0 44160 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_455
timestamp 1679581782
transform 1 0 44832 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_462
timestamp 1679581782
transform 1 0 45504 0 -1 6048
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_469
timestamp 1677580104
transform 1 0 46176 0 -1 6048
box -48 -56 240 834
use sg13g2_decap_8  FILLER_5_475
timestamp 1679581782
transform 1 0 46752 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_482
timestamp 1679581782
transform 1 0 47424 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_489
timestamp 1679581782
transform 1 0 48096 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_496
timestamp 1679577901
transform 1 0 48768 0 -1 6048
box -48 -56 432 834
use sg13g2_decap_8  FILLER_5_504
timestamp 1679581782
transform 1 0 49536 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_511
timestamp 1679581782
transform 1 0 50208 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_518
timestamp 1679577901
transform 1 0 50880 0 -1 6048
box -48 -56 432 834
use sg13g2_fill_1  FILLER_5_522
timestamp 1677579658
transform 1 0 51264 0 -1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_0
timestamp 1679581782
transform 1 0 1152 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_7
timestamp 1679581782
transform 1 0 1824 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_14
timestamp 1679581782
transform 1 0 2496 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_21
timestamp 1679581782
transform 1 0 3168 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_28
timestamp 1679581782
transform 1 0 3840 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_35
timestamp 1679581782
transform 1 0 4512 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_42
timestamp 1679581782
transform 1 0 5184 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_49
timestamp 1679581782
transform 1 0 5856 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_56
timestamp 1679581782
transform 1 0 6528 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_63
timestamp 1679581782
transform 1 0 7200 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_70
timestamp 1679581782
transform 1 0 7872 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_77
timestamp 1679581782
transform 1 0 8544 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_84
timestamp 1679581782
transform 1 0 9216 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_91
timestamp 1679581782
transform 1 0 9888 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_98
timestamp 1679581782
transform 1 0 10560 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_105
timestamp 1679581782
transform 1 0 11232 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_112
timestamp 1679581782
transform 1 0 11904 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_119
timestamp 1679581782
transform 1 0 12576 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_126
timestamp 1679581782
transform 1 0 13248 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_133
timestamp 1679581782
transform 1 0 13920 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_140
timestamp 1679581782
transform 1 0 14592 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_147
timestamp 1679581782
transform 1 0 15264 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_154
timestamp 1679581782
transform 1 0 15936 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_161
timestamp 1679581782
transform 1 0 16608 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_168
timestamp 1679581782
transform 1 0 17280 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_175
timestamp 1679581782
transform 1 0 17952 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_182
timestamp 1679581782
transform 1 0 18624 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_189
timestamp 1679581782
transform 1 0 19296 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_196
timestamp 1679581782
transform 1 0 19968 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_203
timestamp 1679581782
transform 1 0 20640 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_210
timestamp 1679581782
transform 1 0 21312 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_217
timestamp 1679581782
transform 1 0 21984 0 1 6048
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_224
timestamp 1679577901
transform 1 0 22656 0 1 6048
box -48 -56 432 834
use sg13g2_fill_1  FILLER_6_228
timestamp 1677579658
transform 1 0 23040 0 1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_237
timestamp 1679581782
transform 1 0 23904 0 1 6048
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_244
timestamp 1679577901
transform 1 0 24576 0 1 6048
box -48 -56 432 834
use sg13g2_fill_2  FILLER_6_252
timestamp 1677580104
transform 1 0 25344 0 1 6048
box -48 -56 240 834
use sg13g2_decap_8  FILLER_6_258
timestamp 1679581782
transform 1 0 25920 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_265
timestamp 1679581782
transform 1 0 26592 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_272
timestamp 1679581782
transform 1 0 27264 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_279
timestamp 1679581782
transform 1 0 27936 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_286
timestamp 1679581782
transform 1 0 28608 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_293
timestamp 1679581782
transform 1 0 29280 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_300
timestamp 1679581782
transform 1 0 29952 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_307
timestamp 1679581782
transform 1 0 30624 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_314
timestamp 1679581782
transform 1 0 31296 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_321
timestamp 1679581782
transform 1 0 31968 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_328
timestamp 1679581782
transform 1 0 32640 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_335
timestamp 1679581782
transform 1 0 33312 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_342
timestamp 1679581782
transform 1 0 33984 0 1 6048
box -48 -56 720 834
use sg13g2_fill_1  FILLER_6_349
timestamp 1677579658
transform 1 0 34656 0 1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_354
timestamp 1679581782
transform 1 0 35136 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_361
timestamp 1679581782
transform 1 0 35808 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_368
timestamp 1679581782
transform 1 0 36480 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_375
timestamp 1679581782
transform 1 0 37152 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_382
timestamp 1679581782
transform 1 0 37824 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_389
timestamp 1679581782
transform 1 0 38496 0 1 6048
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_396
timestamp 1679577901
transform 1 0 39168 0 1 6048
box -48 -56 432 834
use sg13g2_decap_8  FILLER_6_404
timestamp 1679581782
transform 1 0 39936 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_411
timestamp 1679581782
transform 1 0 40608 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_418
timestamp 1679581782
transform 1 0 41280 0 1 6048
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_425
timestamp 1677580104
transform 1 0 41952 0 1 6048
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_427
timestamp 1677579658
transform 1 0 42144 0 1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_432
timestamp 1679581782
transform 1 0 42624 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_439
timestamp 1679581782
transform 1 0 43296 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_446
timestamp 1679581782
transform 1 0 43968 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_453
timestamp 1679581782
transform 1 0 44640 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_460
timestamp 1679581782
transform 1 0 45312 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_467
timestamp 1679581782
transform 1 0 45984 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_474
timestamp 1679581782
transform 1 0 46656 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_481
timestamp 1679581782
transform 1 0 47328 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_488
timestamp 1679581782
transform 1 0 48000 0 1 6048
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_495
timestamp 1679577901
transform 1 0 48672 0 1 6048
box -48 -56 432 834
use sg13g2_fill_2  FILLER_6_499
timestamp 1677580104
transform 1 0 49056 0 1 6048
box -48 -56 240 834
use sg13g2_decap_8  FILLER_6_505
timestamp 1679581782
transform 1 0 49632 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_512
timestamp 1679581782
transform 1 0 50304 0 1 6048
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_519
timestamp 1679577901
transform 1 0 50976 0 1 6048
box -48 -56 432 834
use sg13g2_decap_8  FILLER_7_0
timestamp 1679581782
transform 1 0 1152 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_7
timestamp 1679581782
transform 1 0 1824 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_14
timestamp 1679581782
transform 1 0 2496 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_21
timestamp 1679581782
transform 1 0 3168 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_28
timestamp 1679581782
transform 1 0 3840 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_35
timestamp 1679581782
transform 1 0 4512 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_42
timestamp 1679581782
transform 1 0 5184 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_49
timestamp 1679581782
transform 1 0 5856 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_56
timestamp 1679581782
transform 1 0 6528 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_63
timestamp 1679581782
transform 1 0 7200 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_70
timestamp 1679581782
transform 1 0 7872 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_77
timestamp 1679581782
transform 1 0 8544 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_84
timestamp 1679581782
transform 1 0 9216 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_91
timestamp 1679581782
transform 1 0 9888 0 -1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_7_98
timestamp 1677580104
transform 1 0 10560 0 -1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_100
timestamp 1677579658
transform 1 0 10752 0 -1 7560
box -48 -56 144 834
use sg13g2_fill_1  FILLER_7_109
timestamp 1677579658
transform 1 0 11616 0 -1 7560
box -48 -56 144 834
use sg13g2_fill_2  FILLER_7_114
timestamp 1677580104
transform 1 0 12096 0 -1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_116
timestamp 1677579658
transform 1 0 12288 0 -1 7560
box -48 -56 144 834
use sg13g2_decap_4  FILLER_7_121
timestamp 1679577901
transform 1 0 12768 0 -1 7560
box -48 -56 432 834
use sg13g2_fill_2  FILLER_7_125
timestamp 1677580104
transform 1 0 13152 0 -1 7560
box -48 -56 240 834
use sg13g2_decap_4  FILLER_7_135
timestamp 1679577901
transform 1 0 14112 0 -1 7560
box -48 -56 432 834
use sg13g2_fill_1  FILLER_7_139
timestamp 1677579658
transform 1 0 14496 0 -1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_148
timestamp 1679581782
transform 1 0 15360 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_155
timestamp 1679581782
transform 1 0 16032 0 -1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_7_162
timestamp 1677580104
transform 1 0 16704 0 -1 7560
box -48 -56 240 834
use sg13g2_decap_8  FILLER_7_168
timestamp 1679581782
transform 1 0 17280 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_175
timestamp 1679581782
transform 1 0 17952 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_182
timestamp 1679581782
transform 1 0 18624 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_189
timestamp 1679581782
transform 1 0 19296 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_196
timestamp 1679581782
transform 1 0 19968 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_203
timestamp 1679581782
transform 1 0 20640 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_210
timestamp 1679581782
transform 1 0 21312 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_217
timestamp 1679581782
transform 1 0 21984 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_224
timestamp 1679581782
transform 1 0 22656 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_231
timestamp 1679581782
transform 1 0 23328 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_238
timestamp 1679581782
transform 1 0 24000 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_245
timestamp 1679581782
transform 1 0 24672 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_252
timestamp 1679581782
transform 1 0 25344 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_259
timestamp 1679581782
transform 1 0 26016 0 -1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_7_266
timestamp 1677580104
transform 1 0 26688 0 -1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_268
timestamp 1677579658
transform 1 0 26880 0 -1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_277
timestamp 1679581782
transform 1 0 27744 0 -1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_7_284
timestamp 1677580104
transform 1 0 28416 0 -1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_286
timestamp 1677579658
transform 1 0 28608 0 -1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_291
timestamp 1679581782
transform 1 0 29088 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_298
timestamp 1679581782
transform 1 0 29760 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_305
timestamp 1679581782
transform 1 0 30432 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_312
timestamp 1679581782
transform 1 0 31104 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_319
timestamp 1679581782
transform 1 0 31776 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_326
timestamp 1679581782
transform 1 0 32448 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_333
timestamp 1679581782
transform 1 0 33120 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_340
timestamp 1679581782
transform 1 0 33792 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_347
timestamp 1679581782
transform 1 0 34464 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_354
timestamp 1679581782
transform 1 0 35136 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_361
timestamp 1679581782
transform 1 0 35808 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_368
timestamp 1679581782
transform 1 0 36480 0 -1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_7_375
timestamp 1677580104
transform 1 0 37152 0 -1 7560
box -48 -56 240 834
use sg13g2_fill_2  FILLER_7_381
timestamp 1677580104
transform 1 0 37728 0 -1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_383
timestamp 1677579658
transform 1 0 37920 0 -1 7560
box -48 -56 144 834
use sg13g2_decap_4  FILLER_7_388
timestamp 1679577901
transform 1 0 38400 0 -1 7560
box -48 -56 432 834
use sg13g2_fill_1  FILLER_7_392
timestamp 1677579658
transform 1 0 38784 0 -1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_397
timestamp 1679581782
transform 1 0 39264 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_404
timestamp 1679581782
transform 1 0 39936 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_411
timestamp 1679581782
transform 1 0 40608 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_418
timestamp 1679581782
transform 1 0 41280 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_425
timestamp 1679581782
transform 1 0 41952 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_432
timestamp 1679581782
transform 1 0 42624 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_439
timestamp 1679581782
transform 1 0 43296 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_446
timestamp 1679581782
transform 1 0 43968 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_453
timestamp 1679581782
transform 1 0 44640 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_460
timestamp 1679581782
transform 1 0 45312 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_467
timestamp 1679581782
transform 1 0 45984 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_474
timestamp 1679581782
transform 1 0 46656 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_481
timestamp 1679581782
transform 1 0 47328 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_488
timestamp 1679581782
transform 1 0 48000 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_495
timestamp 1679581782
transform 1 0 48672 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_502
timestamp 1679581782
transform 1 0 49344 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_509
timestamp 1679581782
transform 1 0 50016 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_516
timestamp 1679581782
transform 1 0 50688 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_0
timestamp 1679581782
transform 1 0 1152 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_7
timestamp 1679581782
transform 1 0 1824 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_14
timestamp 1679581782
transform 1 0 2496 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_25
timestamp 1679581782
transform 1 0 3552 0 1 7560
box -48 -56 720 834
use sg13g2_fill_1  FILLER_8_32
timestamp 1677579658
transform 1 0 4224 0 1 7560
box -48 -56 144 834
use sg13g2_decap_4  FILLER_8_37
timestamp 1679577901
transform 1 0 4704 0 1 7560
box -48 -56 432 834
use sg13g2_fill_1  FILLER_8_41
timestamp 1677579658
transform 1 0 5088 0 1 7560
box -48 -56 144 834
use sg13g2_decap_4  FILLER_8_46
timestamp 1679577901
transform 1 0 5568 0 1 7560
box -48 -56 432 834
use sg13g2_fill_1  FILLER_8_50
timestamp 1677579658
transform 1 0 5952 0 1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_55
timestamp 1679581782
transform 1 0 6432 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_62
timestamp 1679581782
transform 1 0 7104 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_77
timestamp 1679581782
transform 1 0 8544 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_84
timestamp 1679581782
transform 1 0 9216 0 1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_8_91
timestamp 1677580104
transform 1 0 9888 0 1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_93
timestamp 1677579658
transform 1 0 10080 0 1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_102
timestamp 1679581782
transform 1 0 10944 0 1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_8_109
timestamp 1677580104
transform 1 0 11616 0 1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_111
timestamp 1677579658
transform 1 0 11808 0 1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_116
timestamp 1679581782
transform 1 0 12288 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_123
timestamp 1679581782
transform 1 0 12960 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_130
timestamp 1679581782
transform 1 0 13632 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_137
timestamp 1679581782
transform 1 0 14304 0 1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_8_144
timestamp 1677580104
transform 1 0 14976 0 1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_146
timestamp 1677579658
transform 1 0 15168 0 1 7560
box -48 -56 144 834
use sg13g2_fill_2  FILLER_8_183
timestamp 1677580104
transform 1 0 18720 0 1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_185
timestamp 1677579658
transform 1 0 18912 0 1 7560
box -48 -56 144 834
use sg13g2_decap_4  FILLER_8_194
timestamp 1679577901
transform 1 0 19776 0 1 7560
box -48 -56 432 834
use sg13g2_fill_1  FILLER_8_198
timestamp 1677579658
transform 1 0 20160 0 1 7560
box -48 -56 144 834
use sg13g2_fill_1  FILLER_8_203
timestamp 1677579658
transform 1 0 20640 0 1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_208
timestamp 1679581782
transform 1 0 21120 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_215
timestamp 1679581782
transform 1 0 21792 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_222
timestamp 1679581782
transform 1 0 22464 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_229
timestamp 1679581782
transform 1 0 23136 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_236
timestamp 1679581782
transform 1 0 23808 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_243
timestamp 1679581782
transform 1 0 24480 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_250
timestamp 1679581782
transform 1 0 25152 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_257
timestamp 1679581782
transform 1 0 25824 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_264
timestamp 1679581782
transform 1 0 26496 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_271
timestamp 1679581782
transform 1 0 27168 0 1 7560
box -48 -56 720 834
use sg13g2_decap_4  FILLER_8_278
timestamp 1679577901
transform 1 0 27840 0 1 7560
box -48 -56 432 834
use sg13g2_fill_1  FILLER_8_282
timestamp 1677579658
transform 1 0 28224 0 1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_287
timestamp 1679581782
transform 1 0 28704 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_294
timestamp 1679581782
transform 1 0 29376 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_301
timestamp 1679581782
transform 1 0 30048 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_308
timestamp 1679581782
transform 1 0 30720 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_315
timestamp 1679581782
transform 1 0 31392 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_322
timestamp 1679581782
transform 1 0 32064 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_341
timestamp 1679581782
transform 1 0 33888 0 1 7560
box -48 -56 720 834
use sg13g2_fill_1  FILLER_8_348
timestamp 1677579658
transform 1 0 34560 0 1 7560
box -48 -56 144 834
use sg13g2_fill_1  FILLER_8_365
timestamp 1677579658
transform 1 0 36192 0 1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_406
timestamp 1679581782
transform 1 0 40128 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_413
timestamp 1679581782
transform 1 0 40800 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_420
timestamp 1679581782
transform 1 0 41472 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_427
timestamp 1679581782
transform 1 0 42144 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_434
timestamp 1679581782
transform 1 0 42816 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_441
timestamp 1679581782
transform 1 0 43488 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_448
timestamp 1679581782
transform 1 0 44160 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_455
timestamp 1679581782
transform 1 0 44832 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_462
timestamp 1679581782
transform 1 0 45504 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_469
timestamp 1679581782
transform 1 0 46176 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_476
timestamp 1679581782
transform 1 0 46848 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_483
timestamp 1679581782
transform 1 0 47520 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_490
timestamp 1679581782
transform 1 0 48192 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_497
timestamp 1679581782
transform 1 0 48864 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_504
timestamp 1679581782
transform 1 0 49536 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_511
timestamp 1679581782
transform 1 0 50208 0 1 7560
box -48 -56 720 834
use sg13g2_fill_1  FILLER_8_518
timestamp 1677579658
transform 1 0 50880 0 1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_0
timestamp 1679581782
transform 1 0 1152 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_7
timestamp 1679581782
transform 1 0 1824 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_14
timestamp 1679581782
transform 1 0 2496 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_21
timestamp 1679581782
transform 1 0 3168 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_28
timestamp 1679581782
transform 1 0 3840 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_35
timestamp 1679581782
transform 1 0 4512 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_42
timestamp 1679581782
transform 1 0 5184 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_49
timestamp 1679581782
transform 1 0 5856 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_56
timestamp 1679581782
transform 1 0 6528 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_63
timestamp 1679581782
transform 1 0 7200 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_70
timestamp 1679581782
transform 1 0 7872 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_77
timestamp 1679581782
transform 1 0 8544 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_84
timestamp 1679581782
transform 1 0 9216 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_91
timestamp 1679581782
transform 1 0 9888 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_98
timestamp 1679581782
transform 1 0 10560 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_105
timestamp 1679581782
transform 1 0 11232 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_112
timestamp 1679581782
transform 1 0 11904 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_119
timestamp 1679581782
transform 1 0 12576 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_126
timestamp 1679581782
transform 1 0 13248 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_133
timestamp 1679581782
transform 1 0 13920 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_140
timestamp 1679581782
transform 1 0 14592 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_147
timestamp 1679581782
transform 1 0 15264 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_154
timestamp 1679581782
transform 1 0 15936 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_161
timestamp 1679581782
transform 1 0 16608 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_168
timestamp 1679581782
transform 1 0 17280 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_175
timestamp 1679581782
transform 1 0 17952 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_182
timestamp 1679581782
transform 1 0 18624 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_189
timestamp 1679581782
transform 1 0 19296 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_196
timestamp 1679581782
transform 1 0 19968 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_203
timestamp 1679581782
transform 1 0 20640 0 -1 9072
box -48 -56 720 834
use sg13g2_fill_2  FILLER_9_210
timestamp 1677580104
transform 1 0 21312 0 -1 9072
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_212
timestamp 1677579658
transform 1 0 21504 0 -1 9072
box -48 -56 144 834
use sg13g2_fill_1  FILLER_9_217
timestamp 1677579658
transform 1 0 21984 0 -1 9072
box -48 -56 144 834
use sg13g2_fill_2  FILLER_9_226
timestamp 1677580104
transform 1 0 22848 0 -1 9072
box -48 -56 240 834
use sg13g2_fill_2  FILLER_9_232
timestamp 1677580104
transform 1 0 23424 0 -1 9072
box -48 -56 240 834
use sg13g2_decap_8  FILLER_9_238
timestamp 1679581782
transform 1 0 24000 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_245
timestamp 1679581782
transform 1 0 24672 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_252
timestamp 1679581782
transform 1 0 25344 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_259
timestamp 1679581782
transform 1 0 26016 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_298
timestamp 1679581782
transform 1 0 29760 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_305
timestamp 1679581782
transform 1 0 30432 0 -1 9072
box -48 -56 720 834
use sg13g2_fill_1  FILLER_9_312
timestamp 1677579658
transform 1 0 31104 0 -1 9072
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_317
timestamp 1679581782
transform 1 0 31584 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_324
timestamp 1679581782
transform 1 0 32256 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_331
timestamp 1679581782
transform 1 0 32928 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_338
timestamp 1679581782
transform 1 0 33600 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_345
timestamp 1679581782
transform 1 0 34272 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_352
timestamp 1679581782
transform 1 0 34944 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_359
timestamp 1679581782
transform 1 0 35616 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_366
timestamp 1679581782
transform 1 0 36288 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_373
timestamp 1679581782
transform 1 0 36960 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_380
timestamp 1679581782
transform 1 0 37632 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_387
timestamp 1679581782
transform 1 0 38304 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_394
timestamp 1679581782
transform 1 0 38976 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_401
timestamp 1679581782
transform 1 0 39648 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_408
timestamp 1679581782
transform 1 0 40320 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_415
timestamp 1679581782
transform 1 0 40992 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_422
timestamp 1679581782
transform 1 0 41664 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_429
timestamp 1679581782
transform 1 0 42336 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_436
timestamp 1679581782
transform 1 0 43008 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_443
timestamp 1679581782
transform 1 0 43680 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_450
timestamp 1679581782
transform 1 0 44352 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_457
timestamp 1679581782
transform 1 0 45024 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_464
timestamp 1679581782
transform 1 0 45696 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_471
timestamp 1679581782
transform 1 0 46368 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_478
timestamp 1679581782
transform 1 0 47040 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_485
timestamp 1679581782
transform 1 0 47712 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_492
timestamp 1679581782
transform 1 0 48384 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_499
timestamp 1679581782
transform 1 0 49056 0 -1 9072
box -48 -56 720 834
use sg13g2_fill_1  FILLER_9_506
timestamp 1677579658
transform 1 0 49728 0 -1 9072
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_0
timestamp 1679581782
transform 1 0 1152 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_7
timestamp 1679581782
transform 1 0 1824 0 1 9072
box -48 -56 720 834
use sg13g2_fill_2  FILLER_10_14
timestamp 1677580104
transform 1 0 2496 0 1 9072
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_16
timestamp 1677579658
transform 1 0 2688 0 1 9072
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_225
timestamp 1679581782
transform 1 0 22752 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_232
timestamp 1679581782
transform 1 0 23424 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_239
timestamp 1679581782
transform 1 0 24096 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_246
timestamp 1679581782
transform 1 0 24768 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_253
timestamp 1679581782
transform 1 0 25440 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_260
timestamp 1679581782
transform 1 0 26112 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_267
timestamp 1679581782
transform 1 0 26784 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_274
timestamp 1679581782
transform 1 0 27456 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_281
timestamp 1679581782
transform 1 0 28128 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_288
timestamp 1679581782
transform 1 0 28800 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_295
timestamp 1679581782
transform 1 0 29472 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_302
timestamp 1679581782
transform 1 0 30144 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_309
timestamp 1679581782
transform 1 0 30816 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_316
timestamp 1679581782
transform 1 0 31488 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_323
timestamp 1679581782
transform 1 0 32160 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_330
timestamp 1679581782
transform 1 0 32832 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_337
timestamp 1679581782
transform 1 0 33504 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_344
timestamp 1679581782
transform 1 0 34176 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_351
timestamp 1679581782
transform 1 0 34848 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_358
timestamp 1679581782
transform 1 0 35520 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_365
timestamp 1679581782
transform 1 0 36192 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_372
timestamp 1679581782
transform 1 0 36864 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_379
timestamp 1679581782
transform 1 0 37536 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_386
timestamp 1679581782
transform 1 0 38208 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_393
timestamp 1679581782
transform 1 0 38880 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_400
timestamp 1679581782
transform 1 0 39552 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_407
timestamp 1679581782
transform 1 0 40224 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_414
timestamp 1679581782
transform 1 0 40896 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_421
timestamp 1679581782
transform 1 0 41568 0 1 9072
box -48 -56 720 834
use sg13g2_decap_4  FILLER_10_428
timestamp 1679577901
transform 1 0 42240 0 1 9072
box -48 -56 432 834
use sg13g2_fill_1  FILLER_10_432
timestamp 1677579658
transform 1 0 42624 0 1 9072
box -48 -56 144 834
use sg13g2_fill_2  FILLER_10_517
timestamp 1677580104
transform 1 0 50784 0 1 9072
box -48 -56 240 834
use sg13g2_buf_1  output1
timestamp 1676381911
transform 1 0 50976 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output2
timestamp 1676381911
transform 1 0 51360 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output3
timestamp 1676381911
transform 1 0 51744 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output4
timestamp 1676381911
transform 1 0 51360 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output5
timestamp 1676381911
transform 1 0 51744 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output6
timestamp 1676381911
transform 1 0 51360 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output7
timestamp 1676381911
transform 1 0 51744 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output8
timestamp 1676381911
transform 1 0 51360 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  output9
timestamp 1676381911
transform 1 0 51744 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  output10
timestamp 1676381911
transform 1 0 51360 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  output11
timestamp 1676381911
transform 1 0 51744 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  output12
timestamp 1676381911
transform 1 0 50592 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output13
timestamp 1676381911
transform 1 0 51744 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  output14
timestamp 1676381911
transform 1 0 51360 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  output15
timestamp 1676381911
transform 1 0 51744 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output16
timestamp 1676381911
transform 1 0 51360 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output17
timestamp 1676381911
transform 1 0 51744 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output18
timestamp 1676381911
transform 1 0 51360 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output19
timestamp 1676381911
transform 1 0 50976 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output20
timestamp 1676381911
transform 1 0 50976 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output21
timestamp 1676381911
transform 1 0 50592 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output22
timestamp 1676381911
transform 1 0 50976 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  output23
timestamp 1676381911
transform 1 0 50208 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output24
timestamp 1676381911
transform 1 0 50208 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output25
timestamp 1676381911
transform 1 0 49824 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output26
timestamp 1676381911
transform 1 0 51360 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output27
timestamp 1676381911
transform 1 0 50976 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output28
timestamp 1676381911
transform 1 0 51744 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output29
timestamp 1676381911
transform 1 0 51360 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output30
timestamp 1676381911
transform 1 0 51744 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output31
timestamp 1676381911
transform 1 0 51360 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output32
timestamp 1676381911
transform 1 0 51744 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output33
timestamp 1676381911
transform -1 0 43488 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output34
timestamp 1676381911
transform -1 0 47328 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output35
timestamp 1676381911
transform -1 0 47712 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output36
timestamp 1676381911
transform -1 0 48096 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output37
timestamp 1676381911
transform -1 0 48480 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output38
timestamp 1676381911
transform -1 0 48864 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output39
timestamp 1676381911
transform -1 0 49248 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output40
timestamp 1676381911
transform -1 0 49632 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output41
timestamp 1676381911
transform -1 0 50016 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output42
timestamp 1676381911
transform -1 0 50400 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output43
timestamp 1676381911
transform -1 0 50784 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output44
timestamp 1676381911
transform -1 0 43872 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output45
timestamp 1676381911
transform -1 0 44256 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output46
timestamp 1676381911
transform -1 0 44640 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output47
timestamp 1676381911
transform -1 0 45024 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output48
timestamp 1676381911
transform -1 0 45408 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output49
timestamp 1676381911
transform -1 0 45792 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output50
timestamp 1676381911
transform -1 0 46176 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output51
timestamp 1676381911
transform -1 0 46560 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output52
timestamp 1676381911
transform -1 0 46944 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output53
timestamp 1676381911
transform -1 0 3168 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output54
timestamp 1676381911
transform -1 0 3552 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output55
timestamp 1676381911
transform -1 0 3936 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output56
timestamp 1676381911
transform -1 0 4320 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output57
timestamp 1676381911
transform -1 0 4704 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output58
timestamp 1676381911
transform -1 0 5088 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output59
timestamp 1676381911
transform -1 0 5472 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output60
timestamp 1676381911
transform -1 0 5856 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output61
timestamp 1676381911
transform -1 0 6240 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output62
timestamp 1676381911
transform -1 0 6624 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output63
timestamp 1676381911
transform -1 0 7008 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output64
timestamp 1676381911
transform -1 0 7392 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output65
timestamp 1676381911
transform -1 0 7776 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output66
timestamp 1676381911
transform -1 0 8160 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output67
timestamp 1676381911
transform -1 0 8544 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output68
timestamp 1676381911
transform -1 0 8928 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output69
timestamp 1676381911
transform -1 0 9312 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output70
timestamp 1676381911
transform -1 0 9696 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output71
timestamp 1676381911
transform -1 0 10080 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output72
timestamp 1676381911
transform -1 0 10464 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output73
timestamp 1676381911
transform -1 0 10848 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output74
timestamp 1676381911
transform -1 0 14688 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output75
timestamp 1676381911
transform -1 0 15072 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output76
timestamp 1676381911
transform -1 0 15456 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output77
timestamp 1676381911
transform -1 0 15840 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output78
timestamp 1676381911
transform -1 0 16224 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output79
timestamp 1676381911
transform -1 0 16608 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output80
timestamp 1676381911
transform -1 0 11232 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output81
timestamp 1676381911
transform -1 0 11616 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output82
timestamp 1676381911
transform -1 0 12000 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output83
timestamp 1676381911
transform -1 0 12384 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output84
timestamp 1676381911
transform -1 0 12768 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output85
timestamp 1676381911
transform -1 0 13152 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output86
timestamp 1676381911
transform -1 0 13536 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output87
timestamp 1676381911
transform -1 0 13920 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output88
timestamp 1676381911
transform -1 0 14304 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output89
timestamp 1676381911
transform -1 0 16992 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output90
timestamp 1676381911
transform -1 0 20832 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output91
timestamp 1676381911
transform -1 0 21216 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output92
timestamp 1676381911
transform -1 0 21600 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output93
timestamp 1676381911
transform -1 0 21984 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output94
timestamp 1676381911
transform -1 0 22368 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output95
timestamp 1676381911
transform -1 0 22752 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output96
timestamp 1676381911
transform -1 0 17376 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output97
timestamp 1676381911
transform -1 0 17760 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output98
timestamp 1676381911
transform -1 0 18144 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output99
timestamp 1676381911
transform -1 0 18528 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output100
timestamp 1676381911
transform -1 0 18912 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output101
timestamp 1676381911
transform -1 0 19296 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output102
timestamp 1676381911
transform -1 0 19680 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output103
timestamp 1676381911
transform -1 0 20064 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output104
timestamp 1676381911
transform -1 0 20448 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output105
timestamp 1676381911
transform -1 0 43104 0 1 9072
box -48 -56 432 834
<< labels >>
flabel metal2 s 0 548 90 628 0 FreeSans 320 0 0 0 FrameData[0]
port 0 nsew signal input
flabel metal2 s 0 3908 90 3988 0 FreeSans 320 0 0 0 FrameData[10]
port 1 nsew signal input
flabel metal2 s 0 4244 90 4324 0 FreeSans 320 0 0 0 FrameData[11]
port 2 nsew signal input
flabel metal2 s 0 4580 90 4660 0 FreeSans 320 0 0 0 FrameData[12]
port 3 nsew signal input
flabel metal2 s 0 4916 90 4996 0 FreeSans 320 0 0 0 FrameData[13]
port 4 nsew signal input
flabel metal2 s 0 5252 90 5332 0 FreeSans 320 0 0 0 FrameData[14]
port 5 nsew signal input
flabel metal2 s 0 5588 90 5668 0 FreeSans 320 0 0 0 FrameData[15]
port 6 nsew signal input
flabel metal2 s 0 5924 90 6004 0 FreeSans 320 0 0 0 FrameData[16]
port 7 nsew signal input
flabel metal2 s 0 6260 90 6340 0 FreeSans 320 0 0 0 FrameData[17]
port 8 nsew signal input
flabel metal2 s 0 6596 90 6676 0 FreeSans 320 0 0 0 FrameData[18]
port 9 nsew signal input
flabel metal2 s 0 6932 90 7012 0 FreeSans 320 0 0 0 FrameData[19]
port 10 nsew signal input
flabel metal2 s 0 884 90 964 0 FreeSans 320 0 0 0 FrameData[1]
port 11 nsew signal input
flabel metal2 s 0 7268 90 7348 0 FreeSans 320 0 0 0 FrameData[20]
port 12 nsew signal input
flabel metal2 s 0 7604 90 7684 0 FreeSans 320 0 0 0 FrameData[21]
port 13 nsew signal input
flabel metal2 s 0 7940 90 8020 0 FreeSans 320 0 0 0 FrameData[22]
port 14 nsew signal input
flabel metal2 s 0 8276 90 8356 0 FreeSans 320 0 0 0 FrameData[23]
port 15 nsew signal input
flabel metal2 s 0 8612 90 8692 0 FreeSans 320 0 0 0 FrameData[24]
port 16 nsew signal input
flabel metal2 s 0 8948 90 9028 0 FreeSans 320 0 0 0 FrameData[25]
port 17 nsew signal input
flabel metal2 s 0 9284 90 9364 0 FreeSans 320 0 0 0 FrameData[26]
port 18 nsew signal input
flabel metal2 s 0 9620 90 9700 0 FreeSans 320 0 0 0 FrameData[27]
port 19 nsew signal input
flabel metal2 s 0 9956 90 10036 0 FreeSans 320 0 0 0 FrameData[28]
port 20 nsew signal input
flabel metal2 s 0 10292 90 10372 0 FreeSans 320 0 0 0 FrameData[29]
port 21 nsew signal input
flabel metal2 s 0 1220 90 1300 0 FreeSans 320 0 0 0 FrameData[2]
port 22 nsew signal input
flabel metal2 s 0 10628 90 10708 0 FreeSans 320 0 0 0 FrameData[30]
port 23 nsew signal input
flabel metal2 s 0 10964 90 11044 0 FreeSans 320 0 0 0 FrameData[31]
port 24 nsew signal input
flabel metal2 s 0 1556 90 1636 0 FreeSans 320 0 0 0 FrameData[3]
port 25 nsew signal input
flabel metal2 s 0 1892 90 1972 0 FreeSans 320 0 0 0 FrameData[4]
port 26 nsew signal input
flabel metal2 s 0 2228 90 2308 0 FreeSans 320 0 0 0 FrameData[5]
port 27 nsew signal input
flabel metal2 s 0 2564 90 2644 0 FreeSans 320 0 0 0 FrameData[6]
port 28 nsew signal input
flabel metal2 s 0 2900 90 2980 0 FreeSans 320 0 0 0 FrameData[7]
port 29 nsew signal input
flabel metal2 s 0 3236 90 3316 0 FreeSans 320 0 0 0 FrameData[8]
port 30 nsew signal input
flabel metal2 s 0 3572 90 3652 0 FreeSans 320 0 0 0 FrameData[9]
port 31 nsew signal input
flabel metal2 s 53190 548 53280 628 0 FreeSans 320 0 0 0 FrameData_O[0]
port 32 nsew signal output
flabel metal2 s 53190 3908 53280 3988 0 FreeSans 320 0 0 0 FrameData_O[10]
port 33 nsew signal output
flabel metal2 s 53190 4244 53280 4324 0 FreeSans 320 0 0 0 FrameData_O[11]
port 34 nsew signal output
flabel metal2 s 53190 4580 53280 4660 0 FreeSans 320 0 0 0 FrameData_O[12]
port 35 nsew signal output
flabel metal2 s 53190 4916 53280 4996 0 FreeSans 320 0 0 0 FrameData_O[13]
port 36 nsew signal output
flabel metal2 s 53190 5252 53280 5332 0 FreeSans 320 0 0 0 FrameData_O[14]
port 37 nsew signal output
flabel metal2 s 53190 5588 53280 5668 0 FreeSans 320 0 0 0 FrameData_O[15]
port 38 nsew signal output
flabel metal2 s 53190 5924 53280 6004 0 FreeSans 320 0 0 0 FrameData_O[16]
port 39 nsew signal output
flabel metal2 s 53190 6260 53280 6340 0 FreeSans 320 0 0 0 FrameData_O[17]
port 40 nsew signal output
flabel metal2 s 53190 6596 53280 6676 0 FreeSans 320 0 0 0 FrameData_O[18]
port 41 nsew signal output
flabel metal2 s 53190 6932 53280 7012 0 FreeSans 320 0 0 0 FrameData_O[19]
port 42 nsew signal output
flabel metal2 s 53190 884 53280 964 0 FreeSans 320 0 0 0 FrameData_O[1]
port 43 nsew signal output
flabel metal2 s 53190 7268 53280 7348 0 FreeSans 320 0 0 0 FrameData_O[20]
port 44 nsew signal output
flabel metal2 s 53190 7604 53280 7684 0 FreeSans 320 0 0 0 FrameData_O[21]
port 45 nsew signal output
flabel metal2 s 53190 7940 53280 8020 0 FreeSans 320 0 0 0 FrameData_O[22]
port 46 nsew signal output
flabel metal2 s 53190 8276 53280 8356 0 FreeSans 320 0 0 0 FrameData_O[23]
port 47 nsew signal output
flabel metal2 s 53190 8612 53280 8692 0 FreeSans 320 0 0 0 FrameData_O[24]
port 48 nsew signal output
flabel metal2 s 53190 8948 53280 9028 0 FreeSans 320 0 0 0 FrameData_O[25]
port 49 nsew signal output
flabel metal2 s 53190 9284 53280 9364 0 FreeSans 320 0 0 0 FrameData_O[26]
port 50 nsew signal output
flabel metal2 s 53190 9620 53280 9700 0 FreeSans 320 0 0 0 FrameData_O[27]
port 51 nsew signal output
flabel metal2 s 53190 9956 53280 10036 0 FreeSans 320 0 0 0 FrameData_O[28]
port 52 nsew signal output
flabel metal2 s 53190 10292 53280 10372 0 FreeSans 320 0 0 0 FrameData_O[29]
port 53 nsew signal output
flabel metal2 s 53190 1220 53280 1300 0 FreeSans 320 0 0 0 FrameData_O[2]
port 54 nsew signal output
flabel metal2 s 53190 10628 53280 10708 0 FreeSans 320 0 0 0 FrameData_O[30]
port 55 nsew signal output
flabel metal2 s 53190 10964 53280 11044 0 FreeSans 320 0 0 0 FrameData_O[31]
port 56 nsew signal output
flabel metal2 s 53190 1556 53280 1636 0 FreeSans 320 0 0 0 FrameData_O[3]
port 57 nsew signal output
flabel metal2 s 53190 1892 53280 1972 0 FreeSans 320 0 0 0 FrameData_O[4]
port 58 nsew signal output
flabel metal2 s 53190 2228 53280 2308 0 FreeSans 320 0 0 0 FrameData_O[5]
port 59 nsew signal output
flabel metal2 s 53190 2564 53280 2644 0 FreeSans 320 0 0 0 FrameData_O[6]
port 60 nsew signal output
flabel metal2 s 53190 2900 53280 2980 0 FreeSans 320 0 0 0 FrameData_O[7]
port 61 nsew signal output
flabel metal2 s 53190 3236 53280 3316 0 FreeSans 320 0 0 0 FrameData_O[8]
port 62 nsew signal output
flabel metal2 s 53190 3572 53280 3652 0 FreeSans 320 0 0 0 FrameData_O[9]
port 63 nsew signal output
flabel metal3 s 4088 0 4168 80 0 FreeSans 320 0 0 0 FrameStrobe[0]
port 64 nsew signal input
flabel metal3 s 29048 0 29128 80 0 FreeSans 320 0 0 0 FrameStrobe[10]
port 65 nsew signal input
flabel metal3 s 31544 0 31624 80 0 FreeSans 320 0 0 0 FrameStrobe[11]
port 66 nsew signal input
flabel metal3 s 34040 0 34120 80 0 FreeSans 320 0 0 0 FrameStrobe[12]
port 67 nsew signal input
flabel metal3 s 36536 0 36616 80 0 FreeSans 320 0 0 0 FrameStrobe[13]
port 68 nsew signal input
flabel metal3 s 39032 0 39112 80 0 FreeSans 320 0 0 0 FrameStrobe[14]
port 69 nsew signal input
flabel metal3 s 41528 0 41608 80 0 FreeSans 320 0 0 0 FrameStrobe[15]
port 70 nsew signal input
flabel metal3 s 44024 0 44104 80 0 FreeSans 320 0 0 0 FrameStrobe[16]
port 71 nsew signal input
flabel metal3 s 46520 0 46600 80 0 FreeSans 320 0 0 0 FrameStrobe[17]
port 72 nsew signal input
flabel metal3 s 49016 0 49096 80 0 FreeSans 320 0 0 0 FrameStrobe[18]
port 73 nsew signal input
flabel metal3 s 51512 0 51592 80 0 FreeSans 320 0 0 0 FrameStrobe[19]
port 74 nsew signal input
flabel metal3 s 6584 0 6664 80 0 FreeSans 320 0 0 0 FrameStrobe[1]
port 75 nsew signal input
flabel metal3 s 9080 0 9160 80 0 FreeSans 320 0 0 0 FrameStrobe[2]
port 76 nsew signal input
flabel metal3 s 11576 0 11656 80 0 FreeSans 320 0 0 0 FrameStrobe[3]
port 77 nsew signal input
flabel metal3 s 14072 0 14152 80 0 FreeSans 320 0 0 0 FrameStrobe[4]
port 78 nsew signal input
flabel metal3 s 16568 0 16648 80 0 FreeSans 320 0 0 0 FrameStrobe[5]
port 79 nsew signal input
flabel metal3 s 19064 0 19144 80 0 FreeSans 320 0 0 0 FrameStrobe[6]
port 80 nsew signal input
flabel metal3 s 21560 0 21640 80 0 FreeSans 320 0 0 0 FrameStrobe[7]
port 81 nsew signal input
flabel metal3 s 24056 0 24136 80 0 FreeSans 320 0 0 0 FrameStrobe[8]
port 82 nsew signal input
flabel metal3 s 26552 0 26632 80 0 FreeSans 320 0 0 0 FrameStrobe[9]
port 83 nsew signal input
flabel metal3 s 43064 11764 43144 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[0]
port 84 nsew signal output
flabel metal3 s 46904 11764 46984 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[10]
port 85 nsew signal output
flabel metal3 s 47288 11764 47368 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[11]
port 86 nsew signal output
flabel metal3 s 47672 11764 47752 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[12]
port 87 nsew signal output
flabel metal3 s 48056 11764 48136 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[13]
port 88 nsew signal output
flabel metal3 s 48440 11764 48520 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[14]
port 89 nsew signal output
flabel metal3 s 48824 11764 48904 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[15]
port 90 nsew signal output
flabel metal3 s 49208 11764 49288 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[16]
port 91 nsew signal output
flabel metal3 s 49592 11764 49672 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[17]
port 92 nsew signal output
flabel metal3 s 49976 11764 50056 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[18]
port 93 nsew signal output
flabel metal3 s 50360 11764 50440 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[19]
port 94 nsew signal output
flabel metal3 s 43448 11764 43528 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[1]
port 95 nsew signal output
flabel metal3 s 43832 11764 43912 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[2]
port 96 nsew signal output
flabel metal3 s 44216 11764 44296 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[3]
port 97 nsew signal output
flabel metal3 s 44600 11764 44680 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[4]
port 98 nsew signal output
flabel metal3 s 44984 11764 45064 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[5]
port 99 nsew signal output
flabel metal3 s 45368 11764 45448 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[6]
port 100 nsew signal output
flabel metal3 s 45752 11764 45832 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[7]
port 101 nsew signal output
flabel metal3 s 46136 11764 46216 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[8]
port 102 nsew signal output
flabel metal3 s 46520 11764 46600 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[9]
port 103 nsew signal output
flabel metal3 s 2744 11764 2824 11844 0 FreeSans 320 0 0 0 N1BEG[0]
port 104 nsew signal output
flabel metal3 s 3128 11764 3208 11844 0 FreeSans 320 0 0 0 N1BEG[1]
port 105 nsew signal output
flabel metal3 s 3512 11764 3592 11844 0 FreeSans 320 0 0 0 N1BEG[2]
port 106 nsew signal output
flabel metal3 s 3896 11764 3976 11844 0 FreeSans 320 0 0 0 N1BEG[3]
port 107 nsew signal output
flabel metal3 s 4280 11764 4360 11844 0 FreeSans 320 0 0 0 N2BEG[0]
port 108 nsew signal output
flabel metal3 s 4664 11764 4744 11844 0 FreeSans 320 0 0 0 N2BEG[1]
port 109 nsew signal output
flabel metal3 s 5048 11764 5128 11844 0 FreeSans 320 0 0 0 N2BEG[2]
port 110 nsew signal output
flabel metal3 s 5432 11764 5512 11844 0 FreeSans 320 0 0 0 N2BEG[3]
port 111 nsew signal output
flabel metal3 s 5816 11764 5896 11844 0 FreeSans 320 0 0 0 N2BEG[4]
port 112 nsew signal output
flabel metal3 s 6200 11764 6280 11844 0 FreeSans 320 0 0 0 N2BEG[5]
port 113 nsew signal output
flabel metal3 s 6584 11764 6664 11844 0 FreeSans 320 0 0 0 N2BEG[6]
port 114 nsew signal output
flabel metal3 s 6968 11764 7048 11844 0 FreeSans 320 0 0 0 N2BEG[7]
port 115 nsew signal output
flabel metal3 s 7352 11764 7432 11844 0 FreeSans 320 0 0 0 N2BEGb[0]
port 116 nsew signal output
flabel metal3 s 7736 11764 7816 11844 0 FreeSans 320 0 0 0 N2BEGb[1]
port 117 nsew signal output
flabel metal3 s 8120 11764 8200 11844 0 FreeSans 320 0 0 0 N2BEGb[2]
port 118 nsew signal output
flabel metal3 s 8504 11764 8584 11844 0 FreeSans 320 0 0 0 N2BEGb[3]
port 119 nsew signal output
flabel metal3 s 8888 11764 8968 11844 0 FreeSans 320 0 0 0 N2BEGb[4]
port 120 nsew signal output
flabel metal3 s 9272 11764 9352 11844 0 FreeSans 320 0 0 0 N2BEGb[5]
port 121 nsew signal output
flabel metal3 s 9656 11764 9736 11844 0 FreeSans 320 0 0 0 N2BEGb[6]
port 122 nsew signal output
flabel metal3 s 10040 11764 10120 11844 0 FreeSans 320 0 0 0 N2BEGb[7]
port 123 nsew signal output
flabel metal3 s 10424 11764 10504 11844 0 FreeSans 320 0 0 0 N4BEG[0]
port 124 nsew signal output
flabel metal3 s 14264 11764 14344 11844 0 FreeSans 320 0 0 0 N4BEG[10]
port 125 nsew signal output
flabel metal3 s 14648 11764 14728 11844 0 FreeSans 320 0 0 0 N4BEG[11]
port 126 nsew signal output
flabel metal3 s 15032 11764 15112 11844 0 FreeSans 320 0 0 0 N4BEG[12]
port 127 nsew signal output
flabel metal3 s 15416 11764 15496 11844 0 FreeSans 320 0 0 0 N4BEG[13]
port 128 nsew signal output
flabel metal3 s 15800 11764 15880 11844 0 FreeSans 320 0 0 0 N4BEG[14]
port 129 nsew signal output
flabel metal3 s 16184 11764 16264 11844 0 FreeSans 320 0 0 0 N4BEG[15]
port 130 nsew signal output
flabel metal3 s 10808 11764 10888 11844 0 FreeSans 320 0 0 0 N4BEG[1]
port 131 nsew signal output
flabel metal3 s 11192 11764 11272 11844 0 FreeSans 320 0 0 0 N4BEG[2]
port 132 nsew signal output
flabel metal3 s 11576 11764 11656 11844 0 FreeSans 320 0 0 0 N4BEG[3]
port 133 nsew signal output
flabel metal3 s 11960 11764 12040 11844 0 FreeSans 320 0 0 0 N4BEG[4]
port 134 nsew signal output
flabel metal3 s 12344 11764 12424 11844 0 FreeSans 320 0 0 0 N4BEG[5]
port 135 nsew signal output
flabel metal3 s 12728 11764 12808 11844 0 FreeSans 320 0 0 0 N4BEG[6]
port 136 nsew signal output
flabel metal3 s 13112 11764 13192 11844 0 FreeSans 320 0 0 0 N4BEG[7]
port 137 nsew signal output
flabel metal3 s 13496 11764 13576 11844 0 FreeSans 320 0 0 0 N4BEG[8]
port 138 nsew signal output
flabel metal3 s 13880 11764 13960 11844 0 FreeSans 320 0 0 0 N4BEG[9]
port 139 nsew signal output
flabel metal3 s 16568 11764 16648 11844 0 FreeSans 320 0 0 0 NN4BEG[0]
port 140 nsew signal output
flabel metal3 s 20408 11764 20488 11844 0 FreeSans 320 0 0 0 NN4BEG[10]
port 141 nsew signal output
flabel metal3 s 20792 11764 20872 11844 0 FreeSans 320 0 0 0 NN4BEG[11]
port 142 nsew signal output
flabel metal3 s 21176 11764 21256 11844 0 FreeSans 320 0 0 0 NN4BEG[12]
port 143 nsew signal output
flabel metal3 s 21560 11764 21640 11844 0 FreeSans 320 0 0 0 NN4BEG[13]
port 144 nsew signal output
flabel metal3 s 21944 11764 22024 11844 0 FreeSans 320 0 0 0 NN4BEG[14]
port 145 nsew signal output
flabel metal3 s 22328 11764 22408 11844 0 FreeSans 320 0 0 0 NN4BEG[15]
port 146 nsew signal output
flabel metal3 s 16952 11764 17032 11844 0 FreeSans 320 0 0 0 NN4BEG[1]
port 147 nsew signal output
flabel metal3 s 17336 11764 17416 11844 0 FreeSans 320 0 0 0 NN4BEG[2]
port 148 nsew signal output
flabel metal3 s 17720 11764 17800 11844 0 FreeSans 320 0 0 0 NN4BEG[3]
port 149 nsew signal output
flabel metal3 s 18104 11764 18184 11844 0 FreeSans 320 0 0 0 NN4BEG[4]
port 150 nsew signal output
flabel metal3 s 18488 11764 18568 11844 0 FreeSans 320 0 0 0 NN4BEG[5]
port 151 nsew signal output
flabel metal3 s 18872 11764 18952 11844 0 FreeSans 320 0 0 0 NN4BEG[6]
port 152 nsew signal output
flabel metal3 s 19256 11764 19336 11844 0 FreeSans 320 0 0 0 NN4BEG[7]
port 153 nsew signal output
flabel metal3 s 19640 11764 19720 11844 0 FreeSans 320 0 0 0 NN4BEG[8]
port 154 nsew signal output
flabel metal3 s 20024 11764 20104 11844 0 FreeSans 320 0 0 0 NN4BEG[9]
port 155 nsew signal output
flabel metal3 s 22712 11764 22792 11844 0 FreeSans 320 0 0 0 S1END[0]
port 156 nsew signal input
flabel metal3 s 23096 11764 23176 11844 0 FreeSans 320 0 0 0 S1END[1]
port 157 nsew signal input
flabel metal3 s 23480 11764 23560 11844 0 FreeSans 320 0 0 0 S1END[2]
port 158 nsew signal input
flabel metal3 s 23864 11764 23944 11844 0 FreeSans 320 0 0 0 S1END[3]
port 159 nsew signal input
flabel metal3 s 27320 11764 27400 11844 0 FreeSans 320 0 0 0 S2END[0]
port 160 nsew signal input
flabel metal3 s 27704 11764 27784 11844 0 FreeSans 320 0 0 0 S2END[1]
port 161 nsew signal input
flabel metal3 s 28088 11764 28168 11844 0 FreeSans 320 0 0 0 S2END[2]
port 162 nsew signal input
flabel metal3 s 28472 11764 28552 11844 0 FreeSans 320 0 0 0 S2END[3]
port 163 nsew signal input
flabel metal3 s 28856 11764 28936 11844 0 FreeSans 320 0 0 0 S2END[4]
port 164 nsew signal input
flabel metal3 s 29240 11764 29320 11844 0 FreeSans 320 0 0 0 S2END[5]
port 165 nsew signal input
flabel metal3 s 29624 11764 29704 11844 0 FreeSans 320 0 0 0 S2END[6]
port 166 nsew signal input
flabel metal3 s 30008 11764 30088 11844 0 FreeSans 320 0 0 0 S2END[7]
port 167 nsew signal input
flabel metal3 s 24248 11764 24328 11844 0 FreeSans 320 0 0 0 S2MID[0]
port 168 nsew signal input
flabel metal3 s 24632 11764 24712 11844 0 FreeSans 320 0 0 0 S2MID[1]
port 169 nsew signal input
flabel metal3 s 25016 11764 25096 11844 0 FreeSans 320 0 0 0 S2MID[2]
port 170 nsew signal input
flabel metal3 s 25400 11764 25480 11844 0 FreeSans 320 0 0 0 S2MID[3]
port 171 nsew signal input
flabel metal3 s 25784 11764 25864 11844 0 FreeSans 320 0 0 0 S2MID[4]
port 172 nsew signal input
flabel metal3 s 26168 11764 26248 11844 0 FreeSans 320 0 0 0 S2MID[5]
port 173 nsew signal input
flabel metal3 s 26552 11764 26632 11844 0 FreeSans 320 0 0 0 S2MID[6]
port 174 nsew signal input
flabel metal3 s 26936 11764 27016 11844 0 FreeSans 320 0 0 0 S2MID[7]
port 175 nsew signal input
flabel metal3 s 30392 11764 30472 11844 0 FreeSans 320 0 0 0 S4END[0]
port 176 nsew signal input
flabel metal3 s 34232 11764 34312 11844 0 FreeSans 320 0 0 0 S4END[10]
port 177 nsew signal input
flabel metal3 s 34616 11764 34696 11844 0 FreeSans 320 0 0 0 S4END[11]
port 178 nsew signal input
flabel metal3 s 35000 11764 35080 11844 0 FreeSans 320 0 0 0 S4END[12]
port 179 nsew signal input
flabel metal3 s 35384 11764 35464 11844 0 FreeSans 320 0 0 0 S4END[13]
port 180 nsew signal input
flabel metal3 s 35768 11764 35848 11844 0 FreeSans 320 0 0 0 S4END[14]
port 181 nsew signal input
flabel metal3 s 36152 11764 36232 11844 0 FreeSans 320 0 0 0 S4END[15]
port 182 nsew signal input
flabel metal3 s 30776 11764 30856 11844 0 FreeSans 320 0 0 0 S4END[1]
port 183 nsew signal input
flabel metal3 s 31160 11764 31240 11844 0 FreeSans 320 0 0 0 S4END[2]
port 184 nsew signal input
flabel metal3 s 31544 11764 31624 11844 0 FreeSans 320 0 0 0 S4END[3]
port 185 nsew signal input
flabel metal3 s 31928 11764 32008 11844 0 FreeSans 320 0 0 0 S4END[4]
port 186 nsew signal input
flabel metal3 s 32312 11764 32392 11844 0 FreeSans 320 0 0 0 S4END[5]
port 187 nsew signal input
flabel metal3 s 32696 11764 32776 11844 0 FreeSans 320 0 0 0 S4END[6]
port 188 nsew signal input
flabel metal3 s 33080 11764 33160 11844 0 FreeSans 320 0 0 0 S4END[7]
port 189 nsew signal input
flabel metal3 s 33464 11764 33544 11844 0 FreeSans 320 0 0 0 S4END[8]
port 190 nsew signal input
flabel metal3 s 33848 11764 33928 11844 0 FreeSans 320 0 0 0 S4END[9]
port 191 nsew signal input
flabel metal3 s 36536 11764 36616 11844 0 FreeSans 320 0 0 0 SS4END[0]
port 192 nsew signal input
flabel metal3 s 40376 11764 40456 11844 0 FreeSans 320 0 0 0 SS4END[10]
port 193 nsew signal input
flabel metal3 s 40760 11764 40840 11844 0 FreeSans 320 0 0 0 SS4END[11]
port 194 nsew signal input
flabel metal3 s 41144 11764 41224 11844 0 FreeSans 320 0 0 0 SS4END[12]
port 195 nsew signal input
flabel metal3 s 41528 11764 41608 11844 0 FreeSans 320 0 0 0 SS4END[13]
port 196 nsew signal input
flabel metal3 s 41912 11764 41992 11844 0 FreeSans 320 0 0 0 SS4END[14]
port 197 nsew signal input
flabel metal3 s 42296 11764 42376 11844 0 FreeSans 320 0 0 0 SS4END[15]
port 198 nsew signal input
flabel metal3 s 36920 11764 37000 11844 0 FreeSans 320 0 0 0 SS4END[1]
port 199 nsew signal input
flabel metal3 s 37304 11764 37384 11844 0 FreeSans 320 0 0 0 SS4END[2]
port 200 nsew signal input
flabel metal3 s 37688 11764 37768 11844 0 FreeSans 320 0 0 0 SS4END[3]
port 201 nsew signal input
flabel metal3 s 38072 11764 38152 11844 0 FreeSans 320 0 0 0 SS4END[4]
port 202 nsew signal input
flabel metal3 s 38456 11764 38536 11844 0 FreeSans 320 0 0 0 SS4END[5]
port 203 nsew signal input
flabel metal3 s 38840 11764 38920 11844 0 FreeSans 320 0 0 0 SS4END[6]
port 204 nsew signal input
flabel metal3 s 39224 11764 39304 11844 0 FreeSans 320 0 0 0 SS4END[7]
port 205 nsew signal input
flabel metal3 s 39608 11764 39688 11844 0 FreeSans 320 0 0 0 SS4END[8]
port 206 nsew signal input
flabel metal3 s 39992 11764 40072 11844 0 FreeSans 320 0 0 0 SS4END[9]
port 207 nsew signal input
flabel metal3 s 1592 0 1672 80 0 FreeSans 320 0 0 0 UserCLK
port 208 nsew signal input
flabel metal3 s 42680 11764 42760 11844 0 FreeSans 320 0 0 0 UserCLKo
port 209 nsew signal output
flabel metal5 s 4892 0 5332 11844 0 FreeSans 2560 90 0 0 VGND
port 210 nsew ground bidirectional
flabel metal5 s 4892 0 5332 40 0 FreeSans 320 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal5 s 4892 11804 5332 11844 0 FreeSans 320 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal5 s 20012 0 20452 11844 0 FreeSans 2560 90 0 0 VGND
port 210 nsew ground bidirectional
flabel metal5 s 20012 0 20452 40 0 FreeSans 320 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal5 s 20012 11804 20452 11844 0 FreeSans 320 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal5 s 35132 0 35572 11844 0 FreeSans 2560 90 0 0 VGND
port 210 nsew ground bidirectional
flabel metal5 s 35132 0 35572 40 0 FreeSans 320 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal5 s 35132 11804 35572 11844 0 FreeSans 320 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal5 s 50252 0 50692 11844 0 FreeSans 2560 90 0 0 VGND
port 210 nsew ground bidirectional
flabel metal5 s 50252 0 50692 40 0 FreeSans 320 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal5 s 50252 11804 50692 11844 0 FreeSans 320 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal5 s 3652 0 4092 11844 0 FreeSans 2560 90 0 0 VPWR
port 211 nsew power bidirectional
flabel metal5 s 3652 0 4092 40 0 FreeSans 320 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal5 s 3652 11804 4092 11844 0 FreeSans 320 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal5 s 18772 0 19212 11844 0 FreeSans 2560 90 0 0 VPWR
port 211 nsew power bidirectional
flabel metal5 s 18772 0 19212 40 0 FreeSans 320 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal5 s 18772 11804 19212 11844 0 FreeSans 320 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal5 s 33892 0 34332 11844 0 FreeSans 2560 90 0 0 VPWR
port 211 nsew power bidirectional
flabel metal5 s 33892 0 34332 40 0 FreeSans 320 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal5 s 33892 11804 34332 11844 0 FreeSans 320 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal5 s 49012 0 49452 11844 0 FreeSans 2560 90 0 0 VPWR
port 211 nsew power bidirectional
flabel metal5 s 49012 0 49452 40 0 FreeSans 320 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal5 s 49012 11804 49452 11844 0 FreeSans 320 0 0 0 VPWR
port 211 nsew power bidirectional
rlabel metal1 26640 9072 26640 9072 0 VGND
rlabel metal1 26640 9828 26640 9828 0 VPWR
rlabel metal2 9008 588 9008 588 0 FrameData[0]
rlabel metal2 22272 3318 22272 3318 0 FrameData[10]
rlabel metal2 24480 4200 24480 4200 0 FrameData[11]
rlabel metal3 22368 3990 22368 3990 0 FrameData[12]
rlabel metal3 21600 4242 21600 4242 0 FrameData[13]
rlabel metal2 80 5292 80 5292 0 FrameData[14]
rlabel metal2 128 5628 128 5628 0 FrameData[15]
rlabel metal2 560 5964 560 5964 0 FrameData[16]
rlabel metal2 752 6300 752 6300 0 FrameData[17]
rlabel metal2 512 6636 512 6636 0 FrameData[18]
rlabel metal2 368 6972 368 6972 0 FrameData[19]
rlabel metal2 9104 924 9104 924 0 FrameData[1]
rlabel metal2 608 7308 608 7308 0 FrameData[20]
rlabel metal2 18720 7182 18720 7182 0 FrameData[21]
rlabel metal2 656 7980 656 7980 0 FrameData[22]
rlabel metal2 128 8316 128 8316 0 FrameData[23]
rlabel metal2 752 8652 752 8652 0 FrameData[24]
rlabel metal3 17472 8862 17472 8862 0 FrameData[25]
rlabel metal2 176 9324 176 9324 0 FrameData[26]
rlabel metal2 1040 9660 1040 9660 0 FrameData[27]
rlabel metal2 752 9996 752 9996 0 FrameData[28]
rlabel metal2 656 10332 656 10332 0 FrameData[29]
rlabel metal2 9200 1260 9200 1260 0 FrameData[2]
rlabel metal2 320 10668 320 10668 0 FrameData[30]
rlabel metal2 416 11004 416 11004 0 FrameData[31]
rlabel metal2 9968 1596 9968 1596 0 FrameData[3]
rlabel metal2 9776 1932 9776 1932 0 FrameData[4]
rlabel metal2 128 2268 128 2268 0 FrameData[5]
rlabel metal2 80 2604 80 2604 0 FrameData[6]
rlabel metal3 24096 3528 24096 3528 0 FrameData[7]
rlabel metal2 22176 3234 22176 3234 0 FrameData[8]
rlabel metal2 22080 3990 22080 3990 0 FrameData[9]
rlabel metal2 52767 588 52767 588 0 FrameData_O[0]
rlabel metal2 52911 3948 52911 3948 0 FrameData_O[10]
rlabel metal2 52647 4284 52647 4284 0 FrameData_O[11]
rlabel metal2 52455 4620 52455 4620 0 FrameData_O[12]
rlabel metal2 52647 4956 52647 4956 0 FrameData_O[13]
rlabel metal2 53151 5292 53151 5292 0 FrameData_O[14]
rlabel metal2 52647 5628 52647 5628 0 FrameData_O[15]
rlabel metal2 53151 5964 53151 5964 0 FrameData_O[16]
rlabel metal2 52647 6300 52647 6300 0 FrameData_O[17]
rlabel metal2 52455 6636 52455 6636 0 FrameData_O[18]
rlabel metal2 52647 6972 52647 6972 0 FrameData_O[19]
rlabel metal2 53103 924 53103 924 0 FrameData_O[1]
rlabel metal2 52959 7308 52959 7308 0 FrameData_O[20]
rlabel metal2 52455 7644 52455 7644 0 FrameData_O[21]
rlabel metal2 52959 7980 52959 7980 0 FrameData_O[22]
rlabel metal2 52575 8316 52575 8316 0 FrameData_O[23]
rlabel metal2 52959 8652 52959 8652 0 FrameData_O[24]
rlabel metal2 53199 8988 53199 8988 0 FrameData_O[25]
rlabel metal2 52263 9324 52263 9324 0 FrameData_O[26]
rlabel metal2 51240 8904 51240 8904 0 FrameData_O[27]
rlabel metal2 51000 8904 51000 8904 0 FrameData_O[28]
rlabel metal2 51816 8148 51816 8148 0 FrameData_O[29]
rlabel via2 53199 1260 53199 1260 0 FrameData_O[2]
rlabel metal2 50664 8904 50664 8904 0 FrameData_O[30]
rlabel metal2 50136 8904 50136 8904 0 FrameData_O[31]
rlabel metal2 52455 1596 52455 1596 0 FrameData_O[3]
rlabel metal2 52575 1932 52575 1932 0 FrameData_O[4]
rlabel metal2 52296 2100 52296 2100 0 FrameData_O[5]
rlabel metal2 52911 2604 52911 2604 0 FrameData_O[6]
rlabel metal2 52392 2856 52392 2856 0 FrameData_O[7]
rlabel metal2 52455 3276 52455 3276 0 FrameData_O[8]
rlabel metal2 52647 3612 52647 3612 0 FrameData_O[9]
rlabel metal2 17952 6426 17952 6426 0 FrameStrobe[0]
rlabel metal3 29088 3348 29088 3348 0 FrameStrobe[10]
rlabel metal3 31584 2970 31584 2970 0 FrameStrobe[11]
rlabel via3 34080 72 34080 72 0 FrameStrobe[12]
rlabel metal2 36480 7980 36480 7980 0 FrameStrobe[13]
rlabel metal2 37920 7560 37920 7560 0 FrameStrobe[14]
rlabel metal2 40608 6468 40608 6468 0 FrameStrobe[15]
rlabel metal2 43200 6468 43200 6468 0 FrameStrobe[16]
rlabel metal2 46512 5628 46512 5628 0 FrameStrobe[17]
rlabel metal3 49056 744 49056 744 0 FrameStrobe[18]
rlabel metal2 50400 5712 50400 5712 0 FrameStrobe[19]
rlabel metal3 6624 3180 6624 3180 0 FrameStrobe[1]
rlabel metal3 9120 3138 9120 3138 0 FrameStrobe[2]
rlabel metal3 11616 3096 11616 3096 0 FrameStrobe[3]
rlabel metal3 14112 2634 14112 2634 0 FrameStrobe[4]
rlabel metal3 16608 2718 16608 2718 0 FrameStrobe[5]
rlabel metal3 19104 114 19104 114 0 FrameStrobe[6]
rlabel metal3 21600 954 21600 954 0 FrameStrobe[7]
rlabel metal3 33312 5460 33312 5460 0 FrameStrobe[8]
rlabel metal2 34848 6300 34848 6300 0 FrameStrobe[9]
rlabel metal2 43128 9660 43128 9660 0 FrameStrobe_O[0]
rlabel metal2 46968 9660 46968 9660 0 FrameStrobe_O[10]
rlabel metal2 47352 9660 47352 9660 0 FrameStrobe_O[11]
rlabel metal2 47736 9660 47736 9660 0 FrameStrobe_O[12]
rlabel metal2 48120 9660 48120 9660 0 FrameStrobe_O[13]
rlabel metal2 48504 9660 48504 9660 0 FrameStrobe_O[14]
rlabel metal2 48888 9660 48888 9660 0 FrameStrobe_O[15]
rlabel metal2 49416 9660 49416 9660 0 FrameStrobe_O[16]
rlabel metal2 49656 9576 49656 9576 0 FrameStrobe_O[17]
rlabel metal2 50040 9660 50040 9660 0 FrameStrobe_O[18]
rlabel metal2 50424 9660 50424 9660 0 FrameStrobe_O[19]
rlabel metal2 43512 9660 43512 9660 0 FrameStrobe_O[1]
rlabel metal2 43896 9660 43896 9660 0 FrameStrobe_O[2]
rlabel metal2 44280 9660 44280 9660 0 FrameStrobe_O[3]
rlabel metal2 44664 9660 44664 9660 0 FrameStrobe_O[4]
rlabel metal2 45048 9660 45048 9660 0 FrameStrobe_O[5]
rlabel metal2 45432 9660 45432 9660 0 FrameStrobe_O[6]
rlabel metal2 45816 9660 45816 9660 0 FrameStrobe_O[7]
rlabel metal2 46200 9660 46200 9660 0 FrameStrobe_O[8]
rlabel metal2 46584 9660 46584 9660 0 FrameStrobe_O[9]
rlabel metal2 2808 9660 2808 9660 0 N1BEG[0]
rlabel metal2 3192 9660 3192 9660 0 N1BEG[1]
rlabel metal2 3576 9660 3576 9660 0 N1BEG[2]
rlabel metal2 4056 9660 4056 9660 0 N1BEG[3]
rlabel metal2 4344 9660 4344 9660 0 N2BEG[0]
rlabel metal2 4728 9660 4728 9660 0 N2BEG[1]
rlabel metal2 5112 9660 5112 9660 0 N2BEG[2]
rlabel metal2 5496 9660 5496 9660 0 N2BEG[3]
rlabel metal2 5880 9660 5880 9660 0 N2BEG[4]
rlabel metal2 6264 9660 6264 9660 0 N2BEG[5]
rlabel metal2 6648 9660 6648 9660 0 N2BEG[6]
rlabel metal2 7032 9660 7032 9660 0 N2BEG[7]
rlabel metal2 7416 9660 7416 9660 0 N2BEGb[0]
rlabel metal2 7800 9660 7800 9660 0 N2BEGb[1]
rlabel metal2 8184 9660 8184 9660 0 N2BEGb[2]
rlabel metal2 8568 9660 8568 9660 0 N2BEGb[3]
rlabel metal2 8952 9660 8952 9660 0 N2BEGb[4]
rlabel metal2 9336 9660 9336 9660 0 N2BEGb[5]
rlabel metal2 9720 9660 9720 9660 0 N2BEGb[6]
rlabel metal2 10104 9660 10104 9660 0 N2BEGb[7]
rlabel metal2 10488 9660 10488 9660 0 N4BEG[0]
rlabel metal2 14328 9660 14328 9660 0 N4BEG[10]
rlabel metal2 14712 9660 14712 9660 0 N4BEG[11]
rlabel metal2 15096 9660 15096 9660 0 N4BEG[12]
rlabel metal2 15480 9660 15480 9660 0 N4BEG[13]
rlabel metal2 15864 9660 15864 9660 0 N4BEG[14]
rlabel metal2 16248 9660 16248 9660 0 N4BEG[15]
rlabel metal2 10872 9660 10872 9660 0 N4BEG[1]
rlabel metal2 11256 9660 11256 9660 0 N4BEG[2]
rlabel metal2 11640 9660 11640 9660 0 N4BEG[3]
rlabel metal2 12024 9660 12024 9660 0 N4BEG[4]
rlabel metal2 12408 9660 12408 9660 0 N4BEG[5]
rlabel metal2 12792 9660 12792 9660 0 N4BEG[6]
rlabel metal2 13176 9660 13176 9660 0 N4BEG[7]
rlabel metal2 13560 9660 13560 9660 0 N4BEG[8]
rlabel metal2 13944 9660 13944 9660 0 N4BEG[9]
rlabel metal2 16632 9660 16632 9660 0 NN4BEG[0]
rlabel metal2 20472 9660 20472 9660 0 NN4BEG[10]
rlabel metal2 20856 9660 20856 9660 0 NN4BEG[11]
rlabel metal2 21240 9660 21240 9660 0 NN4BEG[12]
rlabel metal2 21624 9660 21624 9660 0 NN4BEG[13]
rlabel metal2 22008 9660 22008 9660 0 NN4BEG[14]
rlabel metal2 22392 9660 22392 9660 0 NN4BEG[15]
rlabel metal2 17016 9660 17016 9660 0 NN4BEG[1]
rlabel metal2 17400 9660 17400 9660 0 NN4BEG[2]
rlabel metal2 17784 9660 17784 9660 0 NN4BEG[3]
rlabel metal2 18168 9660 18168 9660 0 NN4BEG[4]
rlabel metal2 18552 9660 18552 9660 0 NN4BEG[5]
rlabel metal2 18840 9576 18840 9576 0 NN4BEG[6]
rlabel metal2 19320 9660 19320 9660 0 NN4BEG[7]
rlabel metal2 19704 9660 19704 9660 0 NN4BEG[8]
rlabel metal2 20088 9660 20088 9660 0 NN4BEG[9]
rlabel metal3 22752 10848 22752 10848 0 S1END[0]
rlabel metal2 20256 7770 20256 7770 0 S1END[1]
rlabel metal2 9984 8190 9984 8190 0 S1END[2]
rlabel metal3 20928 8610 20928 8610 0 S1END[3]
rlabel metal3 11136 6468 11136 6468 0 S2END[0]
rlabel metal3 19344 6636 19344 6636 0 S2END[1]
rlabel metal2 13632 6972 13632 6972 0 S2END[2]
rlabel metal3 15264 6216 15264 6216 0 S2END[3]
rlabel metal2 19296 6678 19296 6678 0 S2END[4]
rlabel metal2 20640 6510 20640 6510 0 S2END[5]
rlabel metal3 22752 7854 22752 7854 0 S2END[6]
rlabel metal2 20160 7854 20160 7854 0 S2END[7]
rlabel metal2 15264 7392 15264 7392 0 S2MID[0]
rlabel metal3 18048 9408 18048 9408 0 S2MID[1]
rlabel metal2 8064 7938 8064 7938 0 S2MID[2]
rlabel metal3 14400 8946 14400 8946 0 S2MID[3]
rlabel metal3 15360 8232 15360 8232 0 S2MID[4]
rlabel metal2 14016 7098 14016 7098 0 S2MID[5]
rlabel metal3 17040 6972 17040 6972 0 S2MID[6]
rlabel metal2 22944 7350 22944 7350 0 S2MID[7]
rlabel metal3 19296 7602 19296 7602 0 S4END[0]
rlabel metal3 21024 8694 21024 8694 0 S4END[10]
rlabel metal3 22656 9282 22656 9282 0 S4END[11]
rlabel metal2 22368 8694 22368 8694 0 S4END[12]
rlabel metal3 22752 8904 22752 8904 0 S4END[13]
rlabel metal3 35808 10932 35808 10932 0 S4END[14]
rlabel metal3 36192 10722 36192 10722 0 S4END[15]
rlabel metal3 19872 9954 19872 9954 0 S4END[1]
rlabel metal3 19584 10584 19584 10584 0 S4END[2]
rlabel metal3 17280 9912 17280 9912 0 S4END[3]
rlabel metal3 17184 9450 17184 9450 0 S4END[4]
rlabel metal2 20064 8064 20064 8064 0 S4END[5]
rlabel metal3 19392 9660 19392 9660 0 S4END[6]
rlabel metal3 18624 8274 18624 8274 0 S4END[7]
rlabel metal2 19680 8148 19680 8148 0 S4END[8]
rlabel metal2 20544 8022 20544 8022 0 S4END[9]
rlabel metal3 36576 9966 36576 9966 0 SS4END[0]
rlabel metal3 40416 10176 40416 10176 0 SS4END[10]
rlabel metal3 40800 9588 40800 9588 0 SS4END[11]
rlabel metal3 41184 9630 41184 9630 0 SS4END[12]
rlabel metal3 41568 10050 41568 10050 0 SS4END[13]
rlabel metal3 41952 9924 41952 9924 0 SS4END[14]
rlabel metal3 42336 10428 42336 10428 0 SS4END[15]
rlabel metal3 36960 10848 36960 10848 0 SS4END[1]
rlabel metal4 37872 9072 37872 9072 0 SS4END[2]
rlabel metal3 37728 10050 37728 10050 0 SS4END[3]
rlabel metal4 38736 7224 38736 7224 0 SS4END[4]
rlabel metal3 38496 9798 38496 9798 0 SS4END[5]
rlabel metal3 38880 9966 38880 9966 0 SS4END[6]
rlabel metal3 39264 9924 39264 9924 0 SS4END[7]
rlabel metal3 39648 10092 39648 10092 0 SS4END[8]
rlabel metal3 40032 10134 40032 10134 0 SS4END[9]
rlabel metal3 1632 2844 1632 2844 0 UserCLK
rlabel metal2 42744 9660 42744 9660 0 UserCLKo
rlabel metal2 21192 3948 21192 3948 0 net1
rlabel metal4 38256 7140 38256 7140 0 net10
rlabel metal2 19104 9618 19104 9618 0 net100
rlabel metal3 22176 9282 22176 9282 0 net101
rlabel metal2 19584 9534 19584 9534 0 net102
rlabel metal3 19968 9324 19968 9324 0 net103
rlabel metal2 39432 8064 39432 8064 0 net104
rlabel metal3 40320 7518 40320 7518 0 net105
rlabel metal3 38112 5460 38112 5460 0 net11
rlabel metal3 22944 3414 22944 3414 0 net12
rlabel metal3 27936 6384 27936 6384 0 net13
rlabel metal3 27552 6468 27552 6468 0 net14
rlabel metal2 38112 6762 38112 6762 0 net15
rlabel metal4 30048 8694 30048 8694 0 net16
rlabel metal3 47136 9282 47136 9282 0 net17
rlabel metal2 29256 8904 29256 8904 0 net18
rlabel metal2 28632 8064 28632 8064 0 net19
rlabel metal2 51456 4074 51456 4074 0 net2
rlabel metal2 28584 8652 28584 8652 0 net20
rlabel metal2 28800 8820 28800 8820 0 net21
rlabel metal2 38976 7266 38976 7266 0 net22
rlabel metal2 24816 2184 24816 2184 0 net23
rlabel metal2 27768 8652 27768 8652 0 net24
rlabel metal4 34752 8904 34752 8904 0 net25
rlabel metal2 50400 2058 50400 2058 0 net26
rlabel metal2 21912 3948 21912 3948 0 net27
rlabel metal2 49536 2226 49536 2226 0 net28
rlabel metal2 51456 2688 51456 2688 0 net29
rlabel metal2 25344 3906 25344 3906 0 net3
rlabel metal2 51168 2604 51168 2604 0 net30
rlabel metal2 31296 4200 31296 4200 0 net31
rlabel metal2 24960 4116 24960 4116 0 net32
rlabel metal3 34896 6384 34896 6384 0 net33
rlabel metal3 47232 8190 47232 8190 0 net34
rlabel metal3 41184 7014 41184 7014 0 net35
rlabel metal2 38472 8148 38472 8148 0 net36
rlabel metal2 36960 7686 36960 7686 0 net37
rlabel metal3 39744 7812 39744 7812 0 net38
rlabel metal3 48960 7560 48960 7560 0 net39
rlabel metal2 25512 3612 25512 3612 0 net4
rlabel metal2 42600 6552 42600 6552 0 net40
rlabel metal2 46728 5628 46728 5628 0 net41
rlabel metal2 49848 6636 49848 6636 0 net42
rlabel metal2 49752 5628 49752 5628 0 net43
rlabel metal4 34944 6216 34944 6216 0 net44
rlabel metal2 38112 6594 38112 6594 0 net45
rlabel metal2 24504 6636 24504 6636 0 net46
rlabel metal3 33216 5292 33216 5292 0 net47
rlabel metal2 35424 5670 35424 5670 0 net48
rlabel metal3 41856 7098 41856 7098 0 net49
rlabel metal2 24648 3612 24648 3612 0 net5
rlabel metal3 46080 7098 46080 7098 0 net50
rlabel metal3 46464 7476 46464 7476 0 net51
rlabel metal3 46848 7896 46848 7896 0 net52
rlabel metal2 10632 7980 10632 7980 0 net53
rlabel metal2 7704 7812 7704 7812 0 net54
rlabel metal2 4344 8148 4344 8148 0 net55
rlabel metal2 3816 8148 3816 8148 0 net56
rlabel metal3 4608 9366 4608 9366 0 net57
rlabel metal2 15048 7140 15048 7140 0 net58
rlabel metal2 13752 6972 13752 6972 0 net59
rlabel metal2 22056 3612 22056 3612 0 net6
rlabel metal2 11736 8064 11736 8064 0 net60
rlabel metal2 10200 8148 10200 8148 0 net61
rlabel metal2 7800 8148 7800 8148 0 net62
rlabel metal2 6648 8148 6648 8148 0 net63
rlabel metal2 6312 8064 6312 8064 0 net64
rlabel metal2 16056 8148 16056 8148 0 net65
rlabel metal2 14184 8148 14184 8148 0 net66
rlabel metal3 14112 6762 14112 6762 0 net67
rlabel metal2 13176 6972 13176 6972 0 net68
rlabel metal2 12168 6972 12168 6972 0 net69
rlabel metal2 23448 3612 23448 3612 0 net7
rlabel metal2 10680 6972 10680 6972 0 net70
rlabel metal2 10632 7056 10632 7056 0 net71
rlabel metal2 10632 7140 10632 7140 0 net72
rlabel metal2 22848 10122 22848 10122 0 net73
rlabel metal2 16824 8148 16824 8148 0 net74
rlabel metal2 16056 6972 16056 6972 0 net75
rlabel metal2 16440 8148 16440 8148 0 net76
rlabel metal2 17160 8064 17160 8064 0 net77
rlabel metal2 17976 8148 17976 8148 0 net78
rlabel metal2 18888 8148 18888 8148 0 net79
rlabel metal2 25608 2856 25608 2856 0 net8
rlabel metal3 22848 9408 22848 9408 0 net80
rlabel metal2 22488 8484 22488 8484 0 net81
rlabel metal2 19968 9030 19968 9030 0 net82
rlabel metal2 17760 8862 17760 8862 0 net83
rlabel metal3 12672 9072 12672 9072 0 net84
rlabel metal3 13248 9114 13248 9114 0 net85
rlabel metal2 18936 8064 18936 8064 0 net86
rlabel metal2 18360 8148 18360 8148 0 net87
rlabel metal2 17592 8148 17592 8148 0 net88
rlabel metal2 16896 9366 16896 9366 0 net89
rlabel metal2 34944 6216 34944 6216 0 net9
rlabel metal3 21792 8652 21792 8652 0 net90
rlabel metal3 21600 8190 21600 8190 0 net91
rlabel metal3 21696 8652 21696 8652 0 net92
rlabel metal2 21888 9534 21888 9534 0 net93
rlabel metal2 37032 8148 37032 8148 0 net94
rlabel metal3 33312 7686 33312 7686 0 net95
rlabel metal4 18576 9408 18576 9408 0 net96
rlabel metal3 20064 8610 20064 8610 0 net97
rlabel metal3 19680 8316 19680 8316 0 net98
rlabel metal3 22560 7518 22560 7518 0 net99
<< properties >>
string FIXED_BBOX 0 0 53280 11844
<< end >>
