* NGSPICE file created from S_term_single2.ext - technology: ihp-sg13g2

* Black-box entry subcircuit for sg13g2_decap_8 abstract view
.subckt sg13g2_decap_8 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_1 abstract view
.subckt sg13g2_buf_1 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_1 abstract view
.subckt sg13g2_fill_1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_decap_4 abstract view
.subckt sg13g2_decap_4 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_2 abstract view
.subckt sg13g2_fill_2 VDD VSS
.ends

.subckt S_term_single2 FrameData[0] FrameData[10] FrameData[11] FrameData[12] FrameData[13]
+ FrameData[14] FrameData[15] FrameData[16] FrameData[17] FrameData[18] FrameData[19]
+ FrameData[1] FrameData[20] FrameData[21] FrameData[22] FrameData[23] FrameData[24]
+ FrameData[25] FrameData[26] FrameData[27] FrameData[28] FrameData[29] FrameData[2]
+ FrameData[30] FrameData[31] FrameData[3] FrameData[4] FrameData[5] FrameData[6]
+ FrameData[7] FrameData[8] FrameData[9] FrameData_O[0] FrameData_O[10] FrameData_O[11]
+ FrameData_O[12] FrameData_O[13] FrameData_O[14] FrameData_O[15] FrameData_O[16]
+ FrameData_O[17] FrameData_O[18] FrameData_O[19] FrameData_O[1] FrameData_O[20] FrameData_O[21]
+ FrameData_O[22] FrameData_O[23] FrameData_O[24] FrameData_O[25] FrameData_O[26]
+ FrameData_O[27] FrameData_O[28] FrameData_O[29] FrameData_O[2] FrameData_O[30] FrameData_O[31]
+ FrameData_O[3] FrameData_O[4] FrameData_O[5] FrameData_O[6] FrameData_O[7] FrameData_O[8]
+ FrameData_O[9] FrameStrobe[0] FrameStrobe[10] FrameStrobe[11] FrameStrobe[12] FrameStrobe[13]
+ FrameStrobe[14] FrameStrobe[15] FrameStrobe[16] FrameStrobe[17] FrameStrobe[18]
+ FrameStrobe[19] FrameStrobe[1] FrameStrobe[2] FrameStrobe[3] FrameStrobe[4] FrameStrobe[5]
+ FrameStrobe[6] FrameStrobe[7] FrameStrobe[8] FrameStrobe[9] FrameStrobe_O[0] FrameStrobe_O[10]
+ FrameStrobe_O[11] FrameStrobe_O[12] FrameStrobe_O[13] FrameStrobe_O[14] FrameStrobe_O[15]
+ FrameStrobe_O[16] FrameStrobe_O[17] FrameStrobe_O[18] FrameStrobe_O[19] FrameStrobe_O[1]
+ FrameStrobe_O[2] FrameStrobe_O[3] FrameStrobe_O[4] FrameStrobe_O[5] FrameStrobe_O[6]
+ FrameStrobe_O[7] FrameStrobe_O[8] FrameStrobe_O[9] N1BEG[0] N1BEG[1] N1BEG[2] N1BEG[3]
+ N2BEG[0] N2BEG[1] N2BEG[2] N2BEG[3] N2BEG[4] N2BEG[5] N2BEG[6] N2BEG[7] N2BEGb[0]
+ N2BEGb[1] N2BEGb[2] N2BEGb[3] N2BEGb[4] N2BEGb[5] N2BEGb[6] N2BEGb[7] N4BEG[0] N4BEG[10]
+ N4BEG[11] N4BEG[12] N4BEG[13] N4BEG[14] N4BEG[15] N4BEG[1] N4BEG[2] N4BEG[3] N4BEG[4]
+ N4BEG[5] N4BEG[6] N4BEG[7] N4BEG[8] N4BEG[9] NN4BEG[0] NN4BEG[10] NN4BEG[11] NN4BEG[12]
+ NN4BEG[13] NN4BEG[14] NN4BEG[15] NN4BEG[1] NN4BEG[2] NN4BEG[3] NN4BEG[4] NN4BEG[5]
+ NN4BEG[6] NN4BEG[7] NN4BEG[8] NN4BEG[9] S1END[0] S1END[1] S1END[2] S1END[3] S2END[0]
+ S2END[1] S2END[2] S2END[3] S2END[4] S2END[5] S2END[6] S2END[7] S2MID[0] S2MID[1]
+ S2MID[2] S2MID[3] S2MID[4] S2MID[5] S2MID[6] S2MID[7] S4END[0] S4END[10] S4END[11]
+ S4END[12] S4END[13] S4END[14] S4END[15] S4END[1] S4END[2] S4END[3] S4END[4] S4END[5]
+ S4END[6] S4END[7] S4END[8] S4END[9] SS4END[0] SS4END[10] SS4END[11] SS4END[12] SS4END[13]
+ SS4END[14] SS4END[15] SS4END[1] SS4END[2] SS4END[3] SS4END[4] SS4END[5] SS4END[6]
+ SS4END[7] SS4END[8] SS4END[9] UserCLK UserCLKo VGND VPWR
XFILLER_7_7 VPWR VGND sg13g2_decap_8
XFILLER_9_126 VPWR VGND sg13g2_decap_8
XFILLER_5_343 VPWR VGND sg13g2_decap_8
XFILLER_5_321 VPWR VGND sg13g2_decap_8
XFILLER_3_56 VPWR VGND sg13g2_decap_8
XFILLER_2_335 VPWR VGND sg13g2_decap_8
XFILLER_5_140 VPWR VGND sg13g2_decap_8
X_062_ S2MID[1] net63 VPWR VGND sg13g2_buf_1
XFILLER_9_77 VPWR VGND sg13g2_decap_8
XFILLER_6_460 VPWR VGND sg13g2_decap_8
XFILLER_0_35 VPWR VGND sg13g2_decap_8
XFILLER_2_154 VPWR VGND sg13g2_decap_8
X_045_ FrameStrobe[13] net37 VPWR VGND sg13g2_buf_1
XFILLER_7_268 VPWR VGND sg13g2_fill_1
XFILLER_7_224 VPWR VGND sg13g2_decap_8
XFILLER_3_430 VPWR VGND sg13g2_decap_8
XFILLER_0_455 VPWR VGND sg13g2_decap_8
XFILLER_4_238 VPWR VGND sg13g2_decap_8
X_028_ FrameData[28] net21 VPWR VGND sg13g2_buf_1
XFILLER_8_511 VPWR VGND sg13g2_decap_8
XFILLER_6_56 VPWR VGND sg13g2_decap_8
Xoutput20 net20 FrameData_O[27] VPWR VGND sg13g2_buf_1
Xoutput42 net42 FrameStrobe_O[18] VPWR VGND sg13g2_buf_1
Xoutput97 net97 NN4BEG[2] VPWR VGND sg13g2_buf_1
Xoutput75 net75 N4BEG[11] VPWR VGND sg13g2_buf_1
Xoutput86 net86 N4BEG[7] VPWR VGND sg13g2_buf_1
Xoutput64 net64 N2BEG[7] VPWR VGND sg13g2_buf_1
Xoutput53 net53 N1BEG[0] VPWR VGND sg13g2_buf_1
XFILLER_8_341 VPWR VGND sg13g2_decap_8
Xoutput7 net7 FrameData_O[15] VPWR VGND sg13g2_buf_1
XFILLER_0_252 VPWR VGND sg13g2_decap_8
Xoutput31 net31 FrameData_O[8] VPWR VGND sg13g2_buf_1
XFILLER_2_517 VPWR VGND sg13g2_decap_4
XFILLER_9_105 VPWR VGND sg13g2_decap_8
XFILLER_5_399 VPWR VGND sg13g2_decap_8
XFILLER_3_35 VPWR VGND sg13g2_decap_8
XFILLER_6_119 VPWR VGND sg13g2_decap_8
XFILLER_2_314 VPWR VGND sg13g2_decap_8
XFILLER_5_196 VPWR VGND sg13g2_decap_8
XFILLER_1_380 VPWR VGND sg13g2_decap_8
XFILLER_9_56 VPWR VGND sg13g2_decap_8
X_061_ S2MID[2] net62 VPWR VGND sg13g2_buf_1
XFILLER_7_439 VPWR VGND sg13g2_decap_8
XFILLER_0_14 VPWR VGND sg13g2_decap_8
XFILLER_2_133 VPWR VGND sg13g2_decap_8
X_044_ FrameStrobe[12] net36 VPWR VGND sg13g2_buf_1
XFILLER_7_203 VPWR VGND sg13g2_decap_8
XFILLER_3_486 VPWR VGND sg13g2_decap_8
XFILLER_0_434 VPWR VGND sg13g2_decap_8
XFILLER_4_217 VPWR VGND sg13g2_decap_8
X_027_ FrameData[27] net20 VPWR VGND sg13g2_buf_1
XFILLER_6_35 VPWR VGND sg13g2_decap_8
XFILLER_3_283 VPWR VGND sg13g2_decap_8
Xoutput43 net43 FrameStrobe_O[19] VPWR VGND sg13g2_buf_1
Xoutput21 net21 FrameData_O[28] VPWR VGND sg13g2_buf_1
Xoutput98 net98 NN4BEG[3] VPWR VGND sg13g2_buf_1
Xoutput76 net76 N4BEG[12] VPWR VGND sg13g2_buf_1
Xoutput87 net87 N4BEG[8] VPWR VGND sg13g2_buf_1
Xoutput65 net65 N2BEGb[0] VPWR VGND sg13g2_buf_1
Xoutput54 net54 N1BEG[1] VPWR VGND sg13g2_buf_1
Xoutput10 net10 FrameData_O[18] VPWR VGND sg13g2_buf_1
Xoutput8 net8 FrameData_O[16] VPWR VGND sg13g2_buf_1
XFILLER_5_504 VPWR VGND sg13g2_decap_8
XFILLER_0_231 VPWR VGND sg13g2_decap_8
Xoutput32 net32 FrameData_O[9] VPWR VGND sg13g2_buf_1
XFILLER_5_378 VPWR VGND sg13g2_decap_8
XFILLER_8_194 VPWR VGND sg13g2_decap_4
XFILLER_8_183 VPWR VGND sg13g2_fill_2
XFILLER_3_14 VPWR VGND sg13g2_decap_8
XFILLER_5_175 VPWR VGND sg13g2_decap_8
XFILLER_9_492 VPWR VGND sg13g2_decap_8
XFILLER_9_35 VPWR VGND sg13g2_decap_8
X_060_ S2MID[3] net61 VPWR VGND sg13g2_buf_1
XFILLER_7_418 VPWR VGND sg13g2_decap_8
XFILLER_2_112 VPWR VGND sg13g2_decap_8
XFILLER_2_189 VPWR VGND sg13g2_decap_8
XFILLER_6_495 VPWR VGND sg13g2_decap_4
X_043_ FrameStrobe[11] net35 VPWR VGND sg13g2_buf_1
XFILLER_7_259 VPWR VGND sg13g2_decap_8
XFILLER_1_0 VPWR VGND sg13g2_decap_8
XFILLER_3_465 VPWR VGND sg13g2_decap_8
XFILLER_1_91 VPWR VGND sg13g2_decap_8
XFILLER_0_413 VPWR VGND sg13g2_decap_8
X_026_ FrameData[26] net19 VPWR VGND sg13g2_buf_1
XFILLER_6_14 VPWR VGND sg13g2_decap_8
XFILLER_3_262 VPWR VGND sg13g2_decap_8
Xoutput44 net44 FrameStrobe_O[1] VPWR VGND sg13g2_buf_1
Xoutput33 net33 FrameStrobe_O[0] VPWR VGND sg13g2_buf_1
Xoutput99 net99 NN4BEG[4] VPWR VGND sg13g2_buf_1
Xoutput77 net77 N4BEG[13] VPWR VGND sg13g2_buf_1
Xoutput88 net88 N4BEG[9] VPWR VGND sg13g2_buf_1
Xoutput66 net66 N2BEGb[1] VPWR VGND sg13g2_buf_1
Xoutput55 net55 N1BEG[2] VPWR VGND sg13g2_buf_1
Xoutput22 net22 FrameData_O[29] VPWR VGND sg13g2_buf_1
Xoutput11 net11 FrameData_O[19] VPWR VGND sg13g2_buf_1
Xoutput9 net9 FrameData_O[17] VPWR VGND sg13g2_buf_1
XFILLER_0_287 VPWR VGND sg13g2_decap_8
XFILLER_0_210 VPWR VGND sg13g2_decap_8
XFILLER_8_365 VPWR VGND sg13g2_fill_1
X_009_ FrameData[9] net32 VPWR VGND sg13g2_buf_1
XFILLER_10_309 VPWR VGND sg13g2_decap_8
XFILLER_5_357 VPWR VGND sg13g2_decap_8
XFILLER_5_302 VPWR VGND sg13g2_decap_8
XFILLER_5_7 VPWR VGND sg13g2_decap_8
XFILLER_5_154 VPWR VGND sg13g2_decap_8
XFILLER_2_349 VPWR VGND sg13g2_decap_8
XFILLER_9_471 VPWR VGND sg13g2_decap_8
XFILLER_4_91 VPWR VGND sg13g2_decap_8
XFILLER_0_49 VPWR VGND sg13g2_decap_8
XFILLER_2_168 VPWR VGND sg13g2_decap_8
XFILLER_9_14 VPWR VGND sg13g2_decap_8
XFILLER_6_474 VPWR VGND sg13g2_decap_8
X_042_ FrameStrobe[10] net34 VPWR VGND sg13g2_buf_1
XFILLER_7_238 VPWR VGND sg13g2_decap_8
XFILLER_3_444 VPWR VGND sg13g2_decap_8
XFILLER_6_293 VPWR VGND sg13g2_decap_8
XFILLER_1_70 VPWR VGND sg13g2_decap_8
X_025_ FrameData[25] net18 VPWR VGND sg13g2_buf_1
XFILLER_0_469 VPWR VGND sg13g2_decap_8
Xoutput34 net34 FrameStrobe_O[10] VPWR VGND sg13g2_buf_1
Xoutput45 net45 FrameStrobe_O[2] VPWR VGND sg13g2_buf_1
Xoutput89 net89 NN4BEG[0] VPWR VGND sg13g2_buf_1
Xoutput78 net78 N4BEG[14] VPWR VGND sg13g2_buf_1
Xoutput67 net67 N2BEGb[2] VPWR VGND sg13g2_buf_1
Xoutput56 net56 N1BEG[3] VPWR VGND sg13g2_buf_1
XFILLER_0_266 VPWR VGND sg13g2_decap_8
Xoutput23 net23 FrameData_O[2] VPWR VGND sg13g2_buf_1
Xoutput12 net12 FrameData_O[1] VPWR VGND sg13g2_buf_1
XFILLER_8_322 VPWR VGND sg13g2_decap_8
X_008_ FrameData[8] net31 VPWR VGND sg13g2_buf_1
XFILLER_7_91 VPWR VGND sg13g2_decap_8
XFILLER_9_119 VPWR VGND sg13g2_decap_8
XFILLER_5_336 VPWR VGND sg13g2_decap_8
XFILLER_3_49 VPWR VGND sg13g2_decap_8
XFILLER_8_185 VPWR VGND sg13g2_fill_1
XFILLER_8_130 VPWR VGND sg13g2_decap_8
XFILLER_5_133 VPWR VGND sg13g2_decap_8
XFILLER_2_328 VPWR VGND sg13g2_decap_8
XFILLER_9_450 VPWR VGND sg13g2_decap_8
XFILLER_1_394 VPWR VGND sg13g2_decap_8
XFILLER_2_147 VPWR VGND sg13g2_decap_8
XFILLER_4_70 VPWR VGND sg13g2_decap_8
XFILLER_6_453 VPWR VGND sg13g2_decap_8
XFILLER_0_28 VPWR VGND sg13g2_decap_8
XFILLER_7_217 VPWR VGND sg13g2_decap_8
X_041_ FrameStrobe[9] net52 VPWR VGND sg13g2_buf_1
XFILLER_3_423 VPWR VGND sg13g2_decap_8
XFILLER_6_272 VPWR VGND sg13g2_decap_8
XFILLER_8_504 VPWR VGND sg13g2_decap_8
XFILLER_0_448 VPWR VGND sg13g2_decap_8
X_024_ FrameData[24] net17 VPWR VGND sg13g2_buf_1
XFILLER_6_49 VPWR VGND sg13g2_decap_8
XFILLER_3_297 VPWR VGND sg13g2_decap_8
Xoutput24 net24 FrameData_O[30] VPWR VGND sg13g2_buf_1
Xoutput35 net35 FrameStrobe_O[11] VPWR VGND sg13g2_buf_1
Xoutput46 net46 FrameStrobe_O[3] VPWR VGND sg13g2_buf_1
Xoutput57 net57 N2BEG[0] VPWR VGND sg13g2_buf_1
Xoutput13 net13 FrameData_O[20] VPWR VGND sg13g2_buf_1
XFILLER_5_518 VPWR VGND sg13g2_decap_4
Xoutput79 net79 N4BEG[15] VPWR VGND sg13g2_buf_1
Xoutput68 net68 N2BEGb[3] VPWR VGND sg13g2_buf_1
XFILLER_8_301 VPWR VGND sg13g2_decap_8
XFILLER_0_245 VPWR VGND sg13g2_decap_8
X_007_ FrameData[7] net30 VPWR VGND sg13g2_buf_1
XFILLER_7_70 VPWR VGND sg13g2_decap_8
XFILLER_3_28 VPWR VGND sg13g2_decap_8
XFILLER_4_392 VPWR VGND sg13g2_decap_8
XFILLER_2_307 VPWR VGND sg13g2_decap_8
XFILLER_5_189 VPWR VGND sg13g2_decap_8
XFILLER_5_112 VPWR VGND sg13g2_decap_8
XFILLER_1_373 VPWR VGND sg13g2_decap_8
XFILLER_9_49 VPWR VGND sg13g2_decap_8
XFILLER_6_432 VPWR VGND sg13g2_decap_8
XFILLER_2_126 VPWR VGND sg13g2_decap_8
X_040_ FrameStrobe[8] net51 VPWR VGND sg13g2_buf_1
XFILLER_3_402 VPWR VGND sg13g2_decap_8
XFILLER_3_479 VPWR VGND sg13g2_decap_8
XFILLER_0_427 VPWR VGND sg13g2_decap_8
X_023_ FrameData[23] net16 VPWR VGND sg13g2_buf_1
XFILLER_6_28 VPWR VGND sg13g2_decap_8
XFILLER_3_221 VPWR VGND sg13g2_fill_1
XFILLER_3_276 VPWR VGND sg13g2_decap_8
Xoutput25 net25 FrameData_O[31] VPWR VGND sg13g2_buf_1
Xoutput36 net36 FrameStrobe_O[12] VPWR VGND sg13g2_buf_1
Xoutput47 net47 FrameStrobe_O[4] VPWR VGND sg13g2_buf_1
Xoutput69 net69 N2BEGb[4] VPWR VGND sg13g2_buf_1
Xoutput58 net58 N2BEG[1] VPWR VGND sg13g2_buf_1
Xoutput14 net14 FrameData_O[21] VPWR VGND sg13g2_buf_1
XFILLER_0_224 VPWR VGND sg13g2_decap_8
X_006_ FrameData[6] net29 VPWR VGND sg13g2_buf_1
XFILLER_5_316 VPWR VGND sg13g2_fill_1
XFILLER_8_198 VPWR VGND sg13g2_fill_1
XFILLER_4_371 VPWR VGND sg13g2_decap_8
XFILLER_5_168 VPWR VGND sg13g2_decap_8
XFILLER_1_352 VPWR VGND sg13g2_decap_8
XFILLER_9_485 VPWR VGND sg13g2_decap_8
XFILLER_9_28 VPWR VGND sg13g2_decap_8
XFILLER_6_411 VPWR VGND sg13g2_decap_8
XFILLER_2_105 VPWR VGND sg13g2_decap_8
XFILLER_3_7 VPWR VGND sg13g2_decap_8
XFILLER_6_499 VPWR VGND sg13g2_fill_2
XFILLER_6_488 VPWR VGND sg13g2_decap_8
XFILLER_1_182 VPWR VGND sg13g2_decap_8
XFILLER_3_458 VPWR VGND sg13g2_decap_8
XFILLER_10_281 VPWR VGND sg13g2_decap_8
X_099_ SS4END[4] net91 VPWR VGND sg13g2_buf_1
XFILLER_6_252 VPWR VGND sg13g2_fill_2
XFILLER_1_84 VPWR VGND sg13g2_decap_8
XFILLER_0_406 VPWR VGND sg13g2_decap_8
X_022_ FrameData[22] net15 VPWR VGND sg13g2_buf_1
XFILLER_3_200 VPWR VGND sg13g2_fill_2
Xoutput15 net15 FrameData_O[22] VPWR VGND sg13g2_buf_1
Xoutput37 net37 FrameStrobe_O[13] VPWR VGND sg13g2_buf_1
Xoutput48 net48 FrameStrobe_O[5] VPWR VGND sg13g2_buf_1
Xoutput59 net59 N2BEG[2] VPWR VGND sg13g2_buf_1
XFILLER_0_203 VPWR VGND sg13g2_decap_8
Xoutput26 net26 FrameData_O[3] VPWR VGND sg13g2_buf_1
X_005_ FrameData[5] net28 VPWR VGND sg13g2_buf_1
XFILLER_5_328 VPWR VGND sg13g2_decap_4
XFILLER_8_144 VPWR VGND sg13g2_fill_2
XFILLER_8_111 VPWR VGND sg13g2_fill_1
XFILLER_4_350 VPWR VGND sg13g2_decap_8
XFILLER_5_147 VPWR VGND sg13g2_decap_8
XFILLER_1_331 VPWR VGND sg13g2_decap_8
XFILLER_9_464 VPWR VGND sg13g2_decap_8
XFILLER_4_84 VPWR VGND sg13g2_decap_8
XFILLER_6_467 VPWR VGND sg13g2_decap_8
XFILLER_1_161 VPWR VGND sg13g2_decap_8
XFILLER_10_260 VPWR VGND sg13g2_decap_8
X_098_ SS4END[5] net90 VPWR VGND sg13g2_buf_1
XFILLER_6_286 VPWR VGND sg13g2_decap_8
XFILLER_3_437 VPWR VGND sg13g2_decap_8
XFILLER_1_63 VPWR VGND sg13g2_decap_8
XFILLER_8_518 VPWR VGND sg13g2_fill_1
X_021_ FrameData[21] net14 VPWR VGND sg13g2_buf_1
XFILLER_3_234 VPWR VGND sg13g2_decap_4
Xoutput16 net16 FrameData_O[23] VPWR VGND sg13g2_buf_1
Xoutput38 net38 FrameStrobe_O[14] VPWR VGND sg13g2_buf_1
Xoutput49 net49 FrameStrobe_O[6] VPWR VGND sg13g2_buf_1
XFILLER_0_259 VPWR VGND sg13g2_decap_8
Xoutput27 net27 FrameData_O[4] VPWR VGND sg13g2_buf_1
XFILLER_8_348 VPWR VGND sg13g2_fill_1
XFILLER_8_315 VPWR VGND sg13g2_decap_8
X_004_ FrameData[4] net27 VPWR VGND sg13g2_buf_1
XFILLER_7_392 VPWR VGND sg13g2_fill_1
XFILLER_7_381 VPWR VGND sg13g2_fill_2
XFILLER_7_84 VPWR VGND sg13g2_decap_8
XFILLER_8_123 VPWR VGND sg13g2_decap_8
XFILLER_1_513 VPWR VGND sg13g2_decap_4
XFILLER_5_126 VPWR VGND sg13g2_decap_8
XFILLER_1_310 VPWR VGND sg13g2_decap_8
XFILLER_9_443 VPWR VGND sg13g2_decap_8
XFILLER_1_387 VPWR VGND sg13g2_decap_8
XFILLER_4_63 VPWR VGND sg13g2_decap_8
XFILLER_6_446 VPWR VGND sg13g2_decap_8
XFILLER_1_140 VPWR VGND sg13g2_decap_8
XFILLER_6_210 VPWR VGND sg13g2_decap_8
XFILLER_3_416 VPWR VGND sg13g2_decap_8
X_097_ SS4END[6] net104 VPWR VGND sg13g2_buf_1
XFILLER_6_265 VPWR VGND sg13g2_decap_8
XFILLER_1_42 VPWR VGND sg13g2_decap_8
XFILLER_2_482 VPWR VGND sg13g2_decap_8
X_020_ FrameData[20] net13 VPWR VGND sg13g2_buf_1
Xoutput17 net17 FrameData_O[24] VPWR VGND sg13g2_buf_1
Xoutput39 net39 FrameStrobe_O[15] VPWR VGND sg13g2_buf_1
XFILLER_0_238 VPWR VGND sg13g2_decap_8
Xoutput28 net28 FrameData_O[5] VPWR VGND sg13g2_buf_1
XFILLER_4_522 VPWR VGND sg13g2_fill_1
XFILLER_4_511 VPWR VGND sg13g2_decap_8
X_003_ FrameData[3] net26 VPWR VGND sg13g2_buf_1
XFILLER_7_63 VPWR VGND sg13g2_decap_8
XFILLER_8_102 VPWR VGND sg13g2_decap_8
XFILLER_8_146 VPWR VGND sg13g2_fill_1
XFILLER_4_385 VPWR VGND sg13g2_decap_8
XFILLER_5_105 VPWR VGND sg13g2_decap_8
XFILLER_9_499 VPWR VGND sg13g2_decap_8
XFILLER_9_422 VPWR VGND sg13g2_decap_8
XFILLER_1_366 VPWR VGND sg13g2_decap_8
XFILLER_4_42 VPWR VGND sg13g2_decap_8
XFILLER_4_182 VPWR VGND sg13g2_decap_8
XFILLER_2_119 VPWR VGND sg13g2_decap_8
XFILLER_10_432 VPWR VGND sg13g2_fill_1
XFILLER_10_421 VPWR VGND sg13g2_decap_8
XFILLER_8_0 VPWR VGND sg13g2_decap_8
XFILLER_6_425 VPWR VGND sg13g2_fill_2
XFILLER_1_196 VPWR VGND sg13g2_decap_8
XFILLER_9_252 VPWR VGND sg13g2_decap_8
XFILLER_1_7 VPWR VGND sg13g2_decap_8
XFILLER_10_295 VPWR VGND sg13g2_decap_8
X_096_ SS4END[7] net103 VPWR VGND sg13g2_buf_1
XFILLER_6_244 VPWR VGND sg13g2_decap_4
XFILLER_1_98 VPWR VGND sg13g2_decap_8
XFILLER_1_21 VPWR VGND sg13g2_decap_8
XFILLER_2_461 VPWR VGND sg13g2_decap_8
XFILLER_3_269 VPWR VGND sg13g2_decap_8
Xoutput18 net18 FrameData_O[25] VPWR VGND sg13g2_buf_1
X_079_ S4END[8] net86 VPWR VGND sg13g2_buf_1
XFILLER_0_217 VPWR VGND sg13g2_decap_8
Xoutput29 net29 FrameData_O[6] VPWR VGND sg13g2_buf_1
X_002_ FrameData[2] net23 VPWR VGND sg13g2_buf_1
XFILLER_7_383 VPWR VGND sg13g2_fill_1
XFILLER_7_361 VPWR VGND sg13g2_decap_8
XFILLER_7_42 VPWR VGND sg13g2_decap_8
XFILLER_5_309 VPWR VGND sg13g2_decap_8
XFILLER_4_364 VPWR VGND sg13g2_decap_8
XFILLER_9_478 VPWR VGND sg13g2_decap_8
XFILLER_9_401 VPWR VGND sg13g2_decap_8
XFILLER_1_345 VPWR VGND sg13g2_decap_8
XFILLER_4_21 VPWR VGND sg13g2_decap_8
XFILLER_4_98 VPWR VGND sg13g2_decap_8
XFILLER_4_161 VPWR VGND sg13g2_decap_8
XFILLER_10_400 VPWR VGND sg13g2_decap_8
XFILLER_6_404 VPWR VGND sg13g2_decap_8
XFILLER_1_175 VPWR VGND sg13g2_decap_8
XFILLER_10_274 VPWR VGND sg13g2_decap_8
X_095_ SS4END[8] net102 VPWR VGND sg13g2_buf_1
XFILLER_1_77 VPWR VGND sg13g2_decap_8
XFILLER_2_440 VPWR VGND sg13g2_decap_8
X_078_ S4END[9] net85 VPWR VGND sg13g2_buf_1
Xoutput19 net19 FrameData_O[26] VPWR VGND sg13g2_buf_1
X_001_ FrameData[1] net12 VPWR VGND sg13g2_buf_1
XFILLER_7_340 VPWR VGND sg13g2_decap_8
XFILLER_7_98 VPWR VGND sg13g2_fill_2
XFILLER_7_21 VPWR VGND sg13g2_decap_8
XFILLER_8_137 VPWR VGND sg13g2_decap_8
XFILLER_4_343 VPWR VGND sg13g2_decap_8
XFILLER_1_324 VPWR VGND sg13g2_decap_8
XFILLER_9_457 VPWR VGND sg13g2_decap_8
XFILLER_4_77 VPWR VGND sg13g2_decap_8
XFILLER_4_140 VPWR VGND sg13g2_decap_8
XFILLER_8_490 VPWR VGND sg13g2_decap_8
XFILLER_6_427 VPWR VGND sg13g2_fill_1
XFILLER_9_298 VPWR VGND sg13g2_decap_8
XFILLER_9_232 VPWR VGND sg13g2_fill_2
XFILLER_9_210 VPWR VGND sg13g2_fill_2
XFILLER_5_482 VPWR VGND sg13g2_decap_8
XFILLER_1_154 VPWR VGND sg13g2_decap_8
XFILLER_10_253 VPWR VGND sg13g2_decap_8
X_094_ SS4END[9] net101 VPWR VGND sg13g2_buf_1
XFILLER_6_279 VPWR VGND sg13g2_decap_8
XFILLER_6_224 VPWR VGND sg13g2_decap_4
XFILLER_2_496 VPWR VGND sg13g2_decap_8
XFILLER_1_56 VPWR VGND sg13g2_decap_8
X_077_ S4END[10] net84 VPWR VGND sg13g2_buf_1
XFILLER_2_293 VPWR VGND sg13g2_decap_8
XFILLER_8_308 VPWR VGND sg13g2_decap_8
XFILLER_7_77 VPWR VGND sg13g2_decap_8
X_000_ FrameData[0] net1 VPWR VGND sg13g2_buf_1
XFILLER_1_506 VPWR VGND sg13g2_decap_8
XFILLER_1_517 VPWR VGND sg13g2_fill_2
XFILLER_8_116 VPWR VGND sg13g2_decap_8
XFILLER_4_399 VPWR VGND sg13g2_decap_8
XFILLER_4_322 VPWR VGND sg13g2_fill_2
XFILLER_7_182 VPWR VGND sg13g2_decap_8
XFILLER_5_119 VPWR VGND sg13g2_decap_8
XFILLER_1_303 VPWR VGND sg13g2_decap_8
XFILLER_9_436 VPWR VGND sg13g2_decap_8
XFILLER_4_56 VPWR VGND sg13g2_decap_8
XFILLER_4_196 VPWR VGND sg13g2_decap_8
XFILLER_6_439 VPWR VGND sg13g2_decap_8
XFILLER_1_133 VPWR VGND sg13g2_decap_8
XFILLER_3_409 VPWR VGND sg13g2_decap_8
XFILLER_10_232 VPWR VGND sg13g2_decap_8
X_093_ SS4END[10] net100 VPWR VGND sg13g2_buf_1
XFILLER_6_258 VPWR VGND sg13g2_decap_8
XFILLER_6_203 VPWR VGND sg13g2_decap_8
XFILLER_6_0 VPWR VGND sg13g2_decap_8
XFILLER_1_35 VPWR VGND sg13g2_decap_8
XFILLER_2_475 VPWR VGND sg13g2_decap_8
XFILLER_3_206 VPWR VGND sg13g2_decap_8
X_076_ S4END[11] net83 VPWR VGND sg13g2_buf_1
XFILLER_2_261 VPWR VGND sg13g2_decap_8
XFILLER_4_504 VPWR VGND sg13g2_decap_8
X_059_ S2MID[4] net60 VPWR VGND sg13g2_buf_1
XFILLER_7_397 VPWR VGND sg13g2_decap_8
XFILLER_7_375 VPWR VGND sg13g2_fill_2
XFILLER_7_56 VPWR VGND sg13g2_decap_8
XFILLER_4_301 VPWR VGND sg13g2_decap_8
XFILLER_4_378 VPWR VGND sg13g2_decap_8
XFILLER_1_359 VPWR VGND sg13g2_decap_8
XFILLER_9_415 VPWR VGND sg13g2_decap_8
XFILLER_0_392 VPWR VGND sg13g2_decap_8
XFILLER_4_35 VPWR VGND sg13g2_decap_8
XFILLER_4_175 VPWR VGND sg13g2_decap_8
XFILLER_10_414 VPWR VGND sg13g2_decap_8
XFILLER_6_418 VPWR VGND sg13g2_decap_8
XFILLER_1_189 VPWR VGND sg13g2_decap_8
XFILLER_1_112 VPWR VGND sg13g2_decap_8
XFILLER_9_245 VPWR VGND sg13g2_decap_8
XFILLER_9_212 VPWR VGND sg13g2_fill_1
XFILLER_5_462 VPWR VGND sg13g2_decap_8
XFILLER_10_288 VPWR VGND sg13g2_decap_8
X_092_ SS4END[11] net99 VPWR VGND sg13g2_buf_1
XFILLER_6_237 VPWR VGND sg13g2_decap_8
XFILLER_1_14 VPWR VGND sg13g2_decap_8
XFILLER_2_454 VPWR VGND sg13g2_decap_8
XFILLER_5_270 VPWR VGND sg13g2_decap_4
X_075_ S4END[12] net82 VPWR VGND sg13g2_buf_1
XFILLER_7_502 VPWR VGND sg13g2_decap_8
XFILLER_7_354 VPWR VGND sg13g2_decap_8
X_058_ S2MID[5] net59 VPWR VGND sg13g2_buf_1
XFILLER_7_35 VPWR VGND sg13g2_decap_8
XFILLER_4_324 VPWR VGND sg13g2_fill_1
XFILLER_4_357 VPWR VGND sg13g2_decap_8
XFILLER_7_162 VPWR VGND sg13g2_fill_2
XFILLER_1_338 VPWR VGND sg13g2_decap_8
XFILLER_4_14 VPWR VGND sg13g2_decap_8
XFILLER_4_154 VPWR VGND sg13g2_decap_8
XFILLER_0_371 VPWR VGND sg13g2_decap_8
XFILLER_1_168 VPWR VGND sg13g2_decap_8
XFILLER_5_496 VPWR VGND sg13g2_decap_4
XFILLER_5_441 VPWR VGND sg13g2_decap_8
XFILLER_10_267 VPWR VGND sg13g2_decap_8
X_091_ SS4END[12] net98 VPWR VGND sg13g2_buf_1
XFILLER_2_433 VPWR VGND sg13g2_decap_8
XFILLER_5_293 VPWR VGND sg13g2_decap_4
X_074_ S4END[13] net81 VPWR VGND sg13g2_buf_1
XFILLER_2_91 VPWR VGND sg13g2_decap_8
XFILLER_7_388 VPWR VGND sg13g2_decap_4
XFILLER_7_333 VPWR VGND sg13g2_decap_8
X_057_ S2MID[6] net58 VPWR VGND sg13g2_buf_1
XFILLER_7_14 VPWR VGND sg13g2_decap_8
XFILLER_4_336 VPWR VGND sg13g2_decap_8
XFILLER_7_196 VPWR VGND sg13g2_decap_8
XFILLER_1_317 VPWR VGND sg13g2_decap_8
XFILLER_8_483 VPWR VGND sg13g2_decap_8
XFILLER_0_350 VPWR VGND sg13g2_decap_8
XFILLER_4_133 VPWR VGND sg13g2_decap_8
XFILLER_1_147 VPWR VGND sg13g2_decap_8
XFILLER_9_203 VPWR VGND sg13g2_decap_8
XFILLER_5_475 VPWR VGND sg13g2_decap_8
XFILLER_5_420 VPWR VGND sg13g2_decap_8
XFILLER_5_91 VPWR VGND sg13g2_decap_8
XFILLER_10_246 VPWR VGND sg13g2_decap_8
X_090_ SS4END[13] net97 VPWR VGND sg13g2_buf_1
XFILLER_6_228 VPWR VGND sg13g2_fill_1
XFILLER_6_217 VPWR VGND sg13g2_decap_8
XFILLER_1_49 VPWR VGND sg13g2_decap_8
XFILLER_2_412 VPWR VGND sg13g2_decap_8
XFILLER_2_489 VPWR VGND sg13g2_decap_8
XFILLER_10_14 VPWR VGND sg13g2_fill_2
X_073_ S4END[14] net80 VPWR VGND sg13g2_buf_1
XFILLER_2_275 VPWR VGND sg13g2_decap_8
XFILLER_2_286 VPWR VGND sg13g2_decap_8
XFILLER_4_0 VPWR VGND sg13g2_decap_8
XFILLER_4_518 VPWR VGND sg13g2_decap_4
XFILLER_2_70 VPWR VGND sg13g2_decap_8
X_056_ S2MID[7] net57 VPWR VGND sg13g2_buf_1
XFILLER_7_312 VPWR VGND sg13g2_decap_8
XFILLER_8_109 VPWR VGND sg13g2_fill_2
XFILLER_4_315 VPWR VGND sg13g2_fill_2
XFILLER_7_175 VPWR VGND sg13g2_decap_8
XFILLER_3_381 VPWR VGND sg13g2_decap_8
X_039_ FrameStrobe[7] net50 VPWR VGND sg13g2_buf_1
XFILLER_8_91 VPWR VGND sg13g2_fill_2
XFILLER_9_429 VPWR VGND sg13g2_decap_8
XFILLER_4_49 VPWR VGND sg13g2_decap_8
XFILLER_4_112 VPWR VGND sg13g2_decap_8
XFILLER_4_189 VPWR VGND sg13g2_decap_8
XFILLER_10_428 VPWR VGND sg13g2_decap_4
XFILLER_8_462 VPWR VGND sg13g2_decap_8
XFILLER_9_259 VPWR VGND sg13g2_decap_8
XFILLER_9_226 VPWR VGND sg13g2_fill_2
XFILLER_8_7 VPWR VGND sg13g2_decap_8
XFILLER_1_126 VPWR VGND sg13g2_decap_8
XFILLER_5_70 VPWR VGND sg13g2_decap_8
XFILLER_10_225 VPWR VGND sg13g2_decap_8
XFILLER_1_28 VPWR VGND sg13g2_decap_8
XFILLER_2_468 VPWR VGND sg13g2_decap_8
X_072_ S4END[15] net73 VPWR VGND sg13g2_buf_1
XFILLER_7_516 VPWR VGND sg13g2_decap_8
XFILLER_2_210 VPWR VGND sg13g2_decap_4
XFILLER_2_232 VPWR VGND sg13g2_decap_8
XFILLER_2_254 VPWR VGND sg13g2_decap_8
X_055_ S1END[0] net56 VPWR VGND sg13g2_buf_1
XFILLER_7_368 VPWR VGND sg13g2_decap_8
XFILLER_7_49 VPWR VGND sg13g2_decap_8
XFILLER_7_121 VPWR VGND sg13g2_decap_4
XFILLER_3_360 VPWR VGND sg13g2_decap_8
X_038_ FrameStrobe[6] net49 VPWR VGND sg13g2_buf_1
XFILLER_9_408 VPWR VGND sg13g2_decap_8
XFILLER_0_385 VPWR VGND sg13g2_decap_8
XFILLER_4_28 VPWR VGND sg13g2_decap_8
XFILLER_4_168 VPWR VGND sg13g2_decap_8
XFILLER_10_407 VPWR VGND sg13g2_decap_8
XFILLER_8_441 VPWR VGND sg13g2_decap_8
XFILLER_9_238 VPWR VGND sg13g2_decap_8
XFILLER_1_105 VPWR VGND sg13g2_decap_8
XFILLER_8_282 VPWR VGND sg13g2_fill_1
XFILLER_8_271 VPWR VGND sg13g2_decap_8
XFILLER_5_455 VPWR VGND sg13g2_decap_8
XFILLER_0_182 VPWR VGND sg13g2_decap_8
XFILLER_2_447 VPWR VGND sg13g2_decap_8
XFILLER_5_274 VPWR VGND sg13g2_fill_1
XFILLER_5_252 VPWR VGND sg13g2_decap_8
XFILLER_10_16 VPWR VGND sg13g2_fill_1
X_071_ S2END[0] net72 VPWR VGND sg13g2_buf_1
XFILLER_2_244 VPWR VGND sg13g2_fill_2
X_054_ S1END[1] net55 VPWR VGND sg13g2_buf_1
XFILLER_7_347 VPWR VGND sg13g2_decap_8
XFILLER_7_28 VPWR VGND sg13g2_decap_8
XFILLER_4_317 VPWR VGND sg13g2_fill_1
XFILLER_7_155 VPWR VGND sg13g2_decap_8
XFILLER_7_100 VPWR VGND sg13g2_fill_1
X_037_ FrameStrobe[5] net48 VPWR VGND sg13g2_buf_1
XFILLER_8_93 VPWR VGND sg13g2_fill_1
XFILLER_0_364 VPWR VGND sg13g2_decap_8
XFILLER_4_147 VPWR VGND sg13g2_decap_8
XFILLER_8_497 VPWR VGND sg13g2_decap_8
XFILLER_8_420 VPWR VGND sg13g2_decap_8
XFILLER_9_217 VPWR VGND sg13g2_fill_1
XFILLER_5_489 VPWR VGND sg13g2_decap_8
XFILLER_5_434 VPWR VGND sg13g2_decap_8
XFILLER_0_161 VPWR VGND sg13g2_decap_8
XFILLER_8_294 VPWR VGND sg13g2_decap_8
XFILLER_8_250 VPWR VGND sg13g2_decap_8
XFILLER_5_231 VPWR VGND sg13g2_decap_8
XFILLER_2_426 VPWR VGND sg13g2_decap_8
XFILLER_5_297 VPWR VGND sg13g2_fill_1
XFILLER_5_286 VPWR VGND sg13g2_decap_8
XFILLER_1_492 VPWR VGND sg13g2_decap_8
X_070_ S2END[1] net71 VPWR VGND sg13g2_buf_1
XFILLER_2_84 VPWR VGND sg13g2_decap_8
X_053_ S1END[2] net54 VPWR VGND sg13g2_buf_1
XFILLER_7_326 VPWR VGND sg13g2_decap_8
XFILLER_2_0 VPWR VGND sg13g2_decap_8
XFILLER_3_521 VPWR VGND sg13g2_fill_2
XFILLER_4_329 VPWR VGND sg13g2_decap_8
XFILLER_8_50 VPWR VGND sg13g2_fill_1
XFILLER_7_189 VPWR VGND sg13g2_decap_8
X_036_ FrameStrobe[4] net47 VPWR VGND sg13g2_buf_1
XFILLER_3_395 VPWR VGND sg13g2_decap_8
XFILLER_4_126 VPWR VGND sg13g2_decap_8
XFILLER_8_476 VPWR VGND sg13g2_decap_8
X_019_ FrameData[19] net11 VPWR VGND sg13g2_buf_1
XFILLER_0_343 VPWR VGND sg13g2_decap_8
XFILLER_5_413 VPWR VGND sg13g2_decap_8
XFILLER_0_140 VPWR VGND sg13g2_decap_8
XFILLER_5_84 VPWR VGND sg13g2_decap_8
XFILLER_4_490 VPWR VGND sg13g2_decap_8
XFILLER_10_239 VPWR VGND sg13g2_decap_8
XFILLER_6_7 VPWR VGND sg13g2_decap_8
XFILLER_2_405 VPWR VGND sg13g2_decap_8
XFILLER_5_210 VPWR VGND sg13g2_decap_8
XFILLER_1_471 VPWR VGND sg13g2_decap_8
XFILLER_2_268 VPWR VGND sg13g2_decap_8
XFILLER_2_63 VPWR VGND sg13g2_decap_8
X_052_ S1END[3] net53 VPWR VGND sg13g2_buf_1
XFILLER_7_305 VPWR VGND sg13g2_decap_8
XFILLER_3_500 VPWR VGND sg13g2_decap_8
XFILLER_6_382 VPWR VGND sg13g2_decap_8
XFILLER_4_308 VPWR VGND sg13g2_decap_8
XFILLER_7_168 VPWR VGND sg13g2_decap_8
XFILLER_7_135 VPWR VGND sg13g2_decap_4
X_035_ FrameStrobe[3] net46 VPWR VGND sg13g2_buf_1
X_104_ UserCLK net105 VPWR VGND sg13g2_buf_1
XFILLER_3_374 VPWR VGND sg13g2_decap_8
XFILLER_8_84 VPWR VGND sg13g2_decap_8
XFILLER_8_62 VPWR VGND sg13g2_decap_8
XFILLER_4_105 VPWR VGND sg13g2_decap_8
XFILLER_8_455 VPWR VGND sg13g2_decap_8
XFILLER_0_322 VPWR VGND sg13g2_decap_8
XFILLER_0_399 VPWR VGND sg13g2_decap_8
X_018_ FrameData[18] net10 VPWR VGND sg13g2_buf_1
XFILLER_1_119 VPWR VGND sg13g2_decap_8
XFILLER_3_182 VPWR VGND sg13g2_decap_8
XFILLER_5_469 VPWR VGND sg13g2_fill_2
XFILLER_0_196 VPWR VGND sg13g2_decap_8
XFILLER_10_0 VPWR VGND sg13g2_decap_8
XFILLER_5_63 VPWR VGND sg13g2_decap_8
XFILLER_1_450 VPWR VGND sg13g2_decap_8
XFILLER_7_509 VPWR VGND sg13g2_decap_8
XFILLER_2_203 VPWR VGND sg13g2_decap_8
XFILLER_2_225 VPWR VGND sg13g2_fill_2
XFILLER_9_380 VPWR VGND sg13g2_decap_8
XFILLER_2_42 VPWR VGND sg13g2_decap_8
X_051_ FrameStrobe[19] net43 VPWR VGND sg13g2_buf_1
XFILLER_6_361 VPWR VGND sg13g2_decap_8
XFILLER_0_504 VPWR VGND sg13g2_decap_8
X_103_ SS4END[0] net95 VPWR VGND sg13g2_buf_1
XFILLER_7_125 VPWR VGND sg13g2_fill_2
XFILLER_7_114 VPWR VGND sg13g2_fill_2
X_034_ FrameStrobe[2] net45 VPWR VGND sg13g2_buf_1
XFILLER_3_353 VPWR VGND sg13g2_decap_8
XFILLER_8_41 VPWR VGND sg13g2_fill_1
XFILLER_8_434 VPWR VGND sg13g2_decap_8
XFILLER_0_301 VPWR VGND sg13g2_decap_8
XFILLER_0_378 VPWR VGND sg13g2_decap_8
X_017_ FrameData[17] net9 VPWR VGND sg13g2_buf_1
XFILLER_3_161 VPWR VGND sg13g2_decap_8
XFILLER_5_448 VPWR VGND sg13g2_decap_8
XFILLER_8_264 VPWR VGND sg13g2_decap_8
XFILLER_5_42 VPWR VGND sg13g2_decap_8
XFILLER_0_175 VPWR VGND sg13g2_decap_8
XFILLER_5_245 VPWR VGND sg13g2_decap_8
XFILLER_2_21 VPWR VGND sg13g2_decap_8
XFILLER_2_98 VPWR VGND sg13g2_decap_8
Xoutput100 net100 NN4BEG[5] VPWR VGND sg13g2_buf_1
X_050_ FrameStrobe[18] net42 VPWR VGND sg13g2_buf_1
X_102_ SS4END[1] net94 VPWR VGND sg13g2_buf_1
XFILLER_7_148 VPWR VGND sg13g2_decap_8
X_033_ FrameStrobe[1] net44 VPWR VGND sg13g2_buf_1
XFILLER_0_0 VPWR VGND sg13g2_decap_8
XFILLER_3_332 VPWR VGND sg13g2_decap_8
XFILLER_0_357 VPWR VGND sg13g2_decap_8
XFILLER_8_413 VPWR VGND sg13g2_decap_8
X_016_ FrameData[16] net8 VPWR VGND sg13g2_buf_1
XFILLER_3_140 VPWR VGND sg13g2_decap_8
XFILLER_8_287 VPWR VGND sg13g2_decap_8
XFILLER_8_243 VPWR VGND sg13g2_decap_8
XFILLER_5_427 VPWR VGND sg13g2_decap_8
XFILLER_5_21 VPWR VGND sg13g2_decap_8
XFILLER_0_154 VPWR VGND sg13g2_decap_8
XFILLER_5_98 VPWR VGND sg13g2_decap_8
XFILLER_2_419 VPWR VGND sg13g2_decap_8
XFILLER_5_279 VPWR VGND sg13g2_decap_8
XFILLER_5_224 VPWR VGND sg13g2_decap_8
XFILLER_1_485 VPWR VGND sg13g2_decap_8
XFILLER_2_227 VPWR VGND sg13g2_fill_1
XFILLER_4_7 VPWR VGND sg13g2_decap_8
XFILLER_1_282 VPWR VGND sg13g2_decap_8
XFILLER_2_77 VPWR VGND sg13g2_decap_8
Xoutput101 net101 NN4BEG[6] VPWR VGND sg13g2_buf_1
XFILLER_7_319 VPWR VGND sg13g2_decap_8
XFILLER_3_514 VPWR VGND sg13g2_decap_8
XFILLER_6_396 VPWR VGND sg13g2_decap_4
X_101_ SS4END[2] net93 VPWR VGND sg13g2_buf_1
XFILLER_7_116 VPWR VGND sg13g2_fill_1
X_032_ FrameStrobe[0] net33 VPWR VGND sg13g2_buf_1
XFILLER_3_311 VPWR VGND sg13g2_decap_8
XFILLER_3_388 VPWR VGND sg13g2_decap_8
XFILLER_8_32 VPWR VGND sg13g2_fill_1
XFILLER_6_182 VPWR VGND sg13g2_decap_8
XFILLER_0_336 VPWR VGND sg13g2_decap_8
XFILLER_4_119 VPWR VGND sg13g2_decap_8
XFILLER_8_469 VPWR VGND sg13g2_decap_8
X_015_ FrameData[15] net7 VPWR VGND sg13g2_buf_1
XFILLER_3_196 VPWR VGND sg13g2_decap_4
XFILLER_5_406 VPWR VGND sg13g2_decap_8
XFILLER_0_133 VPWR VGND sg13g2_decap_8
XFILLER_8_222 VPWR VGND sg13g2_decap_8
XFILLER_5_77 VPWR VGND sg13g2_decap_8
XFILLER_4_483 VPWR VGND sg13g2_decap_8
XFILLER_5_203 VPWR VGND sg13g2_decap_8
XFILLER_1_464 VPWR VGND sg13g2_decap_8
XFILLER_4_280 VPWR VGND sg13g2_decap_8
XFILLER_2_239 VPWR VGND sg13g2_fill_1
XFILLER_6_512 VPWR VGND sg13g2_decap_8
XFILLER_1_261 VPWR VGND sg13g2_decap_8
XFILLER_2_56 VPWR VGND sg13g2_decap_8
XFILLER_9_394 VPWR VGND sg13g2_decap_8
Xoutput102 net102 NN4BEG[7] VPWR VGND sg13g2_buf_1
XFILLER_10_393 VPWR VGND sg13g2_decap_8
XFILLER_6_375 VPWR VGND sg13g2_decap_8
XFILLER_6_342 VPWR VGND sg13g2_decap_8
X_031_ FrameData[31] net25 VPWR VGND sg13g2_buf_1
X_100_ SS4END[3] net92 VPWR VGND sg13g2_buf_1
XFILLER_7_139 VPWR VGND sg13g2_fill_1
XFILLER_8_77 VPWR VGND sg13g2_decap_8
XFILLER_8_55 VPWR VGND sg13g2_decap_8
XFILLER_6_161 VPWR VGND sg13g2_decap_8
XFILLER_3_367 VPWR VGND sg13g2_decap_8
XFILLER_0_315 VPWR VGND sg13g2_decap_8
XFILLER_8_448 VPWR VGND sg13g2_decap_8
X_014_ FrameData[14] net6 VPWR VGND sg13g2_buf_1
XFILLER_3_175 VPWR VGND sg13g2_decap_8
XFILLER_7_481 VPWR VGND sg13g2_decap_8
XFILLER_0_189 VPWR VGND sg13g2_decap_8
XFILLER_0_112 VPWR VGND sg13g2_decap_8
XFILLER_8_278 VPWR VGND sg13g2_decap_4
XFILLER_5_56 VPWR VGND sg13g2_decap_8
XFILLER_4_462 VPWR VGND sg13g2_decap_8
XFILLER_5_259 VPWR VGND sg13g2_decap_8
XFILLER_1_443 VPWR VGND sg13g2_decap_8
XFILLER_2_218 VPWR VGND sg13g2_decap_8
XFILLER_9_373 VPWR VGND sg13g2_decap_8
Xoutput103 net103 NN4BEG[8] VPWR VGND sg13g2_buf_1
XFILLER_2_35 VPWR VGND sg13g2_decap_8
XFILLER_10_372 VPWR VGND sg13g2_decap_8
XFILLER_6_354 VPWR VGND sg13g2_decap_8
XFILLER_6_321 VPWR VGND sg13g2_decap_8
X_030_ FrameData[30] net24 VPWR VGND sg13g2_buf_1
XFILLER_3_346 VPWR VGND sg13g2_decap_8
XFILLER_6_140 VPWR VGND sg13g2_decap_8
XFILLER_8_427 VPWR VGND sg13g2_decap_8
X_013_ FrameData[13] net5 VPWR VGND sg13g2_buf_1
XFILLER_3_154 VPWR VGND sg13g2_decap_8
XFILLER_7_460 VPWR VGND sg13g2_decap_8
XFILLER_0_168 VPWR VGND sg13g2_decap_8
XFILLER_8_257 VPWR VGND sg13g2_decap_8
XFILLER_5_35 VPWR VGND sg13g2_decap_8
XFILLER_4_441 VPWR VGND sg13g2_decap_8
XFILLER_5_238 VPWR VGND sg13g2_decap_8
XFILLER_1_422 VPWR VGND sg13g2_decap_8
XFILLER_1_499 VPWR VGND sg13g2_decap_8
XFILLER_9_352 VPWR VGND sg13g2_decap_8
Xoutput104 net104 NN4BEG[9] VPWR VGND sg13g2_buf_1
XFILLER_9_0 VPWR VGND sg13g2_decap_8
XFILLER_1_296 VPWR VGND sg13g2_decap_8
XFILLER_2_14 VPWR VGND sg13g2_decap_8
XFILLER_2_7 VPWR VGND sg13g2_decap_8
XFILLER_10_351 VPWR VGND sg13g2_decap_8
XFILLER_6_300 VPWR VGND sg13g2_decap_8
XFILLER_9_182 VPWR VGND sg13g2_decap_8
XFILLER_3_325 VPWR VGND sg13g2_decap_8
X_089_ SS4END[14] net96 VPWR VGND sg13g2_buf_1
XFILLER_8_46 VPWR VGND sg13g2_decap_4
XFILLER_6_196 VPWR VGND sg13g2_decap_8
XFILLER_2_391 VPWR VGND sg13g2_decap_8
XFILLER_8_406 VPWR VGND sg13g2_decap_8
X_012_ FrameData[12] net4 VPWR VGND sg13g2_buf_1
XFILLER_3_133 VPWR VGND sg13g2_decap_8
XFILLER_0_91 VPWR VGND sg13g2_decap_8
XFILLER_8_236 VPWR VGND sg13g2_decap_8
XFILLER_8_203 VPWR VGND sg13g2_fill_1
XFILLER_5_14 VPWR VGND sg13g2_decap_8
XFILLER_4_497 VPWR VGND sg13g2_decap_8
XFILLER_4_420 VPWR VGND sg13g2_decap_8
XFILLER_0_147 VPWR VGND sg13g2_decap_8
XFILLER_7_291 VPWR VGND sg13g2_decap_8
XFILLER_5_217 VPWR VGND sg13g2_decap_8
XFILLER_1_401 VPWR VGND sg13g2_decap_8
XFILLER_1_478 VPWR VGND sg13g2_decap_8
XFILLER_4_294 VPWR VGND sg13g2_decap_8
XFILLER_9_331 VPWR VGND sg13g2_decap_8
XFILLER_1_275 VPWR VGND sg13g2_decap_8
XFILLER_1_231 VPWR VGND sg13g2_decap_8
Xoutput105 net105 UserCLKo VPWR VGND sg13g2_buf_1
XFILLER_3_507 VPWR VGND sg13g2_decap_8
XFILLER_10_330 VPWR VGND sg13g2_decap_8
XFILLER_6_389 VPWR VGND sg13g2_decap_8
XFILLER_9_161 VPWR VGND sg13g2_decap_8
XFILLER_7_109 VPWR VGND sg13g2_fill_1
XFILLER_3_91 VPWR VGND sg13g2_decap_8
XFILLER_3_304 VPWR VGND sg13g2_decap_8
X_088_ SS4END[15] net89 VPWR VGND sg13g2_buf_1
XFILLER_8_25 VPWR VGND sg13g2_decap_8
XFILLER_8_14 VPWR VGND sg13g2_decap_8
XFILLER_6_175 VPWR VGND sg13g2_decap_8
XFILLER_2_370 VPWR VGND sg13g2_decap_8
XFILLER_0_329 VPWR VGND sg13g2_decap_8
XFILLER_3_112 VPWR VGND sg13g2_decap_8
XFILLER_3_189 VPWR VGND sg13g2_decap_8
X_011_ FrameData[11] net3 VPWR VGND sg13g2_buf_1
XFILLER_7_495 VPWR VGND sg13g2_decap_8
XFILLER_0_70 VPWR VGND sg13g2_decap_8
XFILLER_8_215 VPWR VGND sg13g2_decap_8
XFILLER_0_126 VPWR VGND sg13g2_decap_8
XFILLER_10_7 VPWR VGND sg13g2_decap_8
XFILLER_4_476 VPWR VGND sg13g2_decap_8
XFILLER_1_457 VPWR VGND sg13g2_decap_8
XFILLER_0_490 VPWR VGND sg13g2_decap_8
XFILLER_4_273 VPWR VGND sg13g2_decap_8
XFILLER_6_91 VPWR VGND sg13g2_decap_8
XFILLER_6_505 VPWR VGND sg13g2_decap_8
XFILLER_1_254 VPWR VGND sg13g2_decap_8
XFILLER_1_210 VPWR VGND sg13g2_decap_8
XFILLER_2_49 VPWR VGND sg13g2_decap_8
XFILLER_9_387 VPWR VGND sg13g2_decap_8
XFILLER_10_386 VPWR VGND sg13g2_decap_8
XFILLER_6_335 VPWR VGND sg13g2_decap_8
XFILLER_9_140 VPWR VGND sg13g2_decap_8
XFILLER_6_368 VPWR VGND sg13g2_decap_8
XFILLER_3_70 VPWR VGND sg13g2_decap_8
X_087_ S4END[0] net79 VPWR VGND sg13g2_buf_1
XFILLER_8_37 VPWR VGND sg13g2_decap_4
XFILLER_6_154 VPWR VGND sg13g2_decap_8
XFILLER_0_308 VPWR VGND sg13g2_decap_8
XFILLER_3_168 VPWR VGND sg13g2_decap_8
X_010_ FrameData[10] net2 VPWR VGND sg13g2_buf_1
XFILLER_7_474 VPWR VGND sg13g2_decap_8
XFILLER_9_91 VPWR VGND sg13g2_decap_8
XFILLER_0_105 VPWR VGND sg13g2_decap_8
XFILLER_5_49 VPWR VGND sg13g2_decap_8
XFILLER_4_455 VPWR VGND sg13g2_decap_8
XFILLER_1_436 VPWR VGND sg13g2_decap_8
XFILLER_4_252 VPWR VGND sg13g2_decap_8
XFILLER_6_70 VPWR VGND sg13g2_decap_8
XFILLER_2_28 VPWR VGND sg13g2_decap_8
XFILLER_9_366 VPWR VGND sg13g2_decap_8
XFILLER_10_365 VPWR VGND sg13g2_decap_8
XFILLER_7_0 VPWR VGND sg13g2_decap_8
XFILLER_6_314 VPWR VGND sg13g2_decap_8
XFILLER_9_196 VPWR VGND sg13g2_decap_8
X_086_ S4END[1] net78 VPWR VGND sg13g2_buf_1
XFILLER_6_133 VPWR VGND sg13g2_decap_8
XFILLER_0_7 VPWR VGND sg13g2_decap_8
XFILLER_3_339 VPWR VGND sg13g2_decap_8
XFILLER_3_147 VPWR VGND sg13g2_decap_8
XFILLER_7_453 VPWR VGND sg13g2_decap_8
X_069_ S2END[2] net70 VPWR VGND sg13g2_buf_1
XFILLER_9_70 VPWR VGND sg13g2_decap_8
XFILLER_5_28 VPWR VGND sg13g2_decap_8
XFILLER_4_434 VPWR VGND sg13g2_decap_8
XFILLER_1_415 VPWR VGND sg13g2_decap_8
XFILLER_4_231 VPWR VGND sg13g2_decap_8
XFILLER_1_245 VPWR VGND sg13g2_decap_4
XFILLER_9_345 VPWR VGND sg13g2_decap_8
XFILLER_9_312 VPWR VGND sg13g2_fill_1
Xoutput90 net90 NN4BEG[10] VPWR VGND sg13g2_buf_1
XFILLER_1_289 VPWR VGND sg13g2_decap_8
XFILLER_10_344 VPWR VGND sg13g2_decap_8
XFILLER_2_510 VPWR VGND sg13g2_decap_8
XFILLER_2_521 VPWR VGND sg13g2_fill_2
XFILLER_9_175 VPWR VGND sg13g2_decap_8
XFILLER_5_392 VPWR VGND sg13g2_decap_8
XFILLER_3_318 VPWR VGND sg13g2_decap_8
X_085_ S4END[2] net77 VPWR VGND sg13g2_buf_1
XFILLER_6_189 VPWR VGND sg13g2_decap_8
XFILLER_6_112 VPWR VGND sg13g2_decap_8
XFILLER_2_384 VPWR VGND sg13g2_decap_8
XFILLER_3_126 VPWR VGND sg13g2_decap_8
XFILLER_7_432 VPWR VGND sg13g2_decap_8
X_068_ S2END[3] net69 VPWR VGND sg13g2_buf_1
XFILLER_0_84 VPWR VGND sg13g2_decap_8
XFILLER_8_229 VPWR VGND sg13g2_decap_8
XFILLER_4_413 VPWR VGND sg13g2_decap_8
XFILLER_7_284 VPWR VGND sg13g2_fill_2
XFILLER_4_210 VPWR VGND sg13g2_decap_8
XFILLER_4_287 VPWR VGND sg13g2_decap_8
XFILLER_6_519 VPWR VGND sg13g2_decap_4
XFILLER_9_324 VPWR VGND sg13g2_decap_8
XFILLER_1_268 VPWR VGND sg13g2_decap_8
XFILLER_1_224 VPWR VGND sg13g2_decap_8
Xoutput1 net1 FrameData_O[0] VPWR VGND sg13g2_buf_1
Xoutput91 net91 NN4BEG[11] VPWR VGND sg13g2_buf_1
Xoutput80 net80 N4BEG[1] VPWR VGND sg13g2_buf_1
XFILLER_10_323 VPWR VGND sg13g2_decap_8
XFILLER_6_349 VPWR VGND sg13g2_fill_1
XFILLER_9_154 VPWR VGND sg13g2_decap_8
XFILLER_5_371 VPWR VGND sg13g2_decap_8
XFILLER_3_84 VPWR VGND sg13g2_decap_8
X_084_ S4END[3] net76 VPWR VGND sg13g2_buf_1
XFILLER_6_168 VPWR VGND sg13g2_decap_8
XFILLER_2_363 VPWR VGND sg13g2_decap_8
XFILLER_7_488 VPWR VGND sg13g2_decap_8
XFILLER_7_411 VPWR VGND sg13g2_decap_8
XFILLER_3_105 VPWR VGND sg13g2_decap_8
X_067_ S2END[4] net68 VPWR VGND sg13g2_buf_1
XFILLER_0_63 VPWR VGND sg13g2_decap_8
XFILLER_2_182 VPWR VGND sg13g2_decap_8
XFILLER_8_208 VPWR VGND sg13g2_decap_8
XFILLER_4_469 VPWR VGND sg13g2_decap_8
XFILLER_0_119 VPWR VGND sg13g2_decap_8
XFILLER_7_252 VPWR VGND sg13g2_decap_8
XFILLER_9_506 VPWR VGND sg13g2_fill_1
XFILLER_0_483 VPWR VGND sg13g2_decap_8
XFILLER_4_266 VPWR VGND sg13g2_decap_8
XFILLER_6_84 VPWR VGND sg13g2_decap_8
XFILLER_1_203 VPWR VGND sg13g2_decap_8
Xoutput92 net92 NN4BEG[12] VPWR VGND sg13g2_buf_1
Xoutput81 net81 N4BEG[2] VPWR VGND sg13g2_buf_1
Xoutput70 net70 N2BEGb[5] VPWR VGND sg13g2_buf_1
XFILLER_0_280 VPWR VGND sg13g2_decap_8
Xoutput2 net2 FrameData_O[10] VPWR VGND sg13g2_buf_1
XFILLER_10_379 VPWR VGND sg13g2_decap_8
XFILLER_10_302 VPWR VGND sg13g2_decap_8
XFILLER_6_328 VPWR VGND sg13g2_decap_8
XFILLER_9_133 VPWR VGND sg13g2_decap_8
XFILLER_5_350 VPWR VGND sg13g2_decap_8
XFILLER_3_63 VPWR VGND sg13g2_decap_8
X_083_ S4END[4] net75 VPWR VGND sg13g2_buf_1
XFILLER_6_147 VPWR VGND sg13g2_decap_8
XFILLER_5_0 VPWR VGND sg13g2_decap_8
XFILLER_2_342 VPWR VGND sg13g2_decap_8
XFILLER_9_84 VPWR VGND sg13g2_decap_8
XFILLER_7_467 VPWR VGND sg13g2_decap_8
X_066_ S2END[5] net67 VPWR VGND sg13g2_buf_1
XFILLER_0_42 VPWR VGND sg13g2_decap_8
XFILLER_2_161 VPWR VGND sg13g2_decap_8
XFILLER_4_448 VPWR VGND sg13g2_decap_8
XFILLER_7_286 VPWR VGND sg13g2_fill_1
XFILLER_7_231 VPWR VGND sg13g2_decap_8
X_049_ FrameStrobe[17] net41 VPWR VGND sg13g2_buf_1
XFILLER_1_429 VPWR VGND sg13g2_decap_8
XFILLER_0_462 VPWR VGND sg13g2_decap_8
XFILLER_4_245 VPWR VGND sg13g2_decap_8
XFILLER_6_63 VPWR VGND sg13g2_decap_8
XFILLER_10_517 VPWR VGND sg13g2_fill_2
XFILLER_9_7 VPWR VGND sg13g2_decap_8
XFILLER_9_359 VPWR VGND sg13g2_decap_8
Xoutput93 net93 NN4BEG[13] VPWR VGND sg13g2_buf_1
Xoutput82 net82 N4BEG[3] VPWR VGND sg13g2_buf_1
Xoutput71 net71 N2BEGb[6] VPWR VGND sg13g2_buf_1
Xoutput60 net60 N2BEG[3] VPWR VGND sg13g2_buf_1
Xoutput3 net3 FrameData_O[11] VPWR VGND sg13g2_buf_1
XFILLER_10_358 VPWR VGND sg13g2_decap_8
XFILLER_6_307 VPWR VGND sg13g2_decap_8
XFILLER_9_189 VPWR VGND sg13g2_decap_8
XFILLER_9_112 VPWR VGND sg13g2_decap_8
XFILLER_3_42 VPWR VGND sg13g2_decap_8
X_082_ S4END[5] net74 VPWR VGND sg13g2_buf_1
XFILLER_6_126 VPWR VGND sg13g2_decap_8
XFILLER_2_321 VPWR VGND sg13g2_decap_8
XFILLER_2_398 VPWR VGND sg13g2_decap_8
X_065_ S2END[6] net66 VPWR VGND sg13g2_buf_1
XFILLER_7_446 VPWR VGND sg13g2_decap_8
XFILLER_0_98 VPWR VGND sg13g2_decap_8
XFILLER_0_21 VPWR VGND sg13g2_decap_8
XFILLER_2_140 VPWR VGND sg13g2_decap_8
XFILLER_9_63 VPWR VGND sg13g2_decap_8
XFILLER_7_210 VPWR VGND sg13g2_decap_8
XFILLER_4_427 VPWR VGND sg13g2_decap_8
XFILLER_7_298 VPWR VGND sg13g2_decap_8
X_048_ FrameStrobe[16] net40 VPWR VGND sg13g2_buf_1
XFILLER_1_408 VPWR VGND sg13g2_decap_8
XFILLER_3_493 VPWR VGND sg13g2_decap_8
XFILLER_4_224 VPWR VGND sg13g2_decap_8
XFILLER_6_42 VPWR VGND sg13g2_decap_8
XFILLER_0_441 VPWR VGND sg13g2_decap_8
XFILLER_3_290 VPWR VGND sg13g2_decap_8
XFILLER_1_249 VPWR VGND sg13g2_fill_1
XFILLER_1_238 VPWR VGND sg13g2_decap_8
Xoutput50 net50 FrameStrobe_O[7] VPWR VGND sg13g2_buf_1
XFILLER_9_338 VPWR VGND sg13g2_decap_8
XFILLER_9_305 VPWR VGND sg13g2_decap_8
Xoutput94 net94 NN4BEG[14] VPWR VGND sg13g2_buf_1
Xoutput83 net83 N4BEG[4] VPWR VGND sg13g2_buf_1
Xoutput72 net72 N2BEGb[7] VPWR VGND sg13g2_buf_1
Xoutput61 net61 N2BEG[4] VPWR VGND sg13g2_buf_1
XFILLER_5_522 VPWR VGND sg13g2_fill_1
XFILLER_5_511 VPWR VGND sg13g2_decap_8
Xoutput4 net4 FrameData_O[12] VPWR VGND sg13g2_buf_1
XFILLER_10_337 VPWR VGND sg13g2_decap_8
XFILLER_2_503 VPWR VGND sg13g2_decap_8
XFILLER_9_168 VPWR VGND sg13g2_decap_8
XFILLER_5_385 VPWR VGND sg13g2_decap_8
XFILLER_3_21 VPWR VGND sg13g2_decap_8
XFILLER_3_98 VPWR VGND sg13g2_decap_8
X_081_ S4END[6] net88 VPWR VGND sg13g2_buf_1
XFILLER_6_105 VPWR VGND sg13g2_decap_8
XFILLER_2_300 VPWR VGND sg13g2_decap_8
XFILLER_5_182 VPWR VGND sg13g2_decap_8
XFILLER_2_377 VPWR VGND sg13g2_decap_8
XFILLER_3_119 VPWR VGND sg13g2_decap_8
X_064_ S2END[7] net65 VPWR VGND sg13g2_buf_1
XFILLER_7_425 VPWR VGND sg13g2_decap_8
XFILLER_2_196 VPWR VGND sg13g2_decap_8
XFILLER_9_42 VPWR VGND sg13g2_decap_8
XFILLER_0_77 VPWR VGND sg13g2_decap_8
XFILLER_4_406 VPWR VGND sg13g2_decap_8
XFILLER_7_277 VPWR VGND sg13g2_decap_8
XFILLER_7_266 VPWR VGND sg13g2_fill_2
X_047_ FrameStrobe[15] net39 VPWR VGND sg13g2_buf_1
XFILLER_3_472 VPWR VGND sg13g2_decap_8
XFILLER_4_203 VPWR VGND sg13g2_decap_8
XFILLER_6_98 VPWR VGND sg13g2_decap_8
XFILLER_6_21 VPWR VGND sg13g2_decap_8
XFILLER_0_420 VPWR VGND sg13g2_decap_8
XFILLER_0_497 VPWR VGND sg13g2_decap_8
XFILLER_1_217 VPWR VGND sg13g2_decap_8
Xoutput40 net40 FrameStrobe_O[16] VPWR VGND sg13g2_buf_1
Xoutput51 net51 FrameStrobe_O[8] VPWR VGND sg13g2_buf_1
XFILLER_9_317 VPWR VGND sg13g2_decap_8
Xoutput95 net95 NN4BEG[15] VPWR VGND sg13g2_buf_1
Xoutput84 net84 N4BEG[5] VPWR VGND sg13g2_buf_1
Xoutput73 net73 N4BEG[0] VPWR VGND sg13g2_buf_1
Xoutput62 net62 N2BEG[5] VPWR VGND sg13g2_buf_1
Xoutput5 net5 FrameData_O[13] VPWR VGND sg13g2_buf_1
XFILLER_0_294 VPWR VGND sg13g2_decap_8
XFILLER_10_316 VPWR VGND sg13g2_decap_8
XFILLER_9_147 VPWR VGND sg13g2_decap_8
XFILLER_5_364 VPWR VGND sg13g2_decap_8
XFILLER_3_77 VPWR VGND sg13g2_decap_8
X_080_ S4END[7] net87 VPWR VGND sg13g2_buf_1
XFILLER_2_356 VPWR VGND sg13g2_decap_8
XFILLER_5_161 VPWR VGND sg13g2_decap_8
X_063_ S2MID[0] net64 VPWR VGND sg13g2_buf_1
XFILLER_7_404 VPWR VGND sg13g2_decap_8
XFILLER_2_175 VPWR VGND sg13g2_decap_8
XFILLER_3_0 VPWR VGND sg13g2_decap_8
XFILLER_9_98 VPWR VGND sg13g2_decap_8
XFILLER_9_21 VPWR VGND sg13g2_decap_8
XFILLER_6_481 VPWR VGND sg13g2_decap_8
XFILLER_0_56 VPWR VGND sg13g2_decap_8
X_046_ FrameStrobe[14] net38 VPWR VGND sg13g2_buf_1
XFILLER_7_245 VPWR VGND sg13g2_decap_8
XFILLER_3_451 VPWR VGND sg13g2_decap_8
XFILLER_0_476 VPWR VGND sg13g2_decap_8
XFILLER_4_259 VPWR VGND sg13g2_decap_8
X_029_ FrameData[29] net22 VPWR VGND sg13g2_buf_1
XFILLER_6_77 VPWR VGND sg13g2_decap_8
Xoutput41 net41 FrameStrobe_O[17] VPWR VGND sg13g2_buf_1
Xoutput52 net52 FrameStrobe_O[9] VPWR VGND sg13g2_buf_1
Xoutput6 net6 FrameData_O[14] VPWR VGND sg13g2_buf_1
Xoutput30 net30 FrameData_O[7] VPWR VGND sg13g2_buf_1
Xoutput96 net96 NN4BEG[1] VPWR VGND sg13g2_buf_1
Xoutput74 net74 N4BEG[10] VPWR VGND sg13g2_buf_1
Xoutput85 net85 N4BEG[6] VPWR VGND sg13g2_buf_1
Xoutput63 net63 N2BEG[6] VPWR VGND sg13g2_buf_1
XFILLER_0_273 VPWR VGND sg13g2_decap_8
.ends

