module N_term_DSP (UserCLK,
    UserCLKo,
    VPWR,
    VGND,
    FrameData,
    FrameData_O,
    FrameStrobe,
    FrameStrobe_O,
    N1END,
    N2END,
    N2MID,
    N4END,
    NN4END,
    S1BEG,
    S2BEG,
    S2BEGb,
    S4BEG,
    SS4BEG);
 input UserCLK;
 output UserCLKo;
 inout VPWR;
 inout VGND;
 input [31:0] FrameData;
 output [31:0] FrameData_O;
 input [19:0] FrameStrobe;
 output [19:0] FrameStrobe_O;
 input [3:0] N1END;
 input [7:0] N2END;
 input [7:0] N2MID;
 input [15:0] N4END;
 input [15:0] NN4END;
 output [3:0] S1BEG;
 output [7:0] S2BEG;
 output [7:0] S2BEGb;
 output [15:0] S4BEG;
 output [15:0] SS4BEG;

 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;

 sg13g2_buf_1 _000_ (.A(FrameData[0]),
    .X(net1),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _001_ (.A(FrameData[1]),
    .X(net12),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _002_ (.A(FrameData[2]),
    .X(net23),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _003_ (.A(FrameData[3]),
    .X(net26),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _004_ (.A(FrameData[4]),
    .X(net27),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _005_ (.A(FrameData[5]),
    .X(net28),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _006_ (.A(FrameData[6]),
    .X(net29),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _007_ (.A(FrameData[7]),
    .X(net30),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _008_ (.A(FrameData[8]),
    .X(net31),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _009_ (.A(FrameData[9]),
    .X(net32),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _010_ (.A(FrameData[10]),
    .X(net2),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _011_ (.A(FrameData[11]),
    .X(net3),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _012_ (.A(FrameData[12]),
    .X(net4),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _013_ (.A(FrameData[13]),
    .X(net5),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _014_ (.A(FrameData[14]),
    .X(net6),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _015_ (.A(FrameData[15]),
    .X(net7),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _016_ (.A(FrameData[16]),
    .X(net8),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _017_ (.A(FrameData[17]),
    .X(net9),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _018_ (.A(FrameData[18]),
    .X(net10),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _019_ (.A(FrameData[19]),
    .X(net11),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _020_ (.A(FrameData[20]),
    .X(net13),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _021_ (.A(FrameData[21]),
    .X(net14),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _022_ (.A(FrameData[22]),
    .X(net15),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _023_ (.A(FrameData[23]),
    .X(net16),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _024_ (.A(FrameData[24]),
    .X(net17),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _025_ (.A(FrameData[25]),
    .X(net18),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _026_ (.A(FrameData[26]),
    .X(net19),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _027_ (.A(FrameData[27]),
    .X(net20),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _028_ (.A(FrameData[28]),
    .X(net21),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _029_ (.A(FrameData[29]),
    .X(net22),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _030_ (.A(FrameData[30]),
    .X(net24),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _031_ (.A(FrameData[31]),
    .X(net25),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _032_ (.A(FrameStrobe[0]),
    .X(net33),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _033_ (.A(FrameStrobe[1]),
    .X(net44),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _034_ (.A(FrameStrobe[2]),
    .X(net45),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _035_ (.A(FrameStrobe[3]),
    .X(net46),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _036_ (.A(FrameStrobe[4]),
    .X(net47),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _037_ (.A(FrameStrobe[5]),
    .X(net48),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _038_ (.A(FrameStrobe[6]),
    .X(net49),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _039_ (.A(FrameStrobe[7]),
    .X(net50),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _040_ (.A(FrameStrobe[8]),
    .X(net51),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _041_ (.A(FrameStrobe[9]),
    .X(net52),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _042_ (.A(FrameStrobe[10]),
    .X(net34),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _043_ (.A(FrameStrobe[11]),
    .X(net35),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _044_ (.A(FrameStrobe[12]),
    .X(net36),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _045_ (.A(FrameStrobe[13]),
    .X(net37),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _046_ (.A(FrameStrobe[14]),
    .X(net38),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _047_ (.A(FrameStrobe[15]),
    .X(net39),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _048_ (.A(FrameStrobe[16]),
    .X(net40),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _049_ (.A(FrameStrobe[17]),
    .X(net41),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _050_ (.A(FrameStrobe[18]),
    .X(net42),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _051_ (.A(FrameStrobe[19]),
    .X(net43),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _052_ (.A(N1END[3]),
    .X(net53),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _053_ (.A(N1END[2]),
    .X(net54),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _054_ (.A(N1END[1]),
    .X(net55),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _055_ (.A(N1END[0]),
    .X(net56),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _056_ (.A(N2MID[7]),
    .X(net57),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _057_ (.A(N2MID[6]),
    .X(net58),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _058_ (.A(N2MID[5]),
    .X(net59),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _059_ (.A(N2MID[4]),
    .X(net60),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _060_ (.A(N2MID[3]),
    .X(net61),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _061_ (.A(N2MID[2]),
    .X(net62),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _062_ (.A(N2MID[1]),
    .X(net63),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _063_ (.A(N2MID[0]),
    .X(net64),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _064_ (.A(N2END[7]),
    .X(net65),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _065_ (.A(N2END[6]),
    .X(net66),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _066_ (.A(N2END[5]),
    .X(net67),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _067_ (.A(N2END[4]),
    .X(net68),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _068_ (.A(N2END[3]),
    .X(net69),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _069_ (.A(N2END[2]),
    .X(net70),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _070_ (.A(N2END[1]),
    .X(net71),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _071_ (.A(N2END[0]),
    .X(net72),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _072_ (.A(N4END[15]),
    .X(net73),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _073_ (.A(N4END[14]),
    .X(net80),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _074_ (.A(N4END[13]),
    .X(net81),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _075_ (.A(N4END[12]),
    .X(net82),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _076_ (.A(N4END[11]),
    .X(net83),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _077_ (.A(N4END[10]),
    .X(net84),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _078_ (.A(N4END[9]),
    .X(net85),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _079_ (.A(N4END[8]),
    .X(net86),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _080_ (.A(N4END[7]),
    .X(net87),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _081_ (.A(N4END[6]),
    .X(net88),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _082_ (.A(N4END[5]),
    .X(net74),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _083_ (.A(N4END[4]),
    .X(net75),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _084_ (.A(N4END[3]),
    .X(net76),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _085_ (.A(N4END[2]),
    .X(net77),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _086_ (.A(N4END[1]),
    .X(net78),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _087_ (.A(N4END[0]),
    .X(net79),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _088_ (.A(NN4END[15]),
    .X(net89),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _089_ (.A(NN4END[14]),
    .X(net96),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _090_ (.A(NN4END[13]),
    .X(net97),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _091_ (.A(NN4END[12]),
    .X(net98),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _092_ (.A(NN4END[11]),
    .X(net99),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _093_ (.A(NN4END[10]),
    .X(net100),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _094_ (.A(NN4END[9]),
    .X(net101),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _095_ (.A(NN4END[8]),
    .X(net102),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _096_ (.A(NN4END[7]),
    .X(net103),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _097_ (.A(NN4END[6]),
    .X(net104),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _098_ (.A(NN4END[5]),
    .X(net90),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _099_ (.A(NN4END[4]),
    .X(net91),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _100_ (.A(NN4END[3]),
    .X(net92),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _101_ (.A(NN4END[2]),
    .X(net93),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _102_ (.A(NN4END[1]),
    .X(net94),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _103_ (.A(NN4END[0]),
    .X(net95),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _104_ (.A(UserCLK),
    .X(net105),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output1 (.A(net1),
    .X(FrameData_O[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output2 (.A(net2),
    .X(FrameData_O[10]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output3 (.A(net3),
    .X(FrameData_O[11]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output4 (.A(net4),
    .X(FrameData_O[12]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output5 (.A(net5),
    .X(FrameData_O[13]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output6 (.A(net6),
    .X(FrameData_O[14]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output7 (.A(net7),
    .X(FrameData_O[15]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output8 (.A(net8),
    .X(FrameData_O[16]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output9 (.A(net9),
    .X(FrameData_O[17]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output10 (.A(net10),
    .X(FrameData_O[18]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output11 (.A(net11),
    .X(FrameData_O[19]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output12 (.A(net12),
    .X(FrameData_O[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output13 (.A(net13),
    .X(FrameData_O[20]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output14 (.A(net14),
    .X(FrameData_O[21]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output15 (.A(net15),
    .X(FrameData_O[22]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output16 (.A(net16),
    .X(FrameData_O[23]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output17 (.A(net17),
    .X(FrameData_O[24]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output18 (.A(net18),
    .X(FrameData_O[25]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output19 (.A(net19),
    .X(FrameData_O[26]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output20 (.A(net20),
    .X(FrameData_O[27]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output21 (.A(net21),
    .X(FrameData_O[28]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output22 (.A(net22),
    .X(FrameData_O[29]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output23 (.A(net23),
    .X(FrameData_O[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output24 (.A(net24),
    .X(FrameData_O[30]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output25 (.A(net25),
    .X(FrameData_O[31]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output26 (.A(net26),
    .X(FrameData_O[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output27 (.A(net27),
    .X(FrameData_O[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output28 (.A(net28),
    .X(FrameData_O[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output29 (.A(net29),
    .X(FrameData_O[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output30 (.A(net30),
    .X(FrameData_O[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output31 (.A(net31),
    .X(FrameData_O[8]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output32 (.A(net32),
    .X(FrameData_O[9]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output33 (.A(net33),
    .X(FrameStrobe_O[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output34 (.A(net34),
    .X(FrameStrobe_O[10]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output35 (.A(net35),
    .X(FrameStrobe_O[11]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output36 (.A(net36),
    .X(FrameStrobe_O[12]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output37 (.A(net37),
    .X(FrameStrobe_O[13]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output38 (.A(net38),
    .X(FrameStrobe_O[14]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output39 (.A(net39),
    .X(FrameStrobe_O[15]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output40 (.A(net40),
    .X(FrameStrobe_O[16]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output41 (.A(net41),
    .X(FrameStrobe_O[17]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output42 (.A(net42),
    .X(FrameStrobe_O[18]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output43 (.A(net43),
    .X(FrameStrobe_O[19]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output44 (.A(net44),
    .X(FrameStrobe_O[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output45 (.A(net45),
    .X(FrameStrobe_O[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output46 (.A(net46),
    .X(FrameStrobe_O[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output47 (.A(net47),
    .X(FrameStrobe_O[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output48 (.A(net48),
    .X(FrameStrobe_O[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output49 (.A(net49),
    .X(FrameStrobe_O[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output50 (.A(net50),
    .X(FrameStrobe_O[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output51 (.A(net51),
    .X(FrameStrobe_O[8]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output52 (.A(net52),
    .X(FrameStrobe_O[9]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output53 (.A(net53),
    .X(S1BEG[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output54 (.A(net54),
    .X(S1BEG[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output55 (.A(net55),
    .X(S1BEG[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output56 (.A(net56),
    .X(S1BEG[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output57 (.A(net57),
    .X(S2BEG[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output58 (.A(net58),
    .X(S2BEG[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output59 (.A(net59),
    .X(S2BEG[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output60 (.A(net60),
    .X(S2BEG[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output61 (.A(net61),
    .X(S2BEG[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output62 (.A(net62),
    .X(S2BEG[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output63 (.A(net63),
    .X(S2BEG[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output64 (.A(net64),
    .X(S2BEG[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output65 (.A(net65),
    .X(S2BEGb[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output66 (.A(net66),
    .X(S2BEGb[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output67 (.A(net67),
    .X(S2BEGb[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output68 (.A(net68),
    .X(S2BEGb[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output69 (.A(net69),
    .X(S2BEGb[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output70 (.A(net70),
    .X(S2BEGb[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output71 (.A(net71),
    .X(S2BEGb[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output72 (.A(net72),
    .X(S2BEGb[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output73 (.A(net73),
    .X(S4BEG[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output74 (.A(net74),
    .X(S4BEG[10]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output75 (.A(net75),
    .X(S4BEG[11]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output76 (.A(net76),
    .X(S4BEG[12]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output77 (.A(net77),
    .X(S4BEG[13]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output78 (.A(net78),
    .X(S4BEG[14]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output79 (.A(net79),
    .X(S4BEG[15]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output80 (.A(net80),
    .X(S4BEG[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output81 (.A(net81),
    .X(S4BEG[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output82 (.A(net82),
    .X(S4BEG[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output83 (.A(net83),
    .X(S4BEG[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output84 (.A(net84),
    .X(S4BEG[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output85 (.A(net85),
    .X(S4BEG[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output86 (.A(net86),
    .X(S4BEG[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output87 (.A(net87),
    .X(S4BEG[8]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output88 (.A(net88),
    .X(S4BEG[9]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output89 (.A(net89),
    .X(SS4BEG[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output90 (.A(net90),
    .X(SS4BEG[10]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output91 (.A(net91),
    .X(SS4BEG[11]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output92 (.A(net92),
    .X(SS4BEG[12]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output93 (.A(net93),
    .X(SS4BEG[13]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output94 (.A(net94),
    .X(SS4BEG[14]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output95 (.A(net95),
    .X(SS4BEG[15]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output96 (.A(net96),
    .X(SS4BEG[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output97 (.A(net97),
    .X(SS4BEG[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output98 (.A(net98),
    .X(SS4BEG[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output99 (.A(net99),
    .X(SS4BEG[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output100 (.A(net100),
    .X(SS4BEG[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output101 (.A(net101),
    .X(SS4BEG[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output102 (.A(net102),
    .X(SS4BEG[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output103 (.A(net103),
    .X(SS4BEG[8]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output104 (.A(net104),
    .X(SS4BEG[9]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output105 (.A(net105),
    .X(UserCLKo),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_341 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_265 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_293 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_90 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_370 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_71 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_97 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_19 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_26 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_341 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_19 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_26 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_52 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_59 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_66 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_73 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_80 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_136 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_157 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_164 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_171 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_178 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_227 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_265 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_58 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_65 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_69 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_136 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_265 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_15 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_22 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_51 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_58 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_69 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_328 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_375 (.VDD(VPWR),
    .VSS(VGND));
endmodule
