* NGSPICE file created from LUT4AB.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlxtp_1 abstract view
.subckt sky130_fd_sc_hd__dlxtp_1 D GATE VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_1 abstract view
.subckt sky130_fd_sc_hd__inv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd1_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd1_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

.subckt LUT4AB Ci Co E1BEG[0] E1BEG[1] E1BEG[2] E1BEG[3] E1END[0] E1END[1] E1END[2]
+ E1END[3] E2BEG[0] E2BEG[1] E2BEG[2] E2BEG[3] E2BEG[4] E2BEG[5] E2BEG[6] E2BEG[7]
+ E2BEGb[0] E2BEGb[1] E2BEGb[2] E2BEGb[3] E2BEGb[4] E2BEGb[5] E2BEGb[6] E2BEGb[7]
+ E2END[0] E2END[1] E2END[2] E2END[3] E2END[4] E2END[5] E2END[6] E2END[7] E2MID[0]
+ E2MID[1] E2MID[2] E2MID[3] E2MID[4] E2MID[5] E2MID[6] E2MID[7] E6BEG[0] E6BEG[10]
+ E6BEG[11] E6BEG[1] E6BEG[2] E6BEG[3] E6BEG[4] E6BEG[5] E6BEG[6] E6BEG[7] E6BEG[8]
+ E6BEG[9] E6END[0] E6END[10] E6END[11] E6END[1] E6END[2] E6END[3] E6END[4] E6END[5]
+ E6END[6] E6END[7] E6END[8] E6END[9] EE4BEG[0] EE4BEG[10] EE4BEG[11] EE4BEG[12] EE4BEG[13]
+ EE4BEG[14] EE4BEG[15] EE4BEG[1] EE4BEG[2] EE4BEG[3] EE4BEG[4] EE4BEG[5] EE4BEG[6]
+ EE4BEG[7] EE4BEG[8] EE4BEG[9] EE4END[0] EE4END[10] EE4END[11] EE4END[12] EE4END[13]
+ EE4END[14] EE4END[15] EE4END[1] EE4END[2] EE4END[3] EE4END[4] EE4END[5] EE4END[6]
+ EE4END[7] EE4END[8] EE4END[9] FrameData[0] FrameData[10] FrameData[11] FrameData[12]
+ FrameData[13] FrameData[14] FrameData[15] FrameData[16] FrameData[17] FrameData[18]
+ FrameData[19] FrameData[1] FrameData[20] FrameData[21] FrameData[22] FrameData[23]
+ FrameData[24] FrameData[25] FrameData[26] FrameData[27] FrameData[28] FrameData[29]
+ FrameData[2] FrameData[30] FrameData[31] FrameData[3] FrameData[4] FrameData[5]
+ FrameData[6] FrameData[7] FrameData[8] FrameData[9] FrameData_O[0] FrameData_O[10]
+ FrameData_O[11] FrameData_O[12] FrameData_O[13] FrameData_O[14] FrameData_O[15]
+ FrameData_O[16] FrameData_O[17] FrameData_O[18] FrameData_O[19] FrameData_O[1] FrameData_O[20]
+ FrameData_O[21] FrameData_O[22] FrameData_O[23] FrameData_O[24] FrameData_O[25]
+ FrameData_O[26] FrameData_O[27] FrameData_O[28] FrameData_O[29] FrameData_O[2] FrameData_O[30]
+ FrameData_O[31] FrameData_O[3] FrameData_O[4] FrameData_O[5] FrameData_O[6] FrameData_O[7]
+ FrameData_O[8] FrameData_O[9] FrameStrobe[0] FrameStrobe[10] FrameStrobe[11] FrameStrobe[12]
+ FrameStrobe[13] FrameStrobe[14] FrameStrobe[15] FrameStrobe[16] FrameStrobe[17]
+ FrameStrobe[18] FrameStrobe[19] FrameStrobe[1] FrameStrobe[2] FrameStrobe[3] FrameStrobe[4]
+ FrameStrobe[5] FrameStrobe[6] FrameStrobe[7] FrameStrobe[8] FrameStrobe[9] FrameStrobe_O[0]
+ FrameStrobe_O[10] FrameStrobe_O[11] FrameStrobe_O[12] FrameStrobe_O[13] FrameStrobe_O[14]
+ FrameStrobe_O[15] FrameStrobe_O[16] FrameStrobe_O[17] FrameStrobe_O[18] FrameStrobe_O[19]
+ FrameStrobe_O[1] FrameStrobe_O[2] FrameStrobe_O[3] FrameStrobe_O[4] FrameStrobe_O[5]
+ FrameStrobe_O[6] FrameStrobe_O[7] FrameStrobe_O[8] FrameStrobe_O[9] N1BEG[0] N1BEG[1]
+ N1BEG[2] N1BEG[3] N1END[0] N1END[1] N1END[2] N1END[3] N2BEG[0] N2BEG[1] N2BEG[2]
+ N2BEG[3] N2BEG[4] N2BEG[5] N2BEG[6] N2BEG[7] N2BEGb[0] N2BEGb[1] N2BEGb[2] N2BEGb[3]
+ N2BEGb[4] N2BEGb[5] N2BEGb[6] N2BEGb[7] N2END[0] N2END[1] N2END[2] N2END[3] N2END[4]
+ N2END[5] N2END[6] N2END[7] N2MID[0] N2MID[1] N2MID[2] N2MID[3] N2MID[4] N2MID[5]
+ N2MID[6] N2MID[7] N4BEG[0] N4BEG[10] N4BEG[11] N4BEG[12] N4BEG[13] N4BEG[14] N4BEG[15]
+ N4BEG[1] N4BEG[2] N4BEG[3] N4BEG[4] N4BEG[5] N4BEG[6] N4BEG[7] N4BEG[8] N4BEG[9]
+ N4END[0] N4END[10] N4END[11] N4END[12] N4END[13] N4END[14] N4END[15] N4END[1] N4END[2]
+ N4END[3] N4END[4] N4END[5] N4END[6] N4END[7] N4END[8] N4END[9] NN4BEG[0] NN4BEG[10]
+ NN4BEG[11] NN4BEG[12] NN4BEG[13] NN4BEG[14] NN4BEG[15] NN4BEG[1] NN4BEG[2] NN4BEG[3]
+ NN4BEG[4] NN4BEG[5] NN4BEG[6] NN4BEG[7] NN4BEG[8] NN4BEG[9] NN4END[0] NN4END[10]
+ NN4END[11] NN4END[12] NN4END[13] NN4END[14] NN4END[15] NN4END[1] NN4END[2] NN4END[3]
+ NN4END[4] NN4END[5] NN4END[6] NN4END[7] NN4END[8] NN4END[9] S1BEG[0] S1BEG[1] S1BEG[2]
+ S1BEG[3] S1END[0] S1END[1] S1END[2] S1END[3] S2BEG[0] S2BEG[1] S2BEG[2] S2BEG[3]
+ S2BEG[4] S2BEG[5] S2BEG[6] S2BEG[7] S2BEGb[0] S2BEGb[1] S2BEGb[2] S2BEGb[3] S2BEGb[4]
+ S2BEGb[5] S2BEGb[6] S2BEGb[7] S2END[0] S2END[1] S2END[2] S2END[3] S2END[4] S2END[5]
+ S2END[6] S2END[7] S2MID[0] S2MID[1] S2MID[2] S2MID[3] S2MID[4] S2MID[5] S2MID[6]
+ S2MID[7] S4BEG[0] S4BEG[10] S4BEG[11] S4BEG[12] S4BEG[13] S4BEG[14] S4BEG[15] S4BEG[1]
+ S4BEG[2] S4BEG[3] S4BEG[4] S4BEG[5] S4BEG[6] S4BEG[7] S4BEG[8] S4BEG[9] S4END[0]
+ S4END[10] S4END[11] S4END[12] S4END[13] S4END[14] S4END[15] S4END[1] S4END[2] S4END[3]
+ S4END[4] S4END[5] S4END[6] S4END[7] S4END[8] S4END[9] SS4BEG[0] SS4BEG[10] SS4BEG[11]
+ SS4BEG[12] SS4BEG[13] SS4BEG[14] SS4BEG[15] SS4BEG[1] SS4BEG[2] SS4BEG[3] SS4BEG[4]
+ SS4BEG[5] SS4BEG[6] SS4BEG[7] SS4BEG[8] SS4BEG[9] SS4END[0] SS4END[10] SS4END[11]
+ SS4END[12] SS4END[13] SS4END[14] SS4END[15] SS4END[1] SS4END[2] SS4END[3] SS4END[4]
+ SS4END[5] SS4END[6] SS4END[7] SS4END[8] SS4END[9] UserCLK UserCLKo VGND VPWR W1BEG[0]
+ W1BEG[1] W1BEG[2] W1BEG[3] W1END[0] W1END[1] W1END[2] W1END[3] W2BEG[0] W2BEG[1]
+ W2BEG[2] W2BEG[3] W2BEG[4] W2BEG[5] W2BEG[6] W2BEG[7] W2BEGb[0] W2BEGb[1] W2BEGb[2]
+ W2BEGb[3] W2BEGb[4] W2BEGb[5] W2BEGb[6] W2BEGb[7] W2END[0] W2END[1] W2END[2] W2END[3]
+ W2END[4] W2END[5] W2END[6] W2END[7] W2MID[0] W2MID[1] W2MID[2] W2MID[3] W2MID[4]
+ W2MID[5] W2MID[6] W2MID[7] W6BEG[0] W6BEG[10] W6BEG[11] W6BEG[1] W6BEG[2] W6BEG[3]
+ W6BEG[4] W6BEG[5] W6BEG[6] W6BEG[7] W6BEG[8] W6BEG[9] W6END[0] W6END[10] W6END[11]
+ W6END[1] W6END[2] W6END[3] W6END[4] W6END[5] W6END[6] W6END[7] W6END[8] W6END[9]
+ WW4BEG[0] WW4BEG[10] WW4BEG[11] WW4BEG[12] WW4BEG[13] WW4BEG[14] WW4BEG[15] WW4BEG[1]
+ WW4BEG[2] WW4BEG[3] WW4BEG[4] WW4BEG[5] WW4BEG[6] WW4BEG[7] WW4BEG[8] WW4BEG[9]
+ WW4END[0] WW4END[10] WW4END[11] WW4END[12] WW4END[13] WW4END[14] WW4END[15] WW4END[1]
+ WW4END[2] WW4END[3] WW4END[4] WW4END[5] WW4END[6] WW4END[7] WW4END[8] WW4END[9]
X_2106_ clknet_1_1__leaf_UserCLK_regs _0007_ VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.LUT_flop
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_39_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2037_ net766 net699 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_52_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_20_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1270_ net432 _0393_ _0391_ VGND VGND VPWR VPWR _0394_ sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_59_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_89 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1606_ net791 net719 VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9
+ sky130_fd_sc_hd__dlxtp_1
X_0985_ net83 net7 net90 net118 Inst_LUT4AB_ConfigMem.Inst_frame5_bit16.Q Inst_LUT4AB_ConfigMem.Inst_frame5_bit17.Q
+ VGND VGND VPWR VPWR _0130_ sky130_fd_sc_hd__mux4_2
X_1399_ net60 net815 net665 net661 Inst_LUT4AB_ConfigMem.Inst_frame13_bit5.Q Inst_LUT4AB_ConfigMem.Inst_frame13_bit6.Q
+ VGND VGND VPWR VPWR _0499_ sky130_fd_sc_hd__mux4_1
X_1468_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit0.Q net621 _0535_ Inst_LD_LUT4c_frame_config_dffesr.c_reset_value
+ VGND VGND VPWR VPWR _0537_ sky130_fd_sc_hd__o2bb2a_1
X_1537_ net801 net711 VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.c_out_mux
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_27_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout661 net662 VGND VGND VPWR VPWR net661 sky130_fd_sc_hd__buf_2
Xfanout672 net673 VGND VGND VPWR VPWR net672 sky130_fd_sc_hd__buf_1
XFILLER_37_40 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout683 net686 VGND VGND VPWR VPWR net683 sky130_fd_sc_hd__clkbuf_2
Xfanout650 net651 VGND VGND VPWR VPWR net650 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_5_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout694 FrameStrobe[3] VGND VGND VPWR VPWR net694 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_56_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0770_ _0616_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit5.Q _0618_ VGND VGND VPWR VPWR
+ _0619_ sky130_fd_sc_hd__o21a_1
XFILLER_56_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1253_ _0378_ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.JW2BEG7 sky130_fd_sc_hd__inv_1
X_1322_ _0617_ _0053_ _0120_ net664 Inst_LUT4AB_ConfigMem.Inst_frame11_bit26.Q Inst_LUT4AB_ConfigMem.Inst_frame11_bit27.Q
+ VGND VGND VPWR VPWR _0439_ sky130_fd_sc_hd__mux4_1
X_1184_ Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 _0303_ _0307_ Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14
+ VGND VGND VPWR VPWR _0316_ sky130_fd_sc_hd__o22a_1
XFILLER_49_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_20_Left_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0968_ _0112_ _0113_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit16.Q VGND VGND VPWR VPWR
+ _0114_ sky130_fd_sc_hd__mux2_4
Xoutput231 net231 VGND VGND VPWR VPWR FrameStrobe_O[1] sky130_fd_sc_hd__buf_2
Xoutput220 net220 VGND VGND VPWR VPWR FrameStrobe_O[0] sky130_fd_sc_hd__buf_2
Xoutput253 net253 VGND VGND VPWR VPWR N2BEGb[1] sky130_fd_sc_hd__buf_2
Xoutput242 net242 VGND VGND VPWR VPWR N1BEG[2] sky130_fd_sc_hd__buf_4
Xoutput286 net286 VGND VGND VPWR VPWR NN4BEG[4] sky130_fd_sc_hd__buf_2
Xoutput275 net275 VGND VGND VPWR VPWR N4BEG[9] sky130_fd_sc_hd__buf_2
Xoutput264 Inst_LUT4AB_switch_matrix.N4BEG1 VGND VGND VPWR VPWR N4BEG[13] sky130_fd_sc_hd__buf_6
XFILLER_59_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0899_ net58 net66 net3 net11 Inst_LUT4AB_ConfigMem.Inst_frame3_bit10.Q Inst_LUT4AB_ConfigMem.Inst_frame3_bit11.Q
+ VGND VGND VPWR VPWR _0050_ sky130_fd_sc_hd__mux4_1
XFILLER_59_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput297 net297 VGND VGND VPWR VPWR S2BEG[1] sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_53_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1871_ net770 net675 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame7_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1940_ net790 net687 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0822_ net639 net629 net624 net623 Inst_LUT4AB_ConfigMem.Inst_frame1_bit6.Q Inst_LUT4AB_ConfigMem.Inst_frame1_bit7.Q
+ VGND VGND VPWR VPWR _0667_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_16_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0753_ _0602_ _0603_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit0.Q VGND VGND VPWR VPWR
+ _0604_ sky130_fd_sc_hd__mux2_1
X_2285_ S4END[10] VGND VGND VPWR VPWR net324 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_67_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1236_ _0363_ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.E2BEG7 sky130_fd_sc_hd__inv_6
XFILLER_56_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1305_ _0422_ _0423_ _0593_ VGND VGND VPWR VPWR _0424_ sky130_fd_sc_hd__mux2_1
X_2354_ WW4END[14] VGND VGND VPWR VPWR net378 sky130_fd_sc_hd__clkbuf_2
X_1098_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit20.Q _0234_ VGND VGND VPWR VPWR _0235_
+ sky130_fd_sc_hd__and2b_1
X_1167_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit10.Q _0297_ _0298_ Inst_LH_LUT4c_frame_config_dffesr.c_I0mux
+ _0296_ VGND VGND VPWR VPWR _0299_ sky130_fd_sc_hd__a311oi_1
XFILLER_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2070_ net759 net745 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame0_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_72_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1021_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit12.Q _0162_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit13.Q
+ VGND VGND VPWR VPWR _0163_ sky130_fd_sc_hd__a21bo_1
XFILLER_34_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1854_ net808 net677 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame7_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1785_ net753 net670 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1923_ net797 net683 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame5_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0805_ _0648_ _0646_ _0651_ _0558_ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.JS2BEG3
+ sky130_fd_sc_hd__a22o_1
X_0736_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit28.Q VGND VGND VPWR VPWR _0587_ sky130_fd_sc_hd__inv_1
X_2337_ W6END[7] VGND VGND VPWR VPWR net372 sky130_fd_sc_hd__clkbuf_2
X_2268_ net408 VGND VGND VPWR VPWR net301 sky130_fd_sc_hd__buf_2
X_2199_ net733 VGND VGND VPWR VPWR net223 sky130_fd_sc_hd__buf_1
X_1219_ _0341_ _0338_ _0347_ _0348_ VGND VGND VPWR VPWR _0349_ sky130_fd_sc_hd__a22o_1
XFILLER_25_301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_175 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_33_Left_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_42_Left_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_51_Left_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_5 net171 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_60_Left_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1570_ net799 net712 VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11
+ sky130_fd_sc_hd__dlxtp_1
X_2053_ net794 net701 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_66_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrebuffer17 _0354_ VGND VGND VPWR VPWR net409 sky130_fd_sc_hd__dlygate4sd1_1
XTAP_TAPCELL_ROW_49_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer39 _0107_ VGND VGND VPWR VPWR net431 sky130_fd_sc_hd__buf_6
X_2122_ net17 VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__clkbuf_2
X_1004_ Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 _0124_ _0126_ Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1
+ _0147_ VGND VGND VPWR VPWR _0148_ sky130_fd_sc_hd__o221a_1
X_1837_ net774 net674 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame8_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1906_ net761 net682 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame6_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1768_ net785 net739 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame10_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0719_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit17.Q VGND VGND VPWR VPWR _0570_ sky130_fd_sc_hd__inv_1
X_1699_ net797 net730 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame12_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_25_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_23_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_50 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput131 W2MID[6] VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__clkbuf_2
Xinput120 W2END[3] VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__buf_2
XFILLER_71_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1622_ net760 net723 VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6
+ sky130_fd_sc_hd__dlxtp_1
X_1553_ net46 net710 VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13
+ sky130_fd_sc_hd__dlxtp_1
X_1484_ net777 net55 VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1
+ sky130_fd_sc_hd__dlxtp_1
X_2105_ clknet_1_1__leaf_UserCLK_regs _0006_ VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.LUT_flop
+ sky130_fd_sc_hd__dfxtp_1
X_2036_ net790 net699 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_10_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout810 net29 VGND VGND VPWR VPWR net810 sky130_fd_sc_hd__clkbuf_4
XFILLER_45_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_134 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer8 Inst_LUT4AB_switch_matrix.JS2BEG7 VGND VGND VPWR VPWR net400 sky130_fd_sc_hd__clkbuf_2
XFILLER_42_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0984_ net27 net136 net105 Inst_LUT4AB_switch_matrix.JW2BEG3 Inst_LUT4AB_ConfigMem.Inst_frame0_bit17.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame0_bit16.Q VGND VGND VPWR VPWR _0129_ sky130_fd_sc_hd__mux4_2
X_1605_ net793 net718 VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8
+ sky130_fd_sc_hd__dlxtp_1
X_1536_ net804 net707 VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_8_171 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1398_ _0498_ _0497_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit10.Q VGND VGND VPWR VPWR
+ Inst_LUT4AB_switch_matrix.NN4BEG2 sky130_fd_sc_hd__mux2_1
X_1467_ _0349_ _0535_ VGND VGND VPWR VPWR _0536_ sky130_fd_sc_hd__nand2b_1
X_2019_ net797 net697 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_35_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_66 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout640 net643 VGND VGND VPWR VPWR net640 sky130_fd_sc_hd__buf_8
Xfanout651 C VGND VGND VPWR VPWR net651 sky130_fd_sc_hd__clkbuf_2
XFILLER_2_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_56_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout662 net663 VGND VGND VPWR VPWR net662 sky130_fd_sc_hd__clkbuf_2
Xfanout673 FrameStrobe[8] VGND VGND VPWR VPWR net673 sky130_fd_sc_hd__clkbuf_4
XFILLER_37_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_207 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout684 net686 VGND VGND VPWR VPWR net684 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_5_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout695 net696 VGND VGND VPWR VPWR net695 sky130_fd_sc_hd__clkbuf_2
X_1252_ _0585_ _0373_ _0375_ _0377_ VGND VGND VPWR VPWR _0378_ sky130_fd_sc_hd__a2bb2o_4
X_1321_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit28.Q _0433_ _0436_ _0437_ VGND VGND
+ VPWR VPWR _0438_ sky130_fd_sc_hd__o22a_1
X_1183_ _0300_ _0314_ _0311_ VGND VGND VPWR VPWR _0315_ sky130_fd_sc_hd__a21oi_1
XFILLER_64_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0967_ net646 net632 net410 net623 Inst_LUT4AB_ConfigMem.Inst_frame3_bit14.Q Inst_LUT4AB_ConfigMem.Inst_frame3_bit15.Q
+ VGND VGND VPWR VPWR _0113_ sky130_fd_sc_hd__mux4_2
Xoutput221 net221 VGND VGND VPWR VPWR FrameStrobe_O[10] sky130_fd_sc_hd__buf_2
Xoutput232 net232 VGND VGND VPWR VPWR FrameStrobe_O[2] sky130_fd_sc_hd__buf_2
Xoutput276 net276 VGND VGND VPWR VPWR NN4BEG[0] sky130_fd_sc_hd__buf_2
Xoutput265 Inst_LUT4AB_switch_matrix.N4BEG2 VGND VGND VPWR VPWR N4BEG[14] sky130_fd_sc_hd__buf_4
Xoutput243 net243 VGND VGND VPWR VPWR N1BEG[3] sky130_fd_sc_hd__buf_4
Xoutput287 net287 VGND VGND VPWR VPWR NN4BEG[5] sky130_fd_sc_hd__buf_2
Xoutput254 net254 VGND VGND VPWR VPWR N2BEGb[2] sky130_fd_sc_hd__buf_2
XFILLER_59_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput210 net210 VGND VGND VPWR VPWR FrameData_O[2] sky130_fd_sc_hd__buf_2
X_0898_ net86 net94 net88 net114 Inst_LUT4AB_ConfigMem.Inst_frame3_bit11.Q Inst_LUT4AB_ConfigMem.Inst_frame3_bit10.Q
+ VGND VGND VPWR VPWR _0049_ sky130_fd_sc_hd__mux4_1
Xoutput298 net298 VGND VGND VPWR VPWR S2BEG[2] sky130_fd_sc_hd__buf_6
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1519_ net769 net705 VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.c_I0mux
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_30_Right_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1870_ net771 net678 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame7_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0752_ net814 net91 net119 net138 Inst_LUT4AB_ConfigMem.Inst_frame4_bit30.Q Inst_LUT4AB_ConfigMem.Inst_frame4_bit31.Q
+ VGND VGND VPWR VPWR _0603_ sky130_fd_sc_hd__mux4_1
X_0821_ net426 net430 net649 net644 Inst_LUT4AB_ConfigMem.Inst_frame1_bit6.Q Inst_LUT4AB_ConfigMem.Inst_frame1_bit7.Q
+ VGND VGND VPWR VPWR _0666_ sky130_fd_sc_hd__mux4_2
XFILLER_14_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_16_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2353_ WW4END[13] VGND VGND VPWR VPWR net392 sky130_fd_sc_hd__clkbuf_2
X_2284_ S4END[9] VGND VGND VPWR VPWR net323 sky130_fd_sc_hd__clkbuf_2
X_1235_ _0583_ _0358_ _0360_ _0362_ VGND VGND VPWR VPWR _0363_ sky130_fd_sc_hd__a2bb2o_4
XTAP_TAPCELL_ROW_67_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1166_ _0581_ _0240_ VGND VGND VPWR VPWR _0298_ sky130_fd_sc_hd__nand2_1
X_1304_ net62 net815 net78 net7 Inst_LUT4AB_ConfigMem.Inst_frame5_bit27.Q Inst_LUT4AB_ConfigMem.Inst_frame5_bit26.Q
+ VGND VGND VPWR VPWR _0423_ sky130_fd_sc_hd__mux4_1
X_1097_ net60 net68 net815 net13 Inst_LUT4AB_ConfigMem.Inst_frame4_bit18.Q Inst_LUT4AB_ConfigMem.Inst_frame4_bit19.Q
+ VGND VGND VPWR VPWR _0234_ sky130_fd_sc_hd__mux4_1
XFILLER_52_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1999_ net770 net691 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_28_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_13_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_64_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1020_ net642 net631 net627 net623 Inst_LUT4AB_ConfigMem.Inst_frame4_bit10.Q Inst_LUT4AB_ConfigMem.Inst_frame4_bit11.Q
+ VGND VGND VPWR VPWR _0162_ sky130_fd_sc_hd__mux4_1
XFILLER_15_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1922_ net800 net685 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame5_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_34_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_29_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0735_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit25.Q VGND VGND VPWR VPWR _0586_ sky130_fd_sc_hd__inv_1
X_1853_ net810 net677 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame7_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1784_ net756 net670 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0804_ _0649_ _0650_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit8.Q VGND VGND VPWR VPWR
+ _0651_ sky130_fd_sc_hd__mux2_1
XFILLER_69_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2336_ W6END[6] VGND VGND VPWR VPWR net371 sky130_fd_sc_hd__clkbuf_2
X_2267_ Inst_LUT4AB_switch_matrix.JS2BEG4 VGND VGND VPWR VPWR net300 sky130_fd_sc_hd__clkbuf_2
XFILLER_37_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1218_ _0333_ _0344_ _0338_ VGND VGND VPWR VPWR _0348_ sky130_fd_sc_hd__a21oi_1
X_1149_ _0280_ _0281_ _0272_ _0271_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit5.Q Inst_LUT4AB_ConfigMem.Inst_frame8_bit6.Q
+ VGND VGND VPWR VPWR _0282_ sky130_fd_sc_hd__mux4_2
X_2198_ net738 VGND VGND VPWR VPWR net222 sky130_fd_sc_hd__clkbuf_2
XFILLER_25_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_206 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_26_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_6 E6END[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_73 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2052_ net795 net701 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_49_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1003_ Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 _0122_ _0125_ Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5
+ VGND VGND VPWR VPWR _0147_ sky130_fd_sc_hd__o22a_1
X_2121_ net16 VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__buf_1
XFILLER_30_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1905_ net763 net682 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame6_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1836_ net778 net673 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame8_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0718_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit17.Q VGND VGND VPWR VPWR _0569_ sky130_fd_sc_hd__inv_1
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1767_ net787 net740 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame10_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1698_ net800 net730 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame12_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_57_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2319_ Inst_LUT4AB_switch_matrix.JW2BEG3 VGND VGND VPWR VPWR net352 sky130_fd_sc_hd__clkbuf_1
XFILLER_25_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_23_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput110 SS4END[1] VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__buf_2
XFILLER_0_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput132 W2MID[7] VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput121 W2END[4] VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_59_Right_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1621_ net765 net723 VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5
+ sky130_fd_sc_hd__dlxtp_1
X_1552_ net768 net710 VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_68_Right_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2104_ clknet_1_1__leaf_UserCLK_regs _0005_ VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.LUT_flop
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_39_202 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1483_ net779 net55 VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_37_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2035_ net812 net699 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1819_ net749 net671 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame8_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
Xfanout800 net34 VGND VGND VPWR VPWR net800 sky130_fd_sc_hd__buf_4
Xfanout811 net812 VGND VGND VPWR VPWR net811 sky130_fd_sc_hd__buf_4
XFILLER_42_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_146 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer9 _0355_ VGND VGND VPWR VPWR net401 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_5_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0983_ Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 _0124_ _0126_ Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8
+ _0127_ VGND VGND VPWR VPWR _0128_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_42_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1604_ net796 net717 VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_8_183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1535_ net806 net707 VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_67_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1397_ net57 net113 net2 net658 Inst_LUT4AB_ConfigMem.Inst_frame13_bit9.Q Inst_LUT4AB_ConfigMem.Inst_frame13_bit8.Q
+ VGND VGND VPWR VPWR _0498_ sky130_fd_sc_hd__mux4_1
X_1466_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit9.Q _0522_ VGND VGND VPWR VPWR _0535_
+ sky130_fd_sc_hd__nand2_1
XFILLER_27_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2018_ net800 net697 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_12_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout652 net653 VGND VGND VPWR VPWR net652 sky130_fd_sc_hd__buf_2
Xfanout641 net642 VGND VGND VPWR VPWR net641 sky130_fd_sc_hd__buf_8
Xfanout630 G VGND VGND VPWR VPWR net630 sky130_fd_sc_hd__buf_8
Xfanout674 FrameStrobe[8] VGND VGND VPWR VPWR net674 sky130_fd_sc_hd__buf_2
Xfanout685 net686 VGND VGND VPWR VPWR net685 sky130_fd_sc_hd__buf_2
Xfanout663 A VGND VGND VPWR VPWR net663 sky130_fd_sc_hd__buf_8
XFILLER_58_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout696 FrameStrobe[2] VGND VGND VPWR VPWR net696 sky130_fd_sc_hd__clkbuf_2
XFILLER_33_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1320_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit27.Q _0434_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit28.Q
+ VGND VGND VPWR VPWR _0437_ sky130_fd_sc_hd__a21bo_1
X_1182_ _0312_ _0313_ VGND VGND VPWR VPWR _0314_ sky130_fd_sc_hd__nand2_1
X_1251_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit24.Q _0376_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit25.Q
+ VGND VGND VPWR VPWR _0377_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_62_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_19_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput200 net200 VGND VGND VPWR VPWR FrameData_O[20] sky130_fd_sc_hd__buf_2
X_0966_ net662 net656 net653 net636 Inst_LUT4AB_ConfigMem.Inst_frame3_bit14.Q Inst_LUT4AB_ConfigMem.Inst_frame3_bit15.Q
+ VGND VGND VPWR VPWR _0112_ sky130_fd_sc_hd__mux4_1
X_0897_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit12.Q _0047_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit13.Q
+ VGND VGND VPWR VPWR _0048_ sky130_fd_sc_hd__a21bo_1
Xoutput222 net222 VGND VGND VPWR VPWR FrameStrobe_O[11] sky130_fd_sc_hd__buf_2
Xoutput233 net233 VGND VGND VPWR VPWR FrameStrobe_O[3] sky130_fd_sc_hd__buf_2
Xoutput288 net288 VGND VGND VPWR VPWR NN4BEG[6] sky130_fd_sc_hd__buf_2
Xoutput277 net277 VGND VGND VPWR VPWR NN4BEG[10] sky130_fd_sc_hd__buf_2
Xoutput266 net266 VGND VGND VPWR VPWR N4BEG[15] sky130_fd_sc_hd__buf_4
Xoutput244 net244 VGND VGND VPWR VPWR N2BEG[0] sky130_fd_sc_hd__buf_6
Xoutput255 net255 VGND VGND VPWR VPWR N2BEGb[3] sky130_fd_sc_hd__buf_2
Xoutput211 net211 VGND VGND VPWR VPWR FrameData_O[30] sky130_fd_sc_hd__buf_2
XFILLER_59_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput299 net299 VGND VGND VPWR VPWR S2BEG[3] sky130_fd_sc_hd__buf_4
X_1518_ net771 net704 VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.c_out_mux
+ sky130_fd_sc_hd__dlxtp_1
X_1449_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit28.Q _0516_ _0521_ VGND VGND VPWR VPWR
+ _0522_ sky130_fd_sc_hd__o21a_4
XFILLER_70_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0751_ net57 net63 net79 net8 Inst_LUT4AB_ConfigMem.Inst_frame4_bit30.Q Inst_LUT4AB_ConfigMem.Inst_frame4_bit31.Q
+ VGND VGND VPWR VPWR _0602_ sky130_fd_sc_hd__mux4_1
X_0820_ _0664_ _0644_ _0620_ VGND VGND VPWR VPWR _0665_ sky130_fd_sc_hd__mux2_1
XFILLER_9_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2283_ S4END[8] VGND VGND VPWR VPWR net322 sky130_fd_sc_hd__clkbuf_2
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1303_ net813 net110 net118 net134 Inst_LUT4AB_ConfigMem.Inst_frame5_bit26.Q Inst_LUT4AB_ConfigMem.Inst_frame5_bit27.Q
+ VGND VGND VPWR VPWR _0422_ sky130_fd_sc_hd__mux4_1
X_2352_ WW4END[12] VGND VGND VPWR VPWR net391 sky130_fd_sc_hd__clkbuf_2
X_1096_ net88 net114 net96 net665 Inst_LUT4AB_ConfigMem.Inst_frame4_bit19.Q Inst_LUT4AB_ConfigMem.Inst_frame4_bit18.Q
+ VGND VGND VPWR VPWR _0233_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_67_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1234_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit24.Q _0361_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit25.Q
+ VGND VGND VPWR VPWR _0362_ sky130_fd_sc_hd__a21oi_1
XFILLER_64_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1165_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit9.Q _0239_ VGND VGND VPWR VPWR _0297_
+ sky130_fd_sc_hd__nand2_1
XFILLER_37_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0949_ _0092_ _0093_ _0095_ _0094_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit11.Q Inst_LUT4AB_ConfigMem.Inst_frame9_bit12.Q
+ VGND VGND VPWR VPWR _0096_ sky130_fd_sc_hd__mux4_1
X_1998_ net773 net691 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_7_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_72_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1921_ net802 net685 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame5_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1852_ net748 net675 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame7_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0734_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit25.Q VGND VGND VPWR VPWR _0585_ sky130_fd_sc_hd__inv_1
X_1783_ net757 net670 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_6_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_292 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0803_ net93 net121 net105 net137 Inst_LUT4AB_ConfigMem.Inst_frame2_bit7.Q Inst_LUT4AB_ConfigMem.Inst_frame2_bit6.Q
+ VGND VGND VPWR VPWR _0650_ sky130_fd_sc_hd__mux4_1
XFILLER_69_255 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2335_ W6END[5] VGND VGND VPWR VPWR net370 sky130_fd_sc_hd__clkbuf_2
X_2266_ Inst_LUT4AB_switch_matrix.JS2BEG3 VGND VGND VPWR VPWR net299 sky130_fd_sc_hd__clkbuf_2
X_1079_ _0215_ _0216_ VGND VGND VPWR VPWR _0217_ sky130_fd_sc_hd__or2_1
X_2197_ net742 VGND VGND VPWR VPWR net221 sky130_fd_sc_hd__buf_1
X_1217_ _0345_ _0346_ _0333_ VGND VGND VPWR VPWR _0347_ sky130_fd_sc_hd__a21o_1
X_1148_ net70 net15 net98 net126 Inst_LUT4AB_ConfigMem.Inst_frame6_bit24.Q Inst_LUT4AB_ConfigMem.Inst_frame6_bit25.Q
+ VGND VGND VPWR VPWR _0281_ sky130_fd_sc_hd__mux4_1
XFILLER_4_218 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_7 E6END[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2120_ net15 VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__buf_1
X_2051_ net797 net701 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1002_ Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 _0124_ _0126_ Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0
+ _0145_ VGND VGND VPWR VPWR _0146_ sky130_fd_sc_hd__o221a_1
X_1835_ net780 net673 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame8_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1904_ net768 net679 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame6_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0717_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit17.Q VGND VGND VPWR VPWR _0568_ sky130_fd_sc_hd__inv_1
X_1766_ net791 net740 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame10_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1697_ net802 net730 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame12_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2249_ NN4END[10] VGND VGND VPWR VPWR net288 sky130_fd_sc_hd__buf_1
X_2318_ Inst_LUT4AB_switch_matrix.JW2BEG2 VGND VGND VPWR VPWR net351 sky130_fd_sc_hd__buf_6
Xinput111 SS4END[2] VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__buf_2
Xinput100 S2MID[3] VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__buf_2
XFILLER_48_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput133 W6END[0] VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__clkbuf_4
Xinput122 W2END[5] VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__clkbuf_2
XFILLER_63_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1620_ net789 net723 VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4
+ sky130_fd_sc_hd__dlxtp_1
X_1482_ net481 Inst_LUT4AB_ConfigMem.Inst_frame9_bit30.Q net467 _0547_ VGND VGND VPWR
+ VPWR _0007_ sky130_fd_sc_hd__a31o_1
X_1551_ net44 net710 VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_8_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2103_ clknet_1_0__leaf_UserCLK_regs _0004_ VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.LUT_flop
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_37_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_45_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2034_ net761 net695 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1818_ net751 net671 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame8_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_10_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout801 net802 VGND VGND VPWR VPWR net801 sky130_fd_sc_hd__clkbuf_4
Xfanout812 net28 VGND VGND VPWR VPWR net812 sky130_fd_sc_hd__buf_4
X_1749_ net766 net739 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame10_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_13_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_39_Left_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_59_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_48_Left_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_57_Left_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0982_ Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 _0122_ _0125_ Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12
+ VGND VGND VPWR VPWR _0127_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_42_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1603_ net798 net718 VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6
+ sky130_fd_sc_hd__dlxtp_1
X_1534_ net807 net708 VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13
+ sky130_fd_sc_hd__dlxtp_1
X_1465_ net486 Inst_LUT4AB_ConfigMem.Inst_frame10_bit22.Q net467 _0533_ _0534_ VGND
+ VGND VPWR VPWR _0003_ sky130_fd_sc_hd__a32o_1
XPHY_EDGE_ROW_66_Left_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1396_ net653 _0120_ net664 _0044_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit8.Q Inst_LUT4AB_ConfigMem.Inst_frame13_bit9.Q
+ VGND VGND VPWR VPWR _0497_ sky130_fd_sc_hd__mux4_1
X_2017_ net802 net697 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
Xfanout642 net643 VGND VGND VPWR VPWR net642 sky130_fd_sc_hd__buf_8
Xfanout631 net633 VGND VGND VPWR VPWR net631 sky130_fd_sc_hd__buf_2
Xfanout697 net698 VGND VGND VPWR VPWR net697 sky130_fd_sc_hd__buf_2
Xfanout653 C VGND VGND VPWR VPWR net653 sky130_fd_sc_hd__buf_2
Xfanout675 net678 VGND VGND VPWR VPWR net675 sky130_fd_sc_hd__buf_2
Xfanout686 FrameStrobe[5] VGND VGND VPWR VPWR net686 sky130_fd_sc_hd__clkbuf_2
Xfanout664 _0265_ VGND VGND VPWR VPWR net664 sky130_fd_sc_hd__clkbuf_4
XFILLER_53_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1181_ Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 _0307_ _0308_ Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3
+ VGND VGND VPWR VPWR _0313_ sky130_fd_sc_hd__o22a_1
XFILLER_64_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1250_ net85 net87 net89 net113 Inst_LUT4AB_ConfigMem.Inst_frame1_bit22.Q Inst_LUT4AB_ConfigMem.Inst_frame1_bit23.Q
+ VGND VGND VPWR VPWR _0376_ sky130_fd_sc_hd__mux4_1
XFILLER_32_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput223 net223 VGND VGND VPWR VPWR FrameStrobe_O[12] sky130_fd_sc_hd__buf_2
Xoutput234 net234 VGND VGND VPWR VPWR FrameStrobe_O[4] sky130_fd_sc_hd__buf_2
Xoutput212 net212 VGND VGND VPWR VPWR FrameData_O[31] sky130_fd_sc_hd__buf_2
Xoutput201 net201 VGND VGND VPWR VPWR FrameData_O[21] sky130_fd_sc_hd__buf_2
X_0896_ net641 net632 H Inst_LUT4AB_switch_matrix.M_EF Inst_LUT4AB_ConfigMem.Inst_frame3_bit10.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame3_bit11.Q VGND VGND VPWR VPWR _0047_ sky130_fd_sc_hd__mux4_1
X_0965_ net64 net92 net9 net136 Inst_LUT4AB_ConfigMem.Inst_frame5_bit13.Q Inst_LUT4AB_ConfigMem.Inst_frame5_bit12.Q
+ VGND VGND VPWR VPWR _0111_ sky130_fd_sc_hd__mux4_2
Xoutput278 net278 VGND VGND VPWR VPWR NN4BEG[11] sky130_fd_sc_hd__buf_2
Xoutput245 net245 VGND VGND VPWR VPWR N2BEG[1] sky130_fd_sc_hd__buf_8
Xoutput289 net289 VGND VGND VPWR VPWR NN4BEG[7] sky130_fd_sc_hd__buf_2
Xoutput256 net256 VGND VGND VPWR VPWR N2BEGb[4] sky130_fd_sc_hd__buf_2
Xoutput267 net267 VGND VGND VPWR VPWR N4BEG[1] sky130_fd_sc_hd__buf_2
X_1517_ net774 net703 VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15
+ sky130_fd_sc_hd__dlxtp_1
X_1448_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit27.Q _0517_ _0520_ VGND VGND VPWR VPWR
+ _0521_ sky130_fd_sc_hd__a21o_1
XFILLER_70_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1379_ net647 net431 _0252_ _0640_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit31.Q Inst_LUT4AB_ConfigMem.Inst_frame12_bit0.Q
+ VGND VGND VPWR VPWR _0485_ sky130_fd_sc_hd__mux4_1
XFILLER_23_264 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_24_Left_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0750_ _0555_ _0600_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit1.Q VGND VGND VPWR VPWR
+ _0601_ sky130_fd_sc_hd__o21a_1
X_2282_ S4END[7] VGND VGND VPWR VPWR net321 sky130_fd_sc_hd__clkbuf_2
X_1233_ net85 net87 net109 net135 Inst_LUT4AB_ConfigMem.Inst_frame3_bit22.Q Inst_LUT4AB_ConfigMem.Inst_frame3_bit23.Q
+ VGND VGND VPWR VPWR _0361_ sky130_fd_sc_hd__mux4_1
X_2351_ WW4END[11] VGND VGND VPWR VPWR net390 sky130_fd_sc_hd__clkbuf_2
X_1302_ _0593_ _0420_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit29.Q VGND VGND VPWR VPWR
+ _0421_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_67_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1095_ _0231_ _0230_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit20.Q VGND VGND VPWR VPWR
+ _0232_ sky130_fd_sc_hd__mux2_4
X_1164_ _0581_ _0237_ _0295_ VGND VGND VPWR VPWR _0296_ sky130_fd_sc_hd__a21oi_1
X_0948_ net68 net96 net26 net124 Inst_LUT4AB_ConfigMem.Inst_frame5_bit11.Q Inst_LUT4AB_ConfigMem.Inst_frame5_bit10.Q
+ VGND VGND VPWR VPWR _0095_ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_50_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1997_ net776 net691 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_7_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0879_ Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 _0018_ _0022_ Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7
+ VGND VGND VPWR VPWR _0032_ sky130_fd_sc_hd__o22a_1
XFILLER_11_201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_64_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_72_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1920_ net803 net685 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame5_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1851_ net750 net675 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame7_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_12_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0802_ net65 net816 net10 net814 Inst_LUT4AB_ConfigMem.Inst_frame2_bit6.Q Inst_LUT4AB_ConfigMem.Inst_frame2_bit7.Q
+ VGND VGND VPWR VPWR _0649_ sky130_fd_sc_hd__mux4_1
X_0733_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit25.Q VGND VGND VPWR VPWR _0584_ sky130_fd_sc_hd__inv_1
X_1782_ net759 net670 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_69_267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2196_ net669 VGND VGND VPWR VPWR net239 sky130_fd_sc_hd__buf_1
X_2334_ W6END[4] VGND VGND VPWR VPWR net369 sky130_fd_sc_hd__clkbuf_2
X_1216_ Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 _0074_ _0334_ Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2
+ VGND VGND VPWR VPWR _0346_ sky130_fd_sc_hd__o22a_1
X_2265_ Inst_LUT4AB_switch_matrix.JS2BEG2 VGND VGND VPWR VPWR net298 sky130_fd_sc_hd__clkbuf_2
X_1078_ Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 _0212_ _0214_ Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3
+ VGND VGND VPWR VPWR _0216_ sky130_fd_sc_hd__a22o_1
XFILLER_40_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1147_ net69 net14 net125 Inst_LUT4AB_switch_matrix.JW2BEG6 Inst_LUT4AB_ConfigMem.Inst_frame7_bit24.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame7_bit25.Q VGND VGND VPWR VPWR _0280_ sky130_fd_sc_hd__mux4_2
XFILLER_25_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold88 Inst_LA_LUT4c_frame_config_dffesr.LUT_flop VGND VGND VPWR VPWR net480 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_43_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_26_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_8 E6END[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2050_ net800 net701 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1001_ Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 _0122_ _0125_ Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4
+ VGND VGND VPWR VPWR _0145_ sky130_fd_sc_hd__o22a_1
XFILLER_34_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1834_ net781 net673 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame8_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_32_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1903_ net770 net679 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame6_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1765_ net793 net741 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame10_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0716_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit13.Q VGND VGND VPWR VPWR _0567_ sky130_fd_sc_hd__inv_1
X_1696_ net804 net730 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame12_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2248_ NN4END[9] VGND VGND VPWR VPWR net287 sky130_fd_sc_hd__buf_1
X_2179_ net779 VGND VGND VPWR VPWR net204 sky130_fd_sc_hd__clkbuf_1
XFILLER_65_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2317_ Inst_LUT4AB_switch_matrix.JW2BEG1 VGND VGND VPWR VPWR net350 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_11_Left_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput112 SS4END[3] VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput101 S2MID[4] VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__clkbuf_2
Xinput134 W6END[1] VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput123 W2END[6] VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__clkbuf_2
XFILLER_71_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1481_ _0285_ _0292_ _0545_ _0546_ VGND VGND VPWR VPWR _0547_ sky130_fd_sc_hd__o31a_1
X_1550_ net772 net710 VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_47_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_37_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2102_ clknet_1_0__leaf_UserCLK_regs _0003_ VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.LUT_flop
+ sky130_fd_sc_hd__dfxtp_1
X_2033_ net763 net695 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1748_ net790 net54 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame10_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_30_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1817_ net753 net674 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame8_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1679_ net769 net729 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame13_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
Xfanout802 net33 VGND VGND VPWR VPWR net802 sky130_fd_sc_hd__buf_4
Xfanout813 net23 VGND VGND VPWR VPWR net813 sky130_fd_sc_hd__buf_2
XFILLER_53_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_59_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0981_ _0109_ _0121_ VGND VGND VPWR VPWR _0126_ sky130_fd_sc_hd__or2_4
XFILLER_44_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1602_ net799 net719 VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_8_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1395_ _0495_ _0496_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit13.Q VGND VGND VPWR VPWR
+ Inst_LUT4AB_switch_matrix.NN4BEG3 sky130_fd_sc_hd__mux2_4
X_1464_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit22.Q net621 _0532_ Inst_LC_LUT4c_frame_config_dffesr.c_reset_value
+ VGND VGND VPWR VPWR _0534_ sky130_fd_sc_hd__o2bb2a_1
X_1533_ net809 net707 VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12
+ sky130_fd_sc_hd__dlxtp_1
X_2016_ net803 net697 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_50_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout632 net633 VGND VGND VPWR VPWR net632 sky130_fd_sc_hd__buf_8
XFILLER_58_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout643 F VGND VGND VPWR VPWR net643 sky130_fd_sc_hd__buf_8
Xfanout665 net116 VGND VGND VPWR VPWR net665 sky130_fd_sc_hd__clkbuf_4
Xfanout698 FrameStrobe[2] VGND VGND VPWR VPWR net698 sky130_fd_sc_hd__clkbuf_2
Xfanout676 net677 VGND VGND VPWR VPWR net676 sky130_fd_sc_hd__clkbuf_2
Xfanout621 _0513_ VGND VGND VPWR VPWR net621 sky130_fd_sc_hd__buf_6
Xfanout654 net655 VGND VGND VPWR VPWR net654 sky130_fd_sc_hd__buf_8
Xfanout687 net56 VGND VGND VPWR VPWR net687 sky130_fd_sc_hd__buf_2
XFILLER_73_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1180_ Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 _0303_ _0304_ Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1
+ VGND VGND VPWR VPWR _0312_ sky130_fd_sc_hd__o22a_1
X_0964_ net83 net107 net8 Inst_LUT4AB_switch_matrix.E2BEG3 Inst_LUT4AB_ConfigMem.Inst_frame0_bit13.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame0_bit12.Q VGND VGND VPWR VPWR _0110_ sky130_fd_sc_hd__mux4_2
Xoutput224 net224 VGND VGND VPWR VPWR FrameStrobe_O[13] sky130_fd_sc_hd__buf_2
Xoutput235 net235 VGND VGND VPWR VPWR FrameStrobe_O[5] sky130_fd_sc_hd__buf_2
Xoutput246 net246 VGND VGND VPWR VPWR N2BEG[2] sky130_fd_sc_hd__buf_8
Xoutput257 net257 VGND VGND VPWR VPWR N2BEGb[5] sky130_fd_sc_hd__buf_2
Xoutput268 net268 VGND VGND VPWR VPWR N4BEG[2] sky130_fd_sc_hd__buf_2
Xoutput202 net202 VGND VGND VPWR VPWR FrameData_O[22] sky130_fd_sc_hd__buf_2
X_0895_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit12.Q _0045_ VGND VGND VPWR VPWR _0046_
+ sky130_fd_sc_hd__and2b_1
Xoutput213 net213 VGND VGND VPWR VPWR FrameData_O[3] sky130_fd_sc_hd__buf_2
X_1516_ net777 net703 VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14
+ sky130_fd_sc_hd__dlxtp_1
Xoutput279 net279 VGND VGND VPWR VPWR NN4BEG[12] sky130_fd_sc_hd__buf_4
X_1378_ net58 net3 net86 net638 Inst_LUT4AB_ConfigMem.Inst_frame13_bit31.Q Inst_LUT4AB_ConfigMem.Inst_frame12_bit0.Q
+ VGND VGND VPWR VPWR _0484_ sky130_fd_sc_hd__mux4_1
X_1447_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit27.Q _0519_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit28.Q
+ VGND VGND VPWR VPWR _0520_ sky130_fd_sc_hd__o21ai_1
XFILLER_23_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_298 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2281_ S4END[6] VGND VGND VPWR VPWR net320 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_67_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1232_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit24.Q _0359_ VGND VGND VPWR VPWR _0360_
+ sky130_fd_sc_hd__nand2b_1
X_2350_ WW4END[10] VGND VGND VPWR VPWR net389 sky130_fd_sc_hd__clkbuf_2
X_1301_ net639 net630 net625 net623 Inst_LUT4AB_ConfigMem.Inst_frame5_bit26.Q Inst_LUT4AB_ConfigMem.Inst_frame5_bit27.Q
+ VGND VGND VPWR VPWR _0420_ sky130_fd_sc_hd__mux4_1
X_1094_ net660 net656 net652 net636 Inst_LUT4AB_ConfigMem.Inst_frame4_bit18.Q Inst_LUT4AB_ConfigMem.Inst_frame4_bit19.Q
+ VGND VGND VPWR VPWR _0231_ sky130_fd_sc_hd__mux4_1
X_1163_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit9.Q _0238_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit10.Q
+ VGND VGND VPWR VPWR _0295_ sky130_fd_sc_hd__a21o_1
XFILLER_52_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_50_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1996_ net43 net693 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_60_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0947_ net80 net120 net9 Inst_LUT4AB_switch_matrix.JN2BEG3 Inst_LUT4AB_ConfigMem.Inst_frame0_bit11.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame0_bit10.Q VGND VGND VPWR VPWR _0094_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_15_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0878_ Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 _0019_ _0015_ VGND
+ VGND VPWR VPWR _0031_ sky130_fd_sc_hd__o21ba_1
XFILLER_55_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_72_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_29_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1781_ net765 net670 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1850_ net752 net677 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame7_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_12_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0801_ _0557_ _0647_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit9.Q VGND VGND VPWR VPWR
+ _0648_ sky130_fd_sc_hd__o21a_1
X_0732_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit25.Q VGND VGND VPWR VPWR _0583_ sky130_fd_sc_hd__inv_1
X_2333_ W6END[3] VGND VGND VPWR VPWR net368 sky130_fd_sc_hd__clkbuf_2
X_1146_ _0275_ _0576_ _0278_ _0279_ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.JW2BEG6
+ sky130_fd_sc_hd__o22a_4
XFILLER_69_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2195_ net671 VGND VGND VPWR VPWR net238 sky130_fd_sc_hd__clkbuf_1
X_1215_ Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 _0075_ _0336_ Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4
+ VGND VGND VPWR VPWR _0345_ sky130_fd_sc_hd__o22a_1
X_2264_ Inst_LUT4AB_switch_matrix.JS2BEG1 VGND VGND VPWR VPWR net297 sky130_fd_sc_hd__clkbuf_2
X_1077_ Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 _0210_ _0213_ Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5
+ VGND VGND VPWR VPWR _0215_ sky130_fd_sc_hd__a22o_1
X_1979_ net750 net691 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_29_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold89 Inst_LG_LUT4c_frame_config_dffesr.LUT_flop VGND VGND VPWR VPWR net481 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_16_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_9 E6END[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1000_ _0128_ _0143_ _0097_ VGND VGND VPWR VPWR _0144_ sky130_fd_sc_hd__mux2_4
XFILLER_3_297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1902_ net772 net682 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame6_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_19_187 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1833_ net783 net673 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame8_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0715_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit13.Q VGND VGND VPWR VPWR _0566_ sky130_fd_sc_hd__inv_1
X_1764_ net796 net741 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame10_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2316_ Inst_LUT4AB_switch_matrix.JW2BEG0 VGND VGND VPWR VPWR net349 sky130_fd_sc_hd__clkbuf_1
X_1695_ net806 net730 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame12_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2247_ NN4END[8] VGND VGND VPWR VPWR net286 sky130_fd_sc_hd__buf_1
X_1129_ _0574_ _0259_ _0263_ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.E2BEG6
+ sky130_fd_sc_hd__o21a_4
X_2178_ net782 VGND VGND VPWR VPWR net203 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_48_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput102 S2MID[5] VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput113 W1END[0] VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__buf_4
Xinput124 W2END[7] VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__clkbuf_2
Xinput135 WW4END[0] VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__buf_2
XFILLER_72_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1480_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit30.Q net621 _0544_ Inst_LG_LUT4c_frame_config_dffesr.c_reset_value
+ VGND VGND VPWR VPWR _0546_ sky130_fd_sc_hd__o2bb2a_1
XPHY_EDGE_ROW_28_Right_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_37_Right_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_37_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2032_ net768 net695 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2101_ clknet_1_0__leaf_UserCLK_regs _0002_ VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.LUT_flop
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_45_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1678_ net772 net727 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame13_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_46_Right_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1747_ net812 net54 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame10_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1816_ net755 net674 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame8_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
Xfanout803 net804 VGND VGND VPWR VPWR net803 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_55_Right_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout814 net22 VGND VGND VPWR VPWR net814 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_64_Right_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_73_Right_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0980_ _0121_ _0109_ VGND VGND VPWR VPWR _0125_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_42_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1601_ net801 net718 VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4
+ sky130_fd_sc_hd__dlxtp_1
X_1532_ net747 net708 VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_8_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1394_ net647 net431 _0252_ _0606_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit11.Q Inst_LUT4AB_ConfigMem.Inst_frame13_bit12.Q
+ VGND VGND VPWR VPWR _0496_ sky130_fd_sc_hd__mux4_2
X_1463_ _0203_ _0532_ VGND VGND VPWR VPWR _0533_ sky130_fd_sc_hd__nand2b_1
XFILLER_4_392 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2015_ net805 net697 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_35_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout622 Inst_LUT4AB_switch_matrix.M_EF VGND VGND VPWR VPWR net622 sky130_fd_sc_hd__buf_12
Xfanout633 G VGND VGND VPWR VPWR net633 sky130_fd_sc_hd__buf_8
XFILLER_5_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout688 net690 VGND VGND VPWR VPWR net688 sky130_fd_sc_hd__clkbuf_2
XFILLER_58_344 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout666 net115 VGND VGND VPWR VPWR net666 sky130_fd_sc_hd__clkbuf_4
Xfanout677 net678 VGND VGND VPWR VPWR net677 sky130_fd_sc_hd__buf_2
Xfanout699 FrameStrobe[1] VGND VGND VPWR VPWR net699 sky130_fd_sc_hd__buf_2
Xfanout644 net645 VGND VGND VPWR VPWR net644 sky130_fd_sc_hd__buf_4
Xfanout655 B VGND VGND VPWR VPWR net655 sky130_fd_sc_hd__buf_8
XFILLER_53_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0894_ net661 net656 C net637 Inst_LUT4AB_ConfigMem.Inst_frame3_bit10.Q Inst_LUT4AB_ConfigMem.Inst_frame3_bit11.Q
+ VGND VGND VPWR VPWR _0045_ sky130_fd_sc_hd__mux4_2
X_0963_ net431 _0108_ _0099_ _0098_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit15.Q Inst_LUT4AB_ConfigMem.Inst_frame9_bit16.Q
+ VGND VGND VPWR VPWR _0109_ sky130_fd_sc_hd__mux4_2
XFILLER_32_288 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput225 net225 VGND VGND VPWR VPWR FrameStrobe_O[14] sky130_fd_sc_hd__buf_2
Xoutput236 net236 VGND VGND VPWR VPWR FrameStrobe_O[6] sky130_fd_sc_hd__buf_2
Xoutput247 net247 VGND VGND VPWR VPWR N2BEG[3] sky130_fd_sc_hd__buf_6
Xoutput269 net269 VGND VGND VPWR VPWR N4BEG[3] sky130_fd_sc_hd__buf_2
Xoutput258 net258 VGND VGND VPWR VPWR N2BEGb[6] sky130_fd_sc_hd__buf_2
Xoutput203 net203 VGND VGND VPWR VPWR FrameData_O[23] sky130_fd_sc_hd__buf_2
Xoutput214 net214 VGND VGND VPWR VPWR FrameData_O[4] sky130_fd_sc_hd__buf_2
X_1515_ net779 net703 VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13
+ sky130_fd_sc_hd__dlxtp_1
X_1377_ _0480_ _0483_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit5.Q VGND VGND VPWR VPWR
+ Inst_LUT4AB_switch_matrix.E6BEG0 sky130_fd_sc_hd__mux2_4
X_1446_ _0518_ VGND VGND VPWR VPWR _0519_ sky130_fd_sc_hd__inv_1
XFILLER_63_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2280_ S4END[5] VGND VGND VPWR VPWR net319 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_67_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1231_ net57 net61 net2 net6 Inst_LUT4AB_ConfigMem.Inst_frame3_bit22.Q Inst_LUT4AB_ConfigMem.Inst_frame3_bit23.Q
+ VGND VGND VPWR VPWR _0359_ sky130_fd_sc_hd__mux4_1
XFILLER_64_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1162_ _0211_ _0204_ _0126_ _0212_ _0269_ VGND VGND VPWR VPWR _0294_ sky130_fd_sc_hd__a311o_1
X_1300_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit28.Q _0418_ VGND VGND VPWR VPWR _0419_
+ sky130_fd_sc_hd__or2_1
X_1093_ net646 net627 net641 Inst_LUT4AB_switch_matrix.M_AH Inst_LUT4AB_ConfigMem.Inst_frame4_bit19.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame4_bit18.Q VGND VGND VPWR VPWR _0230_ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_50_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1995_ net42 net693 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0946_ net76 net21 net104 net132 Inst_LUT4AB_ConfigMem.Inst_frame6_bit10.Q Inst_LUT4AB_ConfigMem.Inst_frame6_bit11.Q
+ VGND VGND VPWR VPWR _0093_ sky130_fd_sc_hd__mux4_2
X_0877_ Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 _0018_ _0029_ _0015_
+ VGND VGND VPWR VPWR _0030_ sky130_fd_sc_hd__o211a_1
XFILLER_20_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_7_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1429_ net644 Inst_LUT4AB_switch_matrix.JW2BEG1 net664 _0271_ Inst_LUT4AB_ConfigMem.Inst_frame14_bit23.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame14_bit22.Q VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.N1BEG2
+ sky130_fd_sc_hd__mux4_1
XFILLER_11_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_29_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0731_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit25.Q VGND VGND VPWR VPWR _0582_ sky130_fd_sc_hd__inv_1
X_1780_ net789 net670 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_12_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0800_ net640 net630 net624 net397 Inst_LUT4AB_ConfigMem.Inst_frame2_bit6.Q Inst_LUT4AB_ConfigMem.Inst_frame2_bit7.Q
+ VGND VGND VPWR VPWR _0647_ sky130_fd_sc_hd__mux4_2
XFILLER_69_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2332_ W6END[2] VGND VGND VPWR VPWR net365 sky130_fd_sc_hd__clkbuf_2
X_1145_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit20.Q _0276_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit21.Q
+ VGND VGND VPWR VPWR _0279_ sky130_fd_sc_hd__a21o_1
X_2194_ net676 VGND VGND VPWR VPWR net237 sky130_fd_sc_hd__buf_1
X_1214_ _0342_ _0343_ VGND VGND VPWR VPWR _0344_ sky130_fd_sc_hd__nand2_1
X_2263_ Inst_LUT4AB_switch_matrix.JS2BEG0 VGND VGND VPWR VPWR net296 sky130_fd_sc_hd__buf_6
XFILLER_52_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1076_ _0208_ _0209_ VGND VGND VPWR VPWR _0214_ sky130_fd_sc_hd__and2b_1
XFILLER_18_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0929_ _0052_ _0053_ _0044_ _0043_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit25.Q Inst_LUT4AB_ConfigMem.Inst_frame10_bit26.Q
+ VGND VGND VPWR VPWR _0077_ sky130_fd_sc_hd__mux4_2
X_1978_ net752 net691 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_29_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1832_ net786 net673 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame8_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1901_ net774 net682 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame6_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_22_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0714_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit5.Q VGND VGND VPWR VPWR _0565_ sky130_fd_sc_hd__inv_1
X_1763_ net798 net741 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame10_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1694_ net808 net732 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame12_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2246_ NN4END[7] VGND VGND VPWR VPWR net285 sky130_fd_sc_hd__clkbuf_1
X_1128_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit20.Q _0260_ _0262_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit21.Q
+ VGND VGND VPWR VPWR _0263_ sky130_fd_sc_hd__a211o_1
XFILLER_65_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2177_ net784 VGND VGND VPWR VPWR net202 sky130_fd_sc_hd__clkbuf_2
XFILLER_25_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1059_ Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 _0079_ _0171_ Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5
+ VGND VGND VPWR VPWR _0198_ sky130_fd_sc_hd__a22o_1
XFILLER_40_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput103 S2MID[6] VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput125 W2MID[0] VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__clkbuf_2
Xinput114 W1END[1] VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__clkbuf_4
Xinput136 WW4END[1] VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__clkbuf_2
XFILLER_71_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2100_ clknet_1_0__leaf_UserCLK_regs _0001_ VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.LUT_flop
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_62_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_37_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2031_ net770 net695 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1815_ net758 net672 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame8_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_45_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout815 net5 VGND VGND VPWR VPWR net815 sky130_fd_sc_hd__clkbuf_4
Xfanout804 net32 VGND VGND VPWR VPWR net804 sky130_fd_sc_hd__buf_4
X_1677_ net775 net726 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame13_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1746_ net47 net735 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame11_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_7_82 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2229_ N4END[6] VGND VGND VPWR VPWR net268 sky130_fd_sc_hd__clkbuf_1
XFILLER_53_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_42_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1600_ net32 net719 VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_26_Left_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1462_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit31.Q _0522_ VGND VGND VPWR VPWR _0532_
+ sky130_fd_sc_hd__nand2_1
X_1531_ net749 net707 VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10
+ sky130_fd_sc_hd__dlxtp_1
X_1393_ net58 net3 net114 net638 Inst_LUT4AB_ConfigMem.Inst_frame13_bit11.Q Inst_LUT4AB_ConfigMem.Inst_frame13_bit12.Q
+ VGND VGND VPWR VPWR _0495_ sky130_fd_sc_hd__mux4_1
XFILLER_27_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2014_ net808 net698 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_35_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout656 net657 VGND VGND VPWR VPWR net656 sky130_fd_sc_hd__buf_2
X_1729_ net802 net737 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame11_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
Xfanout623 Inst_LUT4AB_switch_matrix.M_AB VGND VGND VPWR VPWR net623 sky130_fd_sc_hd__buf_6
Xfanout667 net668 VGND VGND VPWR VPWR net667 sky130_fd_sc_hd__clkbuf_2
Xfanout645 net648 VGND VGND VPWR VPWR net645 sky130_fd_sc_hd__buf_2
Xfanout634 D VGND VGND VPWR VPWR net634 sky130_fd_sc_hd__buf_8
XFILLER_73_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout689 net690 VGND VGND VPWR VPWR net689 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_58_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout678 FrameStrobe[7] VGND VGND VPWR VPWR net678 sky130_fd_sc_hd__clkbuf_2
XFILLER_37_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_286 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_323 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_264 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0962_ net74 net19 net102 net130 Inst_LUT4AB_ConfigMem.Inst_frame6_bit14.Q Inst_LUT4AB_ConfigMem.Inst_frame6_bit15.Q
+ VGND VGND VPWR VPWR _0108_ sky130_fd_sc_hd__mux4_1
X_0893_ net63 net8 net91 net137 Inst_LUT4AB_ConfigMem.Inst_frame5_bit4.Q Inst_LUT4AB_ConfigMem.Inst_frame5_bit5.Q
+ VGND VGND VPWR VPWR _0044_ sky130_fd_sc_hd__mux4_2
Xoutput226 net226 VGND VGND VPWR VPWR FrameStrobe_O[15] sky130_fd_sc_hd__buf_2
Xoutput237 net237 VGND VGND VPWR VPWR FrameStrobe_O[7] sky130_fd_sc_hd__buf_2
Xoutput248 net248 VGND VGND VPWR VPWR N2BEG[4] sky130_fd_sc_hd__buf_6
Xoutput204 net204 VGND VGND VPWR VPWR FrameData_O[24] sky130_fd_sc_hd__buf_2
Xoutput259 net259 VGND VGND VPWR VPWR N2BEGb[7] sky130_fd_sc_hd__buf_2
Xoutput215 net215 VGND VGND VPWR VPWR FrameData_O[5] sky130_fd_sc_hd__buf_2
X_1445_ Inst_LUT4AB_switch_matrix.JN2BEG1 Inst_LUT4AB_switch_matrix.E2BEG1 Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q
+ VGND VGND VPWR VPWR _0518_ sky130_fd_sc_hd__mux2_1
X_1514_ net782 net705 VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12
+ sky130_fd_sc_hd__dlxtp_1
X_1376_ _0482_ _0481_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit4.Q VGND VGND VPWR VPWR
+ _0483_ sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_61_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_120 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1230_ _0356_ _0357_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit24.Q VGND VGND VPWR VPWR
+ _0358_ sky130_fd_sc_hd__mux2_4
XFILLER_64_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1161_ _0292_ _0285_ Inst_LG_LUT4c_frame_config_dffesr.c_out_mux _0293_ VGND VGND
+ VPWR VPWR G sky130_fd_sc_hd__o31a_4
X_1092_ _0126_ _0204_ _0211_ _0212_ VGND VGND VPWR VPWR _0229_ sky130_fd_sc_hd__a31o_1
XFILLER_49_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1994_ net781 net693 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_50_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0945_ net75 net131 net20 Inst_LUT4AB_switch_matrix.JN2BEG5 Inst_LUT4AB_ConfigMem.Inst_frame7_bit11.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame7_bit10.Q VGND VGND VPWR VPWR _0092_ sky130_fd_sc_hd__mux4_1
XFILLER_9_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0876_ Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 _0022_ _0023_ Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9
+ _0028_ VGND VGND VPWR VPWR _0029_ sky130_fd_sc_hd__o221a_1
X_1428_ net643 _0653_ Inst_LUT4AB_switch_matrix.JW2BEG2 _0639_ Inst_LUT4AB_ConfigMem.Inst_frame14_bit24.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame14_bit25.Q VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.N1BEG3
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_7_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1359_ _0652_ _0071_ net431 _0252_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit6.Q Inst_LUT4AB_ConfigMem.Inst_frame12_bit7.Q
+ VGND VGND VPWR VPWR _0467_ sky130_fd_sc_hd__mux4_2
XFILLER_55_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0730_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit9.Q VGND VGND VPWR VPWR _0581_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_12_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1213_ Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 _0074_ _0336_ Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5
+ VGND VGND VPWR VPWR _0343_ sky130_fd_sc_hd__o22a_1
X_2331_ net132 VGND VGND VPWR VPWR net364 sky130_fd_sc_hd__clkbuf_2
X_1144_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit20.Q _0277_ VGND VGND VPWR VPWR _0278_
+ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_63_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1075_ _0209_ _0208_ VGND VGND VPWR VPWR _0213_ sky130_fd_sc_hd__and2b_1
X_2193_ net681 VGND VGND VPWR VPWR net236 sky130_fd_sc_hd__buf_1
X_1977_ net754 net691 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0928_ _0075_ VGND VGND VPWR VPWR _0076_ sky130_fd_sc_hd__inv_2
XFILLER_0_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0859_ net1 _0663_ _0608_ _0619_ VGND VGND VPWR VPWR _0012_ sky130_fd_sc_hd__a211o_1
XFILLER_45_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1831_ net788 net673 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame8_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_42_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1900_ net777 net680 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame6_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0713_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit5.Q VGND VGND VPWR VPWR _0564_ sky130_fd_sc_hd__inv_1
X_1762_ net799 net740 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame10_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1693_ net810 net732 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame12_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2245_ NN4END[6] VGND VGND VPWR VPWR net284 sky130_fd_sc_hd__clkbuf_1
XFILLER_57_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2176_ net785 VGND VGND VPWR VPWR net201 sky130_fd_sc_hd__buf_1
X_1127_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit20.Q _0261_ VGND VGND VPWR VPWR _0262_
+ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_48_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1058_ _0196_ _0174_ _0170_ VGND VGND VPWR VPWR _0197_ sky130_fd_sc_hd__mux2_4
XFILLER_25_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_23_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput104 S2MID[7] VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput115 W1END[2] VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__buf_2
Xinput126 W2MID[1] VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_56_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput137 WW4END[2] VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__buf_2
XFILLER_71_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2030_ net773 net695 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_62_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1814_ net760 net672 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame8_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1745_ net764 net735 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame11_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
Xfanout805 net806 VGND VGND VPWR VPWR net805 sky130_fd_sc_hd__clkbuf_4
X_1676_ net43 net726 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame13_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
Xfanout816 net4 VGND VGND VPWR VPWR net816 sky130_fd_sc_hd__clkbuf_4
XFILLER_7_94 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_15_Left_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2159_ net758 VGND VGND VPWR VPWR net214 sky130_fd_sc_hd__clkbuf_1
X_2228_ N4END[5] VGND VGND VPWR VPWR net267 sky130_fd_sc_hd__clkbuf_1
XFILLER_38_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_251 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_70 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1392_ _0494_ _0493_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit24.Q VGND VGND VPWR VPWR
+ Inst_LUT4AB_switch_matrix.EE4BEG0 sky130_fd_sc_hd__mux2_1
X_1530_ net751 net707 VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9
+ sky130_fd_sc_hd__dlxtp_1
X_1461_ net487 Inst_LUT4AB_ConfigMem.Inst_frame10_bit12.Q net467 _0530_ _0531_ VGND
+ VGND VPWR VPWR _0002_ sky130_fd_sc_hd__a32o_1
XFILLER_67_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2013_ net810 net698 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1728_ net804 net738 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame11_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
Xfanout646 net647 VGND VGND VPWR VPWR net646 sky130_fd_sc_hd__buf_2
X_1659_ net750 net727 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame13_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
Xfanout668 net669 VGND VGND VPWR VPWR net668 sky130_fd_sc_hd__clkbuf_2
Xfanout657 net658 VGND VGND VPWR VPWR net657 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout635 D VGND VGND VPWR VPWR net635 sky130_fd_sc_hd__buf_2
Xfanout679 FrameStrobe[6] VGND VGND VPWR VPWR net679 sky130_fd_sc_hd__clkbuf_2
Xfanout624 net625 VGND VGND VPWR VPWR net624 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_56_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0961_ net73 net129 net101 net408 Inst_LUT4AB_ConfigMem.Inst_frame7_bit15.Q Inst_LUT4AB_ConfigMem.Inst_frame7_bit14.Q
+ VGND VGND VPWR VPWR _0107_ sky130_fd_sc_hd__mux4_2
XFILLER_17_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput205 net205 VGND VGND VPWR VPWR FrameData_O[25] sky130_fd_sc_hd__buf_2
Xoutput216 net216 VGND VGND VPWR VPWR FrameData_O[6] sky130_fd_sc_hd__buf_2
X_0892_ net79 net8 net124 Inst_LUT4AB_switch_matrix.E2BEG2 Inst_LUT4AB_ConfigMem.Inst_frame0_bit4.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame0_bit5.Q VGND VGND VPWR VPWR _0043_ sky130_fd_sc_hd__mux4_2
Xoutput249 Inst_LUT4AB_switch_matrix.JN2BEG5 VGND VGND VPWR VPWR N2BEG[5] sky130_fd_sc_hd__buf_6
Xoutput238 net238 VGND VGND VPWR VPWR FrameStrobe_O[8] sky130_fd_sc_hd__buf_2
Xoutput227 net227 VGND VGND VPWR VPWR FrameStrobe_O[16] sky130_fd_sc_hd__buf_2
X_1375_ net413 net628 net623 net427 Inst_LUT4AB_ConfigMem.Inst_frame12_bit2.Q Inst_LUT4AB_ConfigMem.Inst_frame12_bit3.Q
+ VGND VGND VPWR VPWR _0482_ sky130_fd_sc_hd__mux4_2
X_1513_ net784 net705 VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11
+ sky130_fd_sc_hd__dlxtp_1
X_1444_ Inst_LUT4AB_switch_matrix.JS2BEG1 Inst_LUT4AB_switch_matrix.JW2BEG1 Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q
+ VGND VGND VPWR VPWR _0517_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_53_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_45_Left_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_18_Left_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_54_Left_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_63_Left_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1160_ Inst_LG_LUT4c_frame_config_dffesr.LUT_flop Inst_LG_LUT4c_frame_config_dffesr.c_out_mux
+ VGND VGND VPWR VPWR _0293_ sky130_fd_sc_hd__nand2b_1
X_1091_ _0228_ Inst_LF_LUT4c_frame_config_dffesr.LUT_flop Inst_LF_LUT4c_frame_config_dffesr.c_out_mux
+ VGND VGND VPWR VPWR F sky130_fd_sc_hd__mux2_4
XFILLER_49_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_72_Left_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1993_ net783 net693 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0944_ _0087_ _0568_ _0089_ _0091_ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.JN2BEG5
+ sky130_fd_sc_hd__o22a_4
XTAP_TAPCELL_ROW_50_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_238 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0875_ Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 _0019_ VGND VGND
+ VPWR VPWR _0028_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_66_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1358_ _0596_ _0462_ _0466_ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.SS4BEG0
+ sky130_fd_sc_hd__o21a_1
X_1427_ net63 net78 net23 net645 Inst_LUT4AB_ConfigMem.Inst_frame14_bit26.Q Inst_LUT4AB_ConfigMem.Inst_frame14_bit27.Q
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.N4BEG0 sky130_fd_sc_hd__mux4_1
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1289_ _0408_ _0409_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit28.Q VGND VGND VPWR VPWR
+ _0410_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_3_Left_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2192_ net685 VGND VGND VPWR VPWR net235 sky130_fd_sc_hd__buf_1
X_2330_ net131 VGND VGND VPWR VPWR net363 sky130_fd_sc_hd__clkbuf_2
XFILLER_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1212_ Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 _0075_ _0334_ Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3
+ VGND VGND VPWR VPWR _0342_ sky130_fd_sc_hd__o22a_1
X_1143_ net60 net68 net815 net13 Inst_LUT4AB_ConfigMem.Inst_frame1_bit18.Q Inst_LUT4AB_ConfigMem.Inst_frame1_bit19.Q
+ VGND VGND VPWR VPWR _0277_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_63_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1074_ _0208_ _0209_ VGND VGND VPWR VPWR _0212_ sky130_fd_sc_hd__and2_1
X_1976_ net756 net693 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0927_ _0073_ _0054_ VGND VGND VPWR VPWR _0075_ sky130_fd_sc_hd__nand2_4
X_0789_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit0.Q _0636_ VGND VGND VPWR VPWR _0637_
+ sky130_fd_sc_hd__nand2b_1
X_0858_ _0663_ net1 VGND VGND VPWR VPWR _0011_ sky130_fd_sc_hd__or2_4
XFILLER_45_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_168 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1830_ net792 net673 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame8_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_30_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1761_ net801 net742 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame10_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0712_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit21.Q VGND VGND VPWR VPWR _0563_ sky130_fd_sc_hd__inv_1
X_1692_ net53 net733 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame12_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1126_ net60 net68 net815 net13 Inst_LUT4AB_ConfigMem.Inst_frame3_bit18.Q Inst_LUT4AB_ConfigMem.Inst_frame3_bit19.Q
+ VGND VGND VPWR VPWR _0261_ sky130_fd_sc_hd__mux4_1
X_2244_ NN4END[5] VGND VGND VPWR VPWR net283 sky130_fd_sc_hd__clkbuf_1
X_2175_ net787 VGND VGND VPWR VPWR net200 sky130_fd_sc_hd__clkbuf_1
XFILLER_57_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1057_ _0194_ _0195_ VGND VGND VPWR VPWR _0196_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_23_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1959_ net788 net689 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_31_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput105 S4END[0] VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__buf_2
Xinput116 W1END[3] VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__clkbuf_2
Xinput127 W2MID[2] VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__clkbuf_2
Xinput138 WW4END[3] VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_6_Left_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1813_ net765 net671 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame8_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1744_ net768 net735 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame11_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1675_ net779 net727 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame13_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
Xfanout806 net31 VGND VGND VPWR VPWR net806 sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2158_ net760 VGND VGND VPWR VPWR net213 sky130_fd_sc_hd__buf_1
X_1109_ net660 net657 net652 net636 Inst_LUT4AB_ConfigMem.Inst_frame2_bit18.Q Inst_LUT4AB_ConfigMem.Inst_frame2_bit19.Q
+ VGND VGND VPWR VPWR _0245_ sky130_fd_sc_hd__mux4_1
X_2227_ N4END[4] VGND VGND VPWR VPWR net260 sky130_fd_sc_hd__clkbuf_1
X_2089_ net783 net746 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame0_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_33_Right_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_318 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_42_Right_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_51_Right_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1391_ net59 net87 net816 net642 Inst_LUT4AB_ConfigMem.Inst_frame13_bit23.Q Inst_LUT4AB_ConfigMem.Inst_frame13_bit22.Q
+ VGND VGND VPWR VPWR _0494_ sky130_fd_sc_hd__mux4_1
X_1460_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit12.Q net621 _0529_ Inst_LB_LUT4c_frame_config_dffesr.c_reset_value
+ VGND VGND VPWR VPWR _0531_ sky130_fd_sc_hd__o2bb2a_1
XPHY_EDGE_ROW_60_Right_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2012_ net748 net695 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_50_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1658_ net752 net726 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame13_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1727_ net806 net738 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame11_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout636 net637 VGND VGND VPWR VPWR net636 sky130_fd_sc_hd__buf_2
X_1589_ net766 net717 VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11
+ sky130_fd_sc_hd__dlxtp_1
Xfanout669 net670 VGND VGND VPWR VPWR net669 sky130_fd_sc_hd__clkbuf_2
Xfanout647 net648 VGND VGND VPWR VPWR net647 sky130_fd_sc_hd__clkbuf_4
Xfanout658 B VGND VGND VPWR VPWR net658 sky130_fd_sc_hd__clkbuf_4
Xfanout625 net626 VGND VGND VPWR VPWR net625 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_56_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0960_ _0102_ _0570_ _0104_ _0106_ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.JS2BEG5
+ sky130_fd_sc_hd__o22a_1
Xoutput239 net239 VGND VGND VPWR VPWR FrameStrobe_O[9] sky130_fd_sc_hd__buf_2
Xoutput206 net206 VGND VGND VPWR VPWR FrameData_O[26] sky130_fd_sc_hd__buf_2
Xoutput228 net228 VGND VGND VPWR VPWR FrameStrobe_O[17] sky130_fd_sc_hd__buf_2
Xoutput217 net217 VGND VGND VPWR VPWR FrameData_O[7] sky130_fd_sc_hd__buf_2
X_0891_ _0565_ _0038_ _0040_ _0042_ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.E2BEG2
+ sky130_fd_sc_hd__o22a_4
X_1512_ net785 net705 VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10
+ sky130_fd_sc_hd__dlxtp_1
X_1374_ _0617_ _0053_ _0120_ net664 Inst_LUT4AB_ConfigMem.Inst_frame12_bit2.Q Inst_LUT4AB_ConfigMem.Inst_frame12_bit3.Q
+ VGND VGND VPWR VPWR _0481_ sky130_fd_sc_hd__mux4_1
XFILLER_4_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1443_ _0514_ _0515_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit27.Q VGND VGND VPWR VPWR
+ _0516_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_53_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_69_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_328 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1090_ _0222_ _0227_ _0218_ VGND VGND VPWR VPWR _0228_ sky130_fd_sc_hd__mux2_4
XFILLER_37_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1992_ net786 net693 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0943_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit16.Q _0090_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit17.Q
+ VGND VGND VPWR VPWR _0091_ sky130_fd_sc_hd__a21o_1
X_0874_ _0024_ _0026_ _0015_ VGND VGND VPWR VPWR _0027_ sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_15_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1426_ net64 net79 net22 net641 Inst_LUT4AB_ConfigMem.Inst_frame14_bit28.Q Inst_LUT4AB_ConfigMem.Inst_frame14_bit29.Q
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.N4BEG1 sky130_fd_sc_hd__mux4_2
X_1357_ _0463_ _0464_ _0465_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit27.Q Inst_LUT4AB_ConfigMem.Inst_frame12_bit28.Q
+ VGND VGND VPWR VPWR _0466_ sky130_fd_sc_hd__a221o_1
X_1288_ net90 net118 net106 net134 Inst_LUT4AB_ConfigMem.Inst_frame3_bit27.Q Inst_LUT4AB_ConfigMem.Inst_frame3_bit26.Q
+ VGND VGND VPWR VPWR _0409_ sky130_fd_sc_hd__mux4_1
XFILLER_34_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1142_ net86 net88 net96 net665 Inst_LUT4AB_ConfigMem.Inst_frame1_bit18.Q Inst_LUT4AB_ConfigMem.Inst_frame1_bit19.Q
+ VGND VGND VPWR VPWR _0276_ sky130_fd_sc_hd__mux4_1
X_2191_ net690 VGND VGND VPWR VPWR net234 sky130_fd_sc_hd__clkbuf_2
X_1211_ _0337_ _0340_ _0333_ VGND VGND VPWR VPWR _0341_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_63_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1073_ _0210_ VGND VGND VPWR VPWR _0211_ sky130_fd_sc_hd__inv_2
XFILLER_33_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1975_ net758 net693 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0926_ _0054_ _0073_ VGND VGND VPWR VPWR _0074_ sky130_fd_sc_hd__or2_4
X_0857_ _0009_ _0008_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit14.Q VGND VGND VPWR VPWR
+ _0010_ sky130_fd_sc_hd__mux2_2
XFILLER_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0788_ net63 net2 net79 net8 Inst_LUT4AB_ConfigMem.Inst_frame5_bit31.Q Inst_LUT4AB_ConfigMem.Inst_frame5_bit30.Q
+ VGND VGND VPWR VPWR _0636_ sky130_fd_sc_hd__mux4_1
X_1409_ net624 Inst_LUT4AB_switch_matrix.JS2BEG1 net664 _0271_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit11.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame11_bit10.Q VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.W1BEG2
+ sky130_fd_sc_hd__mux4_2
XFILLER_68_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1691_ net52 net733 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame12_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0711_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit1.Q VGND VGND VPWR VPWR _0562_ sky130_fd_sc_hd__inv_1
X_1760_ net804 net742 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame10_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2312_ Inst_LUT4AB_switch_matrix.W1BEG0 VGND VGND VPWR VPWR net345 sky130_fd_sc_hd__buf_1
X_2243_ NN4END[4] VGND VGND VPWR VPWR net276 sky130_fd_sc_hd__buf_1
X_1125_ net86 net88 net96 net665 Inst_LUT4AB_ConfigMem.Inst_frame3_bit18.Q Inst_LUT4AB_ConfigMem.Inst_frame3_bit19.Q
+ VGND VGND VPWR VPWR _0260_ sky130_fd_sc_hd__mux4_1
X_2174_ net791 VGND VGND VPWR VPWR net198 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_48_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1056_ Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 _0079_ _0171_ Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12
+ VGND VGND VPWR VPWR _0195_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_23_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_323 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_356 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1958_ net792 net688 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1889_ net33 net681 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame6_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0909_ net92 net120 net108 net134 Inst_LUT4AB_ConfigMem.Inst_frame2_bit3.Q Inst_LUT4AB_ConfigMem.Inst_frame2_bit2.Q
+ VGND VGND VPWR VPWR _0059_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_31_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput106 S4END[1] VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__buf_2
Xinput128 W2MID[3] VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__clkbuf_2
Xinput117 W2END[0] VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__clkbuf_2
XFILLER_71_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_90 net755 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1674_ net782 net727 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame13_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1812_ net789 net671 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame8_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1743_ net770 net735 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame11_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_30_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout807 net808 VGND VGND VPWR VPWR net807 sky130_fd_sc_hd__clkbuf_4
X_2226_ net76 VGND VGND VPWR VPWR net259 sky130_fd_sc_hd__clkbuf_2
XFILLER_53_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2088_ net786 net746 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame0_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1108_ net82 net94 net11 net122 Inst_LUT4AB_ConfigMem.Inst_frame5_bit23.Q Inst_LUT4AB_ConfigMem.Inst_frame5_bit22.Q
+ VGND VGND VPWR VPWR _0244_ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_36_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1039_ net58 net64 net27 net813 Inst_LUT4AB_ConfigMem.Inst_frame1_bit2.Q Inst_LUT4AB_ConfigMem.Inst_frame1_bit3.Q
+ VGND VGND VPWR VPWR _0180_ sky130_fd_sc_hd__mux4_1
X_2157_ FrameData[2] VGND VGND VPWR VPWR net210 sky130_fd_sc_hd__buf_1
XFILLER_13_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1390_ net413 _0617_ _0053_ _0240_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit22.Q Inst_LUT4AB_ConfigMem.Inst_frame13_bit23.Q
+ VGND VGND VPWR VPWR _0493_ sky130_fd_sc_hd__mux4_1
XFILLER_35_212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2011_ net750 net695 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1657_ net754 net726 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame13_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1588_ net39 net720 VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10
+ sky130_fd_sc_hd__dlxtp_1
X_1726_ net808 net737 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame11_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_73_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout626 H VGND VGND VPWR VPWR net626 sky130_fd_sc_hd__buf_2
Xfanout648 E VGND VGND VPWR VPWR net648 sky130_fd_sc_hd__buf_6
Xfanout637 net638 VGND VGND VPWR VPWR net637 sky130_fd_sc_hd__buf_4
Xfanout659 net663 VGND VGND VPWR VPWR net659 sky130_fd_sc_hd__buf_8
X_2209_ Inst_LUT4AB_switch_matrix.N1BEG2 VGND VGND VPWR VPWR net242 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_56_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_26 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0890_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit4.Q _0041_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit5.Q
+ VGND VGND VPWR VPWR _0042_ sky130_fd_sc_hd__a21o_1
Xoutput207 net207 VGND VGND VPWR VPWR FrameData_O[27] sky130_fd_sc_hd__buf_2
Xoutput229 net229 VGND VGND VPWR VPWR FrameStrobe_O[18] sky130_fd_sc_hd__buf_2
Xoutput218 net218 VGND VGND VPWR VPWR FrameData_O[8] sky130_fd_sc_hd__buf_2
X_1511_ net787 net704 VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9
+ sky130_fd_sc_hd__dlxtp_1
X_1442_ _0168_ _0093_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q VGND VGND VPWR VPWR
+ _0515_ sky130_fd_sc_hd__mux2_1
X_1373_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit4.Q _0475_ _0478_ _0479_ VGND VGND VPWR
+ VPWR _0480_ sky130_fd_sc_hd__o22a_1
XFILLER_67_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_18_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1709_ net774 net734 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame12_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_69_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1991_ net788 net692 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0942_ net87 net113 net95 net666 Inst_LUT4AB_ConfigMem.Inst_frame4_bit15.Q Inst_LUT4AB_ConfigMem.Inst_frame4_bit14.Q
+ VGND VGND VPWR VPWR _0090_ sky130_fd_sc_hd__mux4_1
X_0873_ Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 _0022_ _0023_ Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8
+ _0025_ VGND VGND VPWR VPWR _0026_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_15_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1425_ net61 net80 net134 net632 Inst_LUT4AB_ConfigMem.Inst_frame14_bit30.Q Inst_LUT4AB_ConfigMem.Inst_frame14_bit31.Q
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.N4BEG2 sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_66_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1356_ net666 net424 Inst_LUT4AB_ConfigMem.Inst_frame12_bit26.Q VGND VGND VPWR VPWR
+ _0465_ sky130_fd_sc_hd__mux2_1
X_1287_ net82 net7 net815 net813 Inst_LUT4AB_ConfigMem.Inst_frame3_bit27.Q Inst_LUT4AB_ConfigMem.Inst_frame3_bit26.Q
+ VGND VGND VPWR VPWR _0408_ sky130_fd_sc_hd__mux4_1
XFILLER_36_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2190_ net693 VGND VGND VPWR VPWR net233 sky130_fd_sc_hd__buf_1
X_1141_ _0274_ _0273_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit20.Q VGND VGND VPWR VPWR
+ _0275_ sky130_fd_sc_hd__mux2_4
X_1072_ _0209_ _0208_ VGND VGND VPWR VPWR _0210_ sky130_fd_sc_hd__nor2_4
XFILLER_49_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1210_ Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 _0074_ _0075_ Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15
+ _0339_ VGND VGND VPWR VPWR _0340_ sky130_fd_sc_hd__o221a_1
XFILLER_18_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1974_ net759 net694 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0925_ _0071_ _0072_ _0063_ _0062_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit5.Q Inst_LUT4AB_ConfigMem.Inst_frame9_bit6.Q
+ VGND VGND VPWR VPWR _0073_ sky130_fd_sc_hd__mux4_2
X_0787_ net814 net91 net119 net133 Inst_LUT4AB_ConfigMem.Inst_frame5_bit30.Q Inst_LUT4AB_ConfigMem.Inst_frame5_bit31.Q
+ VGND VGND VPWR VPWR _0635_ sky130_fd_sc_hd__mux4_1
X_0856_ _0628_ _0629_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit13.Q VGND VGND VPWR VPWR
+ _0009_ sky130_fd_sc_hd__mux2_1
X_1408_ net663 _0653_ Inst_LUT4AB_switch_matrix.JS2BEG2 _0639_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit12.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame11_bit13.Q VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.W1BEG3
+ sky130_fd_sc_hd__mux4_2
X_1339_ _0449_ _0450_ _0451_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit15.Q Inst_LUT4AB_ConfigMem.Inst_frame11_bit16.Q
+ VGND VGND VPWR VPWR _0452_ sky130_fd_sc_hd__a221o_1
XFILLER_28_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_203 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput390 net390 VGND VGND VPWR VPWR WW4BEG[7] sky130_fd_sc_hd__buf_2
XFILLER_19_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1690_ net51 net733 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame12_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_51_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0710_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit9.Q VGND VGND VPWR VPWR _0561_ sky130_fd_sc_hd__inv_1
X_2311_ clknet_1_0__leaf_UserCLK VGND VGND VPWR VPWR net344 sky130_fd_sc_hd__buf_2
XFILLER_38_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2242_ Inst_LUT4AB_switch_matrix.N4BEG3 VGND VGND VPWR VPWR net266 sky130_fd_sc_hd__clkbuf_2
X_1124_ _0258_ _0257_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit20.Q VGND VGND VPWR VPWR
+ _0259_ sky130_fd_sc_hd__mux2_4
XPHY_EDGE_ROW_69_Left_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2173_ net793 VGND VGND VPWR VPWR net197 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_48_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1055_ Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 _0081_ _0172_ Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10
+ VGND VGND VPWR VPWR _0194_ sky130_fd_sc_hd__a22o_1
X_1957_ net794 net688 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_33_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_31_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0908_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit4.Q _0057_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit5.Q
+ VGND VGND VPWR VPWR _0058_ sky130_fd_sc_hd__a21bo_1
X_1888_ net804 net679 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame6_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0839_ net77 net814 net105 Inst_LUT4AB_switch_matrix.JW2BEG1 Inst_LUT4AB_ConfigMem.Inst_frame0_bit0.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame0_bit1.Q VGND VGND VPWR VPWR _0682_ sky130_fd_sc_hd__mux4_2
Xinput107 S4END[2] VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__buf_2
XFILLER_56_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput129 W2MID[4] VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__buf_2
Xinput118 W2END[1] VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__buf_2
XFILLER_24_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_91 net772 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_80 _0063_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1811_ net811 net671 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame8_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_15_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1673_ net784 net727 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame13_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1742_ net773 net735 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame11_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
Xfanout808 net30 VGND VGND VPWR VPWR net808 sky130_fd_sc_hd__clkbuf_4
X_2225_ net75 VGND VGND VPWR VPWR net258 sky130_fd_sc_hd__clkbuf_2
X_2156_ net789 VGND VGND VPWR VPWR net199 sky130_fd_sc_hd__buf_1
XFILLER_53_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2087_ net788 net746 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame0_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_36_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1038_ net108 net120 net112 net134 Inst_LUT4AB_ConfigMem.Inst_frame1_bit3.Q Inst_LUT4AB_ConfigMem.Inst_frame1_bit2.Q
+ VGND VGND VPWR VPWR _0179_ sky130_fd_sc_hd__mux4_1
X_1107_ net23 net106 net138 Inst_LUT4AB_switch_matrix.JS2BEG4 Inst_LUT4AB_ConfigMem.Inst_frame0_bit22.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame0_bit23.Q VGND VGND VPWR VPWR _0243_ sky130_fd_sc_hd__mux4_2
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_59_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2010_ net752 net696 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1725_ net810 net737 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame11_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1656_ net756 net726 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame13_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1587_ net811 net720 VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9
+ sky130_fd_sc_hd__dlxtp_1
Xfanout627 net628 VGND VGND VPWR VPWR net627 sky130_fd_sc_hd__buf_6
Xfanout638 D VGND VGND VPWR VPWR net638 sky130_fd_sc_hd__buf_6
Xfanout649 net651 VGND VGND VPWR VPWR net649 sky130_fd_sc_hd__buf_4
XFILLER_37_28 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2208_ Inst_LUT4AB_switch_matrix.N1BEG1 VGND VGND VPWR VPWR net241 sky130_fd_sc_hd__buf_4
X_2139_ EE4END[4] VGND VGND VPWR VPWR net172 sky130_fd_sc_hd__clkbuf_1
XFILLER_53_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_4_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput208 net208 VGND VGND VPWR VPWR FrameData_O[28] sky130_fd_sc_hd__buf_2
XFILLER_64_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput219 net219 VGND VGND VPWR VPWR FrameData_O[9] sky130_fd_sc_hd__buf_2
XFILLER_4_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1510_ net791 net705 VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8
+ sky130_fd_sc_hd__dlxtp_1
X_1441_ _0237_ _0629_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q VGND VGND VPWR VPWR
+ _0514_ sky130_fd_sc_hd__mux2_1
X_1372_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit3.Q _0476_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit4.Q
+ VGND VGND VPWR VPWR _0479_ sky130_fd_sc_hd__a21bo_1
XFILLER_67_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_308 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_61_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1708_ net777 net731 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame12_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_69_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1639_ net788 net721 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame14_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_54_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_32_Left_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1990_ net792 net692 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0941_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit16.Q _0088_ VGND VGND VPWR VPWR _0089_
+ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_15_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_41_Left_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0872_ Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 _0018_ _0019_ Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12
+ VGND VGND VPWR VPWR _0025_ sky130_fd_sc_hd__o22a_1
XPHY_EDGE_ROW_50_Left_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1355_ net59 Inst_LUT4AB_ConfigMem.Inst_frame12_bit26.Q Inst_LUT4AB_ConfigMem.Inst_frame12_bit27.Q
+ VGND VGND VPWR VPWR _0464_ sky130_fd_sc_hd__o21ba_1
X_1424_ net62 net133 net77 net625 Inst_LUT4AB_ConfigMem.Inst_frame13_bit1.Q Inst_LUT4AB_ConfigMem.Inst_frame13_bit0.Q
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.N4BEG3 sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_66_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1286_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit28.Q _0404_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit29.Q
+ VGND VGND VPWR VPWR _0407_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_6_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_29_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1140_ net662 net656 net652 net636 Inst_LUT4AB_ConfigMem.Inst_frame1_bit18.Q Inst_LUT4AB_ConfigMem.Inst_frame1_bit19.Q
+ VGND VGND VPWR VPWR _0274_ sky130_fd_sc_hd__mux4_1
X_1071_ _0119_ _0120_ _0111_ _0110_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit23.Q Inst_LUT4AB_ConfigMem.Inst_frame9_bit24.Q
+ VGND VGND VPWR VPWR _0209_ sky130_fd_sc_hd__mux4_2
XFILLER_60_163 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1973_ net765 net694 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0924_ net74 net19 net102 net130 Inst_LUT4AB_ConfigMem.Inst_frame6_bit6.Q Inst_LUT4AB_ConfigMem.Inst_frame6_bit7.Q
+ VGND VGND VPWR VPWR _0072_ sky130_fd_sc_hd__mux4_1
X_0786_ _0632_ _0633_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit0.Q VGND VGND VPWR VPWR
+ _0634_ sky130_fd_sc_hd__mux2_4
X_0855_ _0640_ _0639_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit13.Q VGND VGND VPWR VPWR
+ _0008_ sky130_fd_sc_hd__mux2_4
X_1407_ _0505_ _0504_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit4.Q VGND VGND VPWR VPWR
+ Inst_LUT4AB_switch_matrix.NN4BEG0 sky130_fd_sc_hd__mux2_1
X_1338_ net666 net642 Inst_LUT4AB_ConfigMem.Inst_frame11_bit14.Q VGND VGND VPWR VPWR
+ _0451_ sky130_fd_sc_hd__mux2_1
X_1269_ net632 net627 _0392_ VGND VGND VPWR VPWR _0393_ sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_26_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput391 net391 VGND VGND VPWR VPWR WW4BEG[8] sky130_fd_sc_hd__buf_2
Xoutput380 net380 VGND VGND VPWR VPWR WW4BEG[12] sky130_fd_sc_hd__buf_4
XFILLER_42_163 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2310_ Inst_LUT4AB_switch_matrix.SS4BEG3 VGND VGND VPWR VPWR net334 sky130_fd_sc_hd__buf_6
X_2172_ net796 VGND VGND VPWR VPWR net196 sky130_fd_sc_hd__buf_1
X_1123_ net661 net658 net653 net638 Inst_LUT4AB_ConfigMem.Inst_frame3_bit18.Q Inst_LUT4AB_ConfigMem.Inst_frame3_bit19.Q
+ VGND VGND VPWR VPWR _0258_ sky130_fd_sc_hd__mux4_1
XFILLER_65_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1054_ _0191_ _0192_ _0183_ _0182_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit29.Q Inst_LUT4AB_ConfigMem.Inst_frame10_bit30.Q
+ VGND VGND VPWR VPWR _0193_ sky130_fd_sc_hd__mux4_1
X_1956_ net795 net688 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_33_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0907_ net424 net630 net626 net623 Inst_LUT4AB_ConfigMem.Inst_frame2_bit2.Q Inst_LUT4AB_ConfigMem.Inst_frame2_bit3.Q
+ VGND VGND VPWR VPWR _0057_ sky130_fd_sc_hd__mux4_1
X_1887_ net806 net679 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame6_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput108 S4END[3] VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__clkbuf_2
X_0838_ _0677_ _0562_ _0679_ _0681_ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.JW2BEG1
+ sky130_fd_sc_hd__o22a_4
X_0769_ _0554_ _0617_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit6.Q VGND VGND VPWR VPWR
+ _0618_ sky130_fd_sc_hd__o21ba_1
XFILLER_56_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput119 W2END[2] VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__buf_2
XFILLER_24_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_92 net772 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_81 _0120_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_70 net362 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1810_ net762 net669 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_30_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1741_ net776 net735 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame11_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_7_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout809 net810 VGND VGND VPWR VPWR net809 sky130_fd_sc_hd__buf_4
X_1672_ net785 net728 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame13_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2155_ net811 VGND VGND VPWR VPWR net188 sky130_fd_sc_hd__buf_1
X_1106_ _0241_ _0229_ Inst_LG_LUT4c_frame_config_dffesr.c_I0mux VGND VGND VPWR VPWR
+ _0242_ sky130_fd_sc_hd__mux2_4
X_2224_ net74 VGND VGND VPWR VPWR net257 sky130_fd_sc_hd__clkbuf_2
XFILLER_38_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2086_ net38 net746 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame0_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_42_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1037_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit4.Q _0175_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit5.Q
+ VGND VGND VPWR VPWR _0178_ sky130_fd_sc_hd__a21bo_1
XFILLER_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f_UserCLK_regs clknet_0_UserCLK_regs VGND VGND VPWR VPWR clknet_1_0__leaf_UserCLK_regs
+ sky130_fd_sc_hd__clkbuf_16
Xinput90 S2END[1] VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__buf_2
X_1939_ net812 net687 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_21_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1724_ net748 net737 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame11_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1655_ net758 net727 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame13_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
Xfanout628 H VGND VGND VPWR VPWR net628 sky130_fd_sc_hd__buf_8
X_1586_ net762 net716 VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8
+ sky130_fd_sc_hd__dlxtp_1
Xfanout639 net640 VGND VGND VPWR VPWR net639 sky130_fd_sc_hd__buf_6
X_2069_ net766 net745 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame0_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2207_ Inst_LUT4AB_switch_matrix.N1BEG0 VGND VGND VPWR VPWR net240 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_4_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1371_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit3.Q _0477_ VGND VGND VPWR VPWR _0478_
+ sky130_fd_sc_hd__and2b_1
Xoutput209 net209 VGND VGND VPWR VPWR FrameData_O[29] sky130_fd_sc_hd__buf_2
X_1440_ _0597_ _0512_ _0509_ VGND VGND VPWR VPWR _0513_ sky130_fd_sc_hd__o21ai_4
XFILLER_67_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_61_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1638_ net792 net721 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame14_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1707_ net779 net731 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame12_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_69_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1569_ net801 net713 VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_52_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0940_ net59 net67 net816 net12 Inst_LUT4AB_ConfigMem.Inst_frame4_bit14.Q Inst_LUT4AB_ConfigMem.Inst_frame4_bit15.Q
+ VGND VGND VPWR VPWR _0088_ sky130_fd_sc_hd__mux4_1
XFILLER_54_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0871_ Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 _0022_ _0023_ Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0
+ _0020_ VGND VGND VPWR VPWR _0024_ sky130_fd_sc_hd__o221a_1
X_1354_ net816 Inst_LUT4AB_ConfigMem.Inst_frame12_bit26.Q VGND VGND VPWR VPWR _0463_
+ sky130_fd_sc_hd__nand2b_1
X_1423_ net635 Inst_LUT4AB_switch_matrix.JN2BEG3 _0192_ _0043_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit15.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame13_bit14.Q VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.E1BEG0
+ sky130_fd_sc_hd__mux4_2
X_1285_ _0405_ _0589_ VGND VGND VPWR VPWR _0406_ sky130_fd_sc_hd__or2_4
XFILLER_36_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_29_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1070_ net431 _0108_ _0099_ _0098_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit25.Q Inst_LUT4AB_ConfigMem.Inst_frame9_bit26.Q
+ VGND VGND VPWR VPWR _0208_ sky130_fd_sc_hd__mux4_2
XFILLER_33_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0923_ net73 net18 net101 Inst_LUT4AB_switch_matrix.JS2BEG4 Inst_LUT4AB_ConfigMem.Inst_frame7_bit6.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame7_bit7.Q VGND VGND VPWR VPWR _0071_ sky130_fd_sc_hd__mux4_2
X_1972_ net790 net694 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0854_ _0696_ Inst_LA_LUT4c_frame_config_dffesr.LUT_flop Inst_LA_LUT4c_frame_config_dffesr.c_out_mux
+ VGND VGND VPWR VPWR A sky130_fd_sc_hd__mux2_4
XPHY_EDGE_ROW_23_Left_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_49_Right_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0785_ net639 net629 net624 net403 Inst_LUT4AB_ConfigMem.Inst_frame5_bit30.Q Inst_LUT4AB_ConfigMem.Inst_frame5_bit31.Q
+ VGND VGND VPWR VPWR _0633_ sky130_fd_sc_hd__mux4_2
X_1268_ _0391_ _0328_ Inst_LUT4AB_ConfigMem.Inst_frame14_bit16.Q VGND VGND VPWR VPWR
+ _0392_ sky130_fd_sc_hd__mux2_4
XFILLER_68_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1337_ net59 Inst_LUT4AB_ConfigMem.Inst_frame11_bit14.Q Inst_LUT4AB_ConfigMem.Inst_frame11_bit15.Q
+ VGND VGND VPWR VPWR _0450_ sky130_fd_sc_hd__o21ba_1
X_1406_ net59 net666 net816 net642 Inst_LUT4AB_ConfigMem.Inst_frame13_bit3.Q Inst_LUT4AB_ConfigMem.Inst_frame13_bit2.Q
+ VGND VGND VPWR VPWR _0505_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_58_Right_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_186 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1199_ _0167_ _0168_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit1.Q VGND VGND VPWR VPWR
+ _0329_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_67_Right_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_34_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput392 net392 VGND VGND VPWR VPWR WW4BEG[9] sky130_fd_sc_hd__buf_2
Xoutput381 Inst_LUT4AB_switch_matrix.WW4BEG1 VGND VGND VPWR VPWR WW4BEG[13] sky130_fd_sc_hd__buf_8
Xoutput370 net370 VGND VGND VPWR VPWR W6BEG[3] sky130_fd_sc_hd__buf_2
XFILLER_59_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1122_ net647 net628 net643 net404 Inst_LUT4AB_ConfigMem.Inst_frame3_bit19.Q Inst_LUT4AB_ConfigMem.Inst_frame3_bit18.Q
+ VGND VGND VPWR VPWR _0257_ sky130_fd_sc_hd__mux4_2
X_2171_ net798 VGND VGND VPWR VPWR net195 sky130_fd_sc_hd__clkbuf_1
XFILLER_65_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_142 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1053_ net70 net15 net98 net126 Inst_LUT4AB_ConfigMem.Inst_frame6_bit8.Q Inst_LUT4AB_ConfigMem.Inst_frame6_bit9.Q
+ VGND VGND VPWR VPWR _0192_ sky130_fd_sc_hd__mux4_2
XFILLER_21_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1955_ net797 net688 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_31_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0906_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit4.Q _0055_ VGND VGND VPWR VPWR _0056_
+ sky130_fd_sc_hd__and2b_1
X_1886_ net807 net682 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame6_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0837_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit0.Q _0680_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit1.Q
+ VGND VGND VPWR VPWR _0681_ sky130_fd_sc_hd__a21o_1
Xinput109 SS4END[0] VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__clkbuf_2
X_0768_ net72 net17 net100 net128 Inst_LUT4AB_ConfigMem.Inst_frame7_bit28.Q Inst_LUT4AB_ConfigMem.Inst_frame7_bit29.Q
+ VGND VGND VPWR VPWR _0617_ sky130_fd_sc_hd__mux4_2
X_0699_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit1.Q VGND VGND VPWR VPWR _0550_ sky130_fd_sc_hd__inv_1
XTAP_TAPCELL_ROW_39_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_82 _0120_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_60 net302 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_71 net364 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_93 net782 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_186 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1740_ net778 net736 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame11_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1671_ net787 net728 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame13_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1105_ _0237_ _0238_ _0240_ _0239_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit31.Q Inst_LUT4AB_ConfigMem.Inst_frame8_bit0.Q
+ VGND VGND VPWR VPWR _0241_ sky130_fd_sc_hd__mux4_1
X_2085_ net37 net746 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame0_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_36_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2223_ net73 VGND VGND VPWR VPWR net256 sky130_fd_sc_hd__buf_1
XFILLER_61_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1036_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit4.Q _0176_ VGND VGND VPWR VPWR _0177_
+ sky130_fd_sc_hd__and2b_1
Xinput91 S2END[2] VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__buf_2
X_1869_ net774 net678 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame7_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput80 N4END[3] VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__clkbuf_2
X_1938_ net761 net683 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame5_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_10_Left_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_42_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_218 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1654_ net759 net726 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame13_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_7_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1723_ net750 net737 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame11_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1585_ net764 net716 VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7
+ sky130_fd_sc_hd__dlxtp_1
X_2206_ net55 VGND VGND VPWR VPWR net230 sky130_fd_sc_hd__clkbuf_2
Xfanout629 net630 VGND VGND VPWR VPWR net629 sky130_fd_sc_hd__buf_2
X_1019_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit12.Q _0160_ VGND VGND VPWR VPWR _0161_
+ sky130_fd_sc_hd__and2b_1
XFILLER_53_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_259 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2068_ net790 net744 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame0_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_1_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_4_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1370_ net653 net638 Inst_LUT4AB_ConfigMem.Inst_frame12_bit2.Q VGND VGND VPWR VPWR
+ _0477_ sky130_fd_sc_hd__mux2_1
XFILLER_4_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1706_ net782 net732 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame12_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1637_ net794 net721 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame14_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_69_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1568_ net804 net712 VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9
+ sky130_fd_sc_hd__dlxtp_1
X_1499_ net749 net704 VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.c_out_mux
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_52_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_255 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0870_ _0016_ _0017_ VGND VGND VPWR VPWR _0023_ sky130_fd_sc_hd__or2_2
X_1422_ net645 _0093_ Inst_LUT4AB_switch_matrix.JN2BEG0 _0098_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit16.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame13_bit17.Q VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.E1BEG1
+ sky130_fd_sc_hd__mux4_1
X_1353_ net399 _0617_ _0053_ _0272_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit26.Q Inst_LUT4AB_ConfigMem.Inst_frame12_bit27.Q
+ VGND VGND VPWR VPWR _0462_ sky130_fd_sc_hd__mux4_1
X_1284_ net639 net629 net624 net416 Inst_LUT4AB_ConfigMem.Inst_frame3_bit26.Q Inst_LUT4AB_ConfigMem.Inst_frame3_bit27.Q
+ VGND VGND VPWR VPWR _0405_ sky130_fd_sc_hd__mux4_2
XFILLER_36_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0999_ Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 _0124_ _0141_ _0142_
+ VGND VGND VPWR VPWR _0143_ sky130_fd_sc_hd__o211a_1
XFILLER_3_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout790 net39 VGND VGND VPWR VPWR net790 sky130_fd_sc_hd__clkbuf_4
XFILLER_45_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_150 net57 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0922_ _0066_ _0566_ _0068_ _0070_ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.JS2BEG4
+ sky130_fd_sc_hd__o22a_4
X_1971_ net812 net694 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0853_ _0695_ _0688_ _0684_ VGND VGND VPWR VPWR _0696_ sky130_fd_sc_hd__mux2_4
X_1405_ net413 _0617_ _0053_ _0256_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit2.Q Inst_LUT4AB_ConfigMem.Inst_frame13_bit3.Q
+ VGND VGND VPWR VPWR _0504_ sky130_fd_sc_hd__mux4_1
X_0784_ net659 net634 net649 net645 Inst_LUT4AB_ConfigMem.Inst_frame5_bit31.Q Inst_LUT4AB_ConfigMem.Inst_frame5_bit30.Q
+ VGND VGND VPWR VPWR _0632_ sky130_fd_sc_hd__mux4_1
X_1267_ _0390_ net412 Inst_LUT4AB_ConfigMem.Inst_frame14_bit17.Q VGND VGND VPWR VPWR
+ _0391_ sky130_fd_sc_hd__mux2_4
XFILLER_68_232 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1198_ net647 net641 _0328_ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.M_EF sky130_fd_sc_hd__mux2_4
X_1336_ net87 Inst_LUT4AB_ConfigMem.Inst_frame11_bit14.Q VGND VGND VPWR VPWR _0449_
+ sky130_fd_sc_hd__nand2b_1
Xinput1 Ci VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__buf_6
XFILLER_51_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_34_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput371 net371 VGND VGND VPWR VPWR W6BEG[4] sky130_fd_sc_hd__buf_2
Xoutput360 net360 VGND VGND VPWR VPWR W2BEGb[3] sky130_fd_sc_hd__buf_2
Xoutput382 net382 VGND VGND VPWR VPWR WW4BEG[14] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_25_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_368 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_29_Left_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2170_ net799 VGND VGND VPWR VPWR net194 sky130_fd_sc_hd__buf_1
XFILLER_65_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1121_ net64 net109 net9 net120 Inst_LUT4AB_ConfigMem.Inst_frame5_bit21.Q Inst_LUT4AB_ConfigMem.Inst_frame5_bit20.Q
+ VGND VGND VPWR VPWR _0256_ sky130_fd_sc_hd__mux4_2
X_1052_ net69 net97 net125 Inst_LUT4AB_switch_matrix.JW2BEG4 Inst_LUT4AB_ConfigMem.Inst_frame7_bit8.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame7_bit9.Q VGND VGND VPWR VPWR _0191_ sky130_fd_sc_hd__mux4_2
X_1954_ net800 net688 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_38_Left_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_47_Left_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_31_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0905_ net659 net655 net635 net648 Inst_LUT4AB_ConfigMem.Inst_frame2_bit2.Q Inst_LUT4AB_ConfigMem.Inst_frame2_bit3.Q
+ VGND VGND VPWR VPWR _0055_ sky130_fd_sc_hd__mux4_2
X_1885_ net809 net682 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame6_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0836_ net91 net119 net107 net133 Inst_LUT4AB_ConfigMem.Inst_frame2_bit31.Q Inst_LUT4AB_ConfigMem.Inst_frame2_bit30.Q
+ VGND VGND VPWR VPWR _0680_ sky130_fd_sc_hd__mux4_1
X_0767_ net16 net99 net127 Inst_LUT4AB_switch_matrix.E2BEG3 Inst_LUT4AB_ConfigMem.Inst_frame8_bit28.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame8_bit29.Q VGND VGND VPWR VPWR _0616_ sky130_fd_sc_hd__mux4_2
X_0698_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit3.Q VGND VGND VPWR VPWR _0549_ sky130_fd_sc_hd__inv_2
X_2299_ SS4END[8] VGND VGND VPWR VPWR net338 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_56_Left_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_39_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1319_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit27.Q _0435_ VGND VGND VPWR VPWR _0436_
+ sky130_fd_sc_hd__and2b_1
XANTENNA_50 NN4END[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_83 _0120_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_61 net308 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_72 net370 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_94 net782 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput190 net190 VGND VGND VPWR VPWR FrameData_O[11] sky130_fd_sc_hd__buf_2
XFILLER_47_246 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f_UserCLK clknet_0_UserCLK VGND VGND VPWR VPWR clknet_1_0__leaf_UserCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_30_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_198 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1670_ net791 net728 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame13_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2222_ net72 VGND VGND VPWR VPWR net255 sky130_fd_sc_hd__buf_4
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1104_ net68 net13 net96 net135 Inst_LUT4AB_ConfigMem.Inst_frame5_bit18.Q Inst_LUT4AB_ConfigMem.Inst_frame5_bit19.Q
+ VGND VGND VPWR VPWR _0240_ sky130_fd_sc_hd__mux4_2
X_2153_ Inst_LUT4AB_switch_matrix.EE4BEG2 VGND VGND VPWR VPWR net177 sky130_fd_sc_hd__buf_1
X_1035_ net426 net655 net635 net648 Inst_LUT4AB_ConfigMem.Inst_frame1_bit2.Q Inst_LUT4AB_ConfigMem.Inst_frame1_bit3.Q
+ VGND VGND VPWR VPWR _0176_ sky130_fd_sc_hd__mux4_2
X_2084_ net795 net743 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame0_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1937_ net763 net683 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame5_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_21_135 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput92 S2END[3] VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__clkbuf_2
X_1799_ net787 net668 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1868_ net778 net675 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame7_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput81 NN4END[0] VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__clkbuf_2
Xinput70 N2MID[1] VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__clkbuf_2
X_0819_ Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14
+ _0643_ VGND VGND VPWR VPWR _0664_ sky130_fd_sc_hd__mux2_4
XFILLER_69_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_58_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1653_ net765 net727 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame13_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1584_ net45 net716 VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1722_ net752 net737 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame11_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_66_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2205_ net706 VGND VGND VPWR VPWR net229 sky130_fd_sc_hd__buf_1
X_2136_ E6END[11] VGND VGND VPWR VPWR net171 sky130_fd_sc_hd__clkbuf_2
X_1018_ net662 net656 net653 net636 Inst_LUT4AB_ConfigMem.Inst_frame4_bit10.Q Inst_LUT4AB_ConfigMem.Inst_frame4_bit11.Q
+ VGND VGND VPWR VPWR _0160_ sky130_fd_sc_hd__mux4_1
X_2067_ net812 net744 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame0_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_57_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclone40 Inst_LUT4AB_switch_matrix.M_EF VGND VGND VPWR VPWR net432 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_4_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1705_ net784 net732 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame12_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1636_ net795 net722 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame14_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1567_ net806 net712 VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8
+ sky130_fd_sc_hd__dlxtp_1
X_2119_ net14 VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__clkbuf_2
X_1498_ net751 net704 VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_1_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_77 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1421_ net424 Inst_LUT4AB_switch_matrix.JN2BEG1 net664 _0271_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit19.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame13_bit18.Q VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.E1BEG2
+ sky130_fd_sc_hd__mux4_2
XFILLER_48_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1283_ net430 net411 net649 net644 Inst_LUT4AB_ConfigMem.Inst_frame3_bit27.Q Inst_LUT4AB_ConfigMem.Inst_frame3_bit26.Q
+ VGND VGND VPWR VPWR _0404_ sky130_fd_sc_hd__mux4_1
X_1352_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit31.Q _0457_ _0460_ _0461_ VGND VGND
+ VPWR VPWR Inst_LUT4AB_switch_matrix.SS4BEG1 sky130_fd_sc_hd__o22a_1
XFILLER_36_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0998_ Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 _0125_ VGND VGND
+ VPWR VPWR _0142_ sky130_fd_sc_hd__or2_1
X_1619_ net811 net723 VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_54_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout780 net42 VGND VGND VPWR VPWR net780 sky130_fd_sc_hd__buf_4
Xfanout791 net792 VGND VGND VPWR VPWR net791 sky130_fd_sc_hd__clkbuf_4
XFILLER_1_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0921_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit12.Q _0069_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit13.Q
+ VGND VGND VPWR VPWR _0070_ sky130_fd_sc_hd__a21o_1
XFILLER_33_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_151 net57 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1970_ net761 net687 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
XANTENNA_140 net137 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0852_ _0694_ _0691_ _0663_ VGND VGND VPWR VPWR _0695_ sky130_fd_sc_hd__mux2_1
X_0783_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit3.Q _0628_ _0630_ VGND VGND VPWR VPWR
+ _0631_ sky130_fd_sc_hd__o21a_1
XFILLER_68_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1335_ net631 _0617_ _0053_ _0244_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit14.Q Inst_LUT4AB_ConfigMem.Inst_frame11_bit15.Q
+ VGND VGND VPWR VPWR _0448_ sky130_fd_sc_hd__mux4_1
X_1404_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit7.Q _0499_ _0501_ _0503_ VGND VGND VPWR
+ VPWR Inst_LUT4AB_switch_matrix.NN4BEG1 sky130_fd_sc_hd__o22a_1
X_1266_ _0389_ VGND VGND VPWR VPWR _0390_ sky130_fd_sc_hd__inv_2
X_1197_ _0326_ net396 Inst_LUT4AB_ConfigMem.Inst_frame14_bit17.Q VGND VGND VPWR VPWR
+ _0328_ sky130_fd_sc_hd__mux2_4
XFILLER_36_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput2 E1END[0] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_4
XFILLER_51_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput350 net350 VGND VGND VPWR VPWR W2BEG[1] sky130_fd_sc_hd__buf_6
XFILLER_10_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput361 net361 VGND VGND VPWR VPWR W2BEGb[4] sky130_fd_sc_hd__buf_2
XFILLER_59_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput383 Inst_LUT4AB_switch_matrix.WW4BEG3 VGND VGND VPWR VPWR WW4BEG[15] sky130_fd_sc_hd__buf_8
Xoutput372 net372 VGND VGND VPWR VPWR W6BEG[5] sky130_fd_sc_hd__buf_2
XFILLER_35_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_25_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1051_ _0567_ _0186_ _0188_ _0190_ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.JW2BEG4
+ sky130_fd_sc_hd__o22a_4
X_1120_ net79 net119 net111 Inst_LUT4AB_switch_matrix.E2BEG4 Inst_LUT4AB_ConfigMem.Inst_frame0_bit21.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame0_bit20.Q VGND VGND VPWR VPWR _0255_ sky130_fd_sc_hd__mux4_2
XFILLER_33_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1953_ net802 net688 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0904_ _0052_ _0053_ _0044_ _0043_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit3.Q Inst_LUT4AB_ConfigMem.Inst_frame9_bit4.Q
+ VGND VGND VPWR VPWR _0054_ sky130_fd_sc_hd__mux4_2
X_1884_ net748 net679 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame6_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_31_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0697_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit9.Q VGND VGND VPWR VPWR _0548_ sky130_fd_sc_hd__inv_1
X_0835_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit0.Q _0678_ VGND VGND VPWR VPWR _0679_
+ sky130_fd_sc_hd__and2b_1
X_0766_ _0612_ _0610_ _0615_ _0553_ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.E2BEG3
+ sky130_fd_sc_hd__a22o_4
X_2298_ SS4END[7] VGND VGND VPWR VPWR net337 sky130_fd_sc_hd__clkbuf_2
XFILLER_56_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1318_ net650 net411 Inst_LUT4AB_ConfigMem.Inst_frame11_bit26.Q VGND VGND VPWR VPWR
+ _0435_ sky130_fd_sc_hd__mux2_1
XFILLER_64_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1249_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit24.Q _0374_ VGND VGND VPWR VPWR _0375_
+ sky130_fd_sc_hd__nand2b_1
XANTENNA_51 NN4END[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_40 N4END[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_73 W6END[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_95 net784 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_84 _0120_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_62 net314 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput191 net191 VGND VGND VPWR VPWR FrameData_O[12] sky130_fd_sc_hd__buf_2
Xoutput180 net180 VGND VGND VPWR VPWR EE4BEG[2] sky130_fd_sc_hd__buf_2
XFILLER_47_258 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2221_ net71 VGND VGND VPWR VPWR net254 sky130_fd_sc_hd__clkbuf_2
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1103_ net80 net24 net108 Inst_LUT4AB_switch_matrix.JN2BEG4 Inst_LUT4AB_ConfigMem.Inst_frame0_bit18.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame0_bit19.Q VGND VGND VPWR VPWR _0239_ sky130_fd_sc_hd__mux4_2
X_1034_ net424 net399 net626 net432 Inst_LUT4AB_ConfigMem.Inst_frame1_bit2.Q Inst_LUT4AB_ConfigMem.Inst_frame1_bit3.Q
+ VGND VGND VPWR VPWR _0175_ sky130_fd_sc_hd__mux4_1
X_2083_ net797 net743 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame0_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1867_ net780 net675 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame7_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1936_ net768 net684 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame5_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_21_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput93 S2END[4] VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__buf_2
X_1798_ net791 net668 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput60 N1END[3] VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__clkbuf_4
Xinput82 NN4END[1] VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__clkbuf_2
Xinput71 N2MID[2] VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__buf_2
X_0749_ net640 net629 net626 net623 Inst_LUT4AB_ConfigMem.Inst_frame4_bit30.Q Inst_LUT4AB_ConfigMem.Inst_frame4_bit31.Q
+ VGND VGND VPWR VPWR _0600_ sky130_fd_sc_hd__mux4_1
X_0818_ _0652_ _0653_ _0662_ _0661_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit7.Q Inst_LUT4AB_ConfigMem.Inst_frame10_bit8.Q
+ VGND VGND VPWR VPWR _0663_ sky130_fd_sc_hd__mux4_2
XFILLER_52_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_58_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1721_ net754 net737 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame11_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1583_ net769 net716 VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5
+ sky130_fd_sc_hd__dlxtp_1
X_1652_ net790 net728 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame13_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2135_ E6END[10] VGND VGND VPWR VPWR net170 sky130_fd_sc_hd__clkbuf_2
X_2204_ net709 VGND VGND VPWR VPWR net228 sky130_fd_sc_hd__buf_1
X_1017_ net84 net95 net12 net123 Inst_LUT4AB_ConfigMem.Inst_frame5_bit3.Q Inst_LUT4AB_ConfigMem.Inst_frame5_bit2.Q
+ VGND VGND VPWR VPWR _0159_ sky130_fd_sc_hd__mux4_2
XFILLER_34_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2066_ net761 net699 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1919_ net805 net685 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame5_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_57_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1704_ net785 net730 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame12_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1635_ net797 net722 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame14_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1566_ net807 net712 VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7
+ sky130_fd_sc_hd__dlxtp_1
X_1497_ net753 net704 VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14
+ sky130_fd_sc_hd__dlxtp_1
X_2049_ net802 net701 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_39_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_1_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_52_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_9_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_89 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_63 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1351_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit30.Q _0458_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit31.Q
+ VGND VGND VPWR VPWR _0461_ sky130_fd_sc_hd__a21bo_1
X_1420_ net399 _0653_ Inst_LUT4AB_switch_matrix.JN2BEG2 _0639_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit20.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame13_bit21.Q VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.E1BEG3
+ sky130_fd_sc_hd__mux4_2
X_1282_ _0398_ _0400_ _0403_ _0588_ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.JW2BEG0
+ sky130_fd_sc_hd__a22o_1
XFILLER_63_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1618_ net762 net719 VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2
+ sky130_fd_sc_hd__dlxtp_1
X_0997_ Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 _0122_ _0126_ Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9
+ VGND VGND VPWR VPWR _0141_ sky130_fd_sc_hd__o22a_1
X_1549_ net775 net710 VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_54_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout781 FrameData[23] VGND VGND VPWR VPWR net781 sky130_fd_sc_hd__clkbuf_4
Xfanout792 net38 VGND VGND VPWR VPWR net792 sky130_fd_sc_hd__buf_4
Xfanout770 net44 VGND VGND VPWR VPWR net770 sky130_fd_sc_hd__buf_4
Xclkbuf_regs_0_UserCLK UserCLK VGND VGND VPWR VPWR UserCLK_regs sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_71_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0920_ net86 net94 net114 net116 Inst_LUT4AB_ConfigMem.Inst_frame2_bit10.Q Inst_LUT4AB_ConfigMem.Inst_frame2_bit11.Q
+ VGND VGND VPWR VPWR _0069_ sky130_fd_sc_hd__mux4_1
XFILLER_45_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_130 net768 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_152 net57 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_141 net137 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_0851_ _0692_ _0693_ _0620_ VGND VGND VPWR VPWR _0694_ sky130_fd_sc_hd__mux2_1
X_0782_ _0549_ _0629_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit4.Q VGND VGND VPWR VPWR
+ _0630_ sky130_fd_sc_hd__o21ba_1
XFILLER_68_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1265_ _0586_ _0388_ _0387_ VGND VGND VPWR VPWR _0389_ sky130_fd_sc_hd__a21oi_2
X_1403_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit6.Q _0502_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit7.Q
+ VGND VGND VPWR VPWR _0503_ sky130_fd_sc_hd__a21bo_1
XFILLER_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1334_ _0447_ _0446_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit19.Q VGND VGND VPWR VPWR
+ Inst_LUT4AB_switch_matrix.WW4BEG1 sky130_fd_sc_hd__mux2_4
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1196_ Inst_LUT4AB_switch_matrix.JN2BEG4 Inst_LUT4AB_switch_matrix.JS2BEG4 Inst_LUT4AB_switch_matrix.E2BEG4
+ Inst_LUT4AB_switch_matrix.JW2BEG4 Inst_LUT4AB_ConfigMem.Inst_frame8_bit19.Q Inst_LUT4AB_ConfigMem.Inst_frame8_bit18.Q
+ VGND VGND VPWR VPWR _0327_ sky130_fd_sc_hd__mux4_2
XFILLER_36_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput3 E1END[1] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_34_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_36_Right_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput340 net340 VGND VGND VPWR VPWR SS4BEG[6] sky130_fd_sc_hd__buf_2
Xoutput351 net351 VGND VGND VPWR VPWR W2BEG[2] sky130_fd_sc_hd__buf_8
XFILLER_10_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput384 net384 VGND VGND VPWR VPWR WW4BEG[1] sky130_fd_sc_hd__buf_2
Xoutput362 net362 VGND VGND VPWR VPWR W2BEGb[5] sky130_fd_sc_hd__buf_2
Xoutput373 net373 VGND VGND VPWR VPWR W6BEG[6] sky130_fd_sc_hd__buf_2
XFILLER_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_45_Right_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_25_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_54_Right_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_63_Right_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1050_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit12.Q _0189_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit13.Q
+ VGND VGND VPWR VPWR _0190_ sky130_fd_sc_hd__a21o_1
X_1952_ net803 net688 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0903_ net72 net17 net100 net128 Inst_LUT4AB_ConfigMem.Inst_frame6_bit4.Q Inst_LUT4AB_ConfigMem.Inst_frame6_bit5.Q
+ VGND VGND VPWR VPWR _0053_ sky130_fd_sc_hd__mux4_2
X_0834_ net57 net8 net63 net814 Inst_LUT4AB_ConfigMem.Inst_frame2_bit31.Q Inst_LUT4AB_ConfigMem.Inst_frame2_bit30.Q
+ VGND VGND VPWR VPWR _0678_ sky130_fd_sc_hd__mux4_1
X_1883_ net750 net679 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame6_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_72_Right_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0765_ _0613_ _0614_ _0552_ VGND VGND VPWR VPWR _0615_ sky130_fd_sc_hd__mux2_1
X_2297_ SS4END[6] VGND VGND VPWR VPWR net336 sky130_fd_sc_hd__clkbuf_2
X_1248_ net57 net81 net2 net6 Inst_LUT4AB_ConfigMem.Inst_frame1_bit22.Q Inst_LUT4AB_ConfigMem.Inst_frame1_bit23.Q
+ VGND VGND VPWR VPWR _0374_ sky130_fd_sc_hd__mux4_1
X_1317_ net645 net640 Inst_LUT4AB_ConfigMem.Inst_frame11_bit26.Q VGND VGND VPWR VPWR
+ _0434_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_47_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1179_ _0280_ _0281_ _0272_ _0271_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit15.Q Inst_LUT4AB_ConfigMem.Inst_frame8_bit16.Q
+ VGND VGND VPWR VPWR _0311_ sky130_fd_sc_hd__mux4_2
XFILLER_12_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_52 NN4END[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_41 N4END[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_74 _0053_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_85 _0120_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_30 FrameStrobe[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_63 net320 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_96 net788 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput192 net192 VGND VGND VPWR VPWR FrameData_O[13] sky130_fd_sc_hd__buf_2
Xoutput170 net170 VGND VGND VPWR VPWR E6BEG[8] sky130_fd_sc_hd__buf_2
Xoutput181 net181 VGND VGND VPWR VPWR EE4BEG[3] sky130_fd_sc_hd__buf_2
XFILLER_62_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_64 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2151_ Inst_LUT4AB_switch_matrix.EE4BEG0 VGND VGND VPWR VPWR net175 sky130_fd_sc_hd__clkbuf_1
XFILLER_38_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1102_ net76 net21 net104 net132 Inst_LUT4AB_ConfigMem.Inst_frame6_bit18.Q Inst_LUT4AB_ConfigMem.Inst_frame6_bit19.Q
+ VGND VGND VPWR VPWR _0238_ sky130_fd_sc_hd__mux4_2
X_2220_ net70 VGND VGND VPWR VPWR net253 sky130_fd_sc_hd__buf_4
X_2082_ net800 net743 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame0_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_53_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1033_ Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 _0079_ _0081_ Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15
+ _0173_ VGND VGND VPWR VPWR _0174_ sky130_fd_sc_hd__a221o_1
Xinput50 FrameData[6] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__buf_1
X_1866_ net781 net677 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame7_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1797_ net793 net667 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0817_ net65 net93 net24 net121 Inst_LUT4AB_ConfigMem.Inst_frame6_bit31.Q Inst_LUT4AB_ConfigMem.Inst_frame6_bit30.Q
+ VGND VGND VPWR VPWR _0662_ sky130_fd_sc_hd__mux4_2
Xinput61 N2END[0] VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__buf_2
Xinput72 N2MID[3] VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__clkbuf_2
X_1935_ net770 net684 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame5_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput94 S2END[5] VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__clkbuf_2
XFILLER_67_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput83 NN4END[2] VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__buf_1
X_0748_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit0.Q _0598_ VGND VGND VPWR VPWR _0599_
+ sky130_fd_sc_hd__or2_1
XFILLER_37_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2349_ WW4END[9] VGND VGND VPWR VPWR net388 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_58_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1720_ net755 net738 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame11_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1651_ net812 net728 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame13_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1582_ net771 net716 VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4
+ sky130_fd_sc_hd__dlxtp_1
X_2134_ E6END[9] VGND VGND VPWR VPWR net169 sky130_fd_sc_hd__buf_1
XFILLER_66_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2203_ FrameStrobe[16] VGND VGND VPWR VPWR net227 sky130_fd_sc_hd__buf_1
X_2065_ net763 net699 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_19_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1016_ net9 net137 net112 Inst_LUT4AB_switch_matrix.JN2BEG2 Inst_LUT4AB_ConfigMem.Inst_frame0_bit3.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame0_bit2.Q VGND VGND VPWR VPWR _0158_ sky130_fd_sc_hd__mux4_1
XFILLER_34_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_14_Left_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1918_ net808 net686 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame5_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1849_ net754 net677 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame7_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_72_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_55_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_232 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclone75 _0513_ VGND VGND VPWR VPWR net467 sky130_fd_sc_hd__buf_6
XFILLER_9_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1634_ net799 net724 VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.c_reset_value
+ sky130_fd_sc_hd__dlxtp_1
X_1703_ net787 net730 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame12_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1565_ net809 net712 VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6
+ sky130_fd_sc_hd__dlxtp_1
X_1496_ net755 net703 VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13
+ sky130_fd_sc_hd__dlxtp_1
X_2117_ Inst_LUT4AB_switch_matrix.E2BEG6 VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_52_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2048_ net803 net702 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_60_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1281_ _0401_ _0402_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit28.Q VGND VGND VPWR VPWR
+ _0403_ sky130_fd_sc_hd__mux2_1
X_1350_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit30.Q _0459_ VGND VGND VPWR VPWR _0460_
+ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_66_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0996_ _0138_ _0139_ _0130_ _0129_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit17.Q Inst_LUT4AB_ConfigMem.Inst_frame9_bit18.Q
+ VGND VGND VPWR VPWR _0140_ sky130_fd_sc_hd__mux4_2
X_1617_ net764 net719 VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1
+ sky130_fd_sc_hd__dlxtp_1
X_1479_ _0544_ VGND VGND VPWR VPWR _0545_ sky130_fd_sc_hd__inv_1
XFILLER_39_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1548_ net777 net709 VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_27_302 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0_UserCLK_regs UserCLK_regs VGND VGND VPWR VPWR clknet_0_UserCLK_regs sky130_fd_sc_hd__clkbuf_16
XFILLER_10_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_17_Left_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_20_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout760 net48 VGND VGND VPWR VPWR net760 sky130_fd_sc_hd__clkbuf_4
XFILLER_2_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout782 FrameData[23] VGND VGND VPWR VPWR net782 sky130_fd_sc_hd__buf_4
XANTENNA_120 net219 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout793 net794 VGND VGND VPWR VPWR net793 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_28_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout771 net773 VGND VGND VPWR VPWR net771 sky130_fd_sc_hd__clkbuf_4
XANTENNA_131 net786 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_142 net397 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_71_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_153 net57 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_198 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0850_ Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0
+ _0643_ VGND VGND VPWR VPWR _0693_ sky130_fd_sc_hd__mux2_1
X_1402_ _0071_ _0111_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit5.Q VGND VGND VPWR VPWR
+ _0502_ sky130_fd_sc_hd__mux2_4
X_0781_ net76 net21 net104 net132 Inst_LUT4AB_ConfigMem.Inst_frame7_bit26.Q Inst_LUT4AB_ConfigMem.Inst_frame7_bit27.Q
+ VGND VGND VPWR VPWR _0629_ sky130_fd_sc_hd__mux4_1
X_1264_ Inst_LUT4AB_switch_matrix.JN2BEG7 Inst_LUT4AB_switch_matrix.E2BEG7 Inst_LUT4AB_ConfigMem.Inst_frame8_bit24.Q
+ VGND VGND VPWR VPWR _0388_ sky130_fd_sc_hd__mux2_1
X_1333_ net60 net88 net665 net660 Inst_LUT4AB_ConfigMem.Inst_frame11_bit17.Q Inst_LUT4AB_ConfigMem.Inst_frame11_bit18.Q
+ VGND VGND VPWR VPWR _0447_ sky130_fd_sc_hd__mux4_1
Xinput4 E1END[2] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__buf_1
X_1195_ _0324_ _0325_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit23.Q VGND VGND VPWR VPWR
+ _0326_ sky130_fd_sc_hd__mux2_4
XFILLER_51_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0979_ _0109_ _0121_ VGND VGND VPWR VPWR _0124_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_34_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput374 net374 VGND VGND VPWR VPWR W6BEG[7] sky130_fd_sc_hd__buf_2
Xoutput352 net352 VGND VGND VPWR VPWR W2BEG[3] sky130_fd_sc_hd__buf_6
Xoutput330 net330 VGND VGND VPWR VPWR SS4BEG[11] sky130_fd_sc_hd__buf_2
Xoutput341 net341 VGND VGND VPWR VPWR SS4BEG[7] sky130_fd_sc_hd__buf_2
Xoutput363 net363 VGND VGND VPWR VPWR W2BEGb[6] sky130_fd_sc_hd__buf_2
Xoutput385 net385 VGND VGND VPWR VPWR WW4BEG[2] sky130_fd_sc_hd__buf_2
XFILLER_19_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_2_Left_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1951_ net805 net688 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0902_ net71 net127 net16 Inst_LUT4AB_switch_matrix.E2BEG4 Inst_LUT4AB_ConfigMem.Inst_frame7_bit5.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame7_bit4.Q VGND VGND VPWR VPWR _0052_ sky130_fd_sc_hd__mux4_2
X_1882_ net751 net681 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame6_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0833_ _0675_ _0676_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit0.Q VGND VGND VPWR VPWR
+ _0677_ sky130_fd_sc_hd__mux2_4
X_0764_ net59 net65 net77 net10 Inst_LUT4AB_ConfigMem.Inst_frame3_bit6.Q Inst_LUT4AB_ConfigMem.Inst_frame3_bit7.Q
+ VGND VGND VPWR VPWR _0614_ sky130_fd_sc_hd__mux4_1
X_1178_ _0305_ _0309_ _0300_ VGND VGND VPWR VPWR _0310_ sky130_fd_sc_hd__a21o_1
X_2296_ SS4END[5] VGND VGND VPWR VPWR net335 sky130_fd_sc_hd__clkbuf_2
XFILLER_56_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1247_ _0372_ _0371_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit24.Q VGND VGND VPWR VPWR
+ _0373_ sky130_fd_sc_hd__mux2_4
X_1316_ net815 net665 net426 net430 Inst_LUT4AB_ConfigMem.Inst_frame11_bit26.Q Inst_LUT4AB_ConfigMem.Inst_frame11_bit27.Q
+ VGND VGND VPWR VPWR _0433_ sky130_fd_sc_hd__mux4_1
XFILLER_64_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_31 FrameStrobe[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_20 EE4END[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_53 NN4END[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_42 N4END[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_97 net796 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_75 _0053_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_64 net321 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_86 _0662_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput193 net193 VGND VGND VPWR VPWR FrameData_O[14] sky130_fd_sc_hd__buf_2
Xoutput171 net171 VGND VGND VPWR VPWR E6BEG[9] sky130_fd_sc_hd__buf_2
Xoutput160 net160 VGND VGND VPWR VPWR E6BEG[0] sky130_fd_sc_hd__buf_2
Xoutput182 net182 VGND VGND VPWR VPWR EE4BEG[4] sky130_fd_sc_hd__buf_2
XFILLER_46_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2150_ EE4END[15] VGND VGND VPWR VPWR net174 sky130_fd_sc_hd__buf_1
X_1101_ net75 net103 net20 Inst_LUT4AB_switch_matrix.JN2BEG6 Inst_LUT4AB_ConfigMem.Inst_frame7_bit19.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame7_bit18.Q VGND VGND VPWR VPWR _0237_ sky130_fd_sc_hd__mux4_2
X_1032_ Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 _0171_ _0172_ Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11
+ VGND VGND VPWR VPWR _0173_ sky130_fd_sc_hd__a22o_1
X_2081_ net802 net743 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame0_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1934_ net773 net683 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame5_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput95 S2END[6] VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__clkbuf_2
Xinput40 FrameData[20] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__buf_1
Xinput51 FrameData[7] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__buf_1
X_1865_ net783 net677 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame7_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1796_ net36 net667 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput62 N2END[1] VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput73 N2MID[4] VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput84 NN4END[3] VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__dlymetal6s2s_1
X_0747_ net663 net635 net651 net644 Inst_LUT4AB_ConfigMem.Inst_frame4_bit31.Q Inst_LUT4AB_ConfigMem.Inst_frame4_bit30.Q
+ VGND VGND VPWR VPWR _0598_ sky130_fd_sc_hd__mux4_1
X_0816_ net78 net813 net134 Inst_LUT4AB_switch_matrix.JS2BEG1 Inst_LUT4AB_ConfigMem.Inst_frame1_bit30.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame1_bit31.Q VGND VGND VPWR VPWR _0661_ sky130_fd_sc_hd__mux4_2
XFILLER_69_374 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2348_ WW4END[8] VGND VGND VPWR VPWR net387 sky130_fd_sc_hd__clkbuf_2
X_2279_ S4END[4] VGND VGND VPWR VPWR net312 sky130_fd_sc_hd__clkbuf_2
XFILLER_29_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_274 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_41_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1581_ net775 net716 VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3
+ sky130_fd_sc_hd__dlxtp_1
X_1650_ net47 net722 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame14_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2202_ net719 VGND VGND VPWR VPWR net226 sky130_fd_sc_hd__clkbuf_1
X_2133_ E6END[8] VGND VGND VPWR VPWR net168 sky130_fd_sc_hd__buf_1
XFILLER_66_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1015_ _0153_ _0564_ _0156_ _0157_ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.JN2BEG2
+ sky130_fd_sc_hd__o22a_4
X_2064_ net767 net700 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1917_ net810 net685 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame5_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1848_ net49 net678 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame7_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1779_ net811 net670 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_4_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclone21 G VGND VGND VPWR VPWR net413 sky130_fd_sc_hd__clkbuf_1
XFILLER_43_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclone32 net643 VGND VGND VPWR VPWR net424 sky130_fd_sc_hd__clkbuf_1
XFILLER_68_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1633_ net801 net724 VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.c_I0mux
+ sky130_fd_sc_hd__dlxtp_1
X_1564_ net747 net713 VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5
+ sky130_fd_sc_hd__dlxtp_1
X_1702_ net792 net730 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame12_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_66_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1495_ net757 net703 VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12
+ sky130_fd_sc_hd__dlxtp_1
X_2116_ Inst_LUT4AB_switch_matrix.E2BEG5 VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__buf_1
XFILLER_54_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2047_ net805 net702 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_17_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_66_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1280_ net90 net118 net106 net134 Inst_LUT4AB_ConfigMem.Inst_frame2_bit27.Q Inst_LUT4AB_ConfigMem.Inst_frame2_bit26.Q
+ VGND VGND VPWR VPWR _0402_ sky130_fd_sc_hd__mux4_1
XFILLER_63_188 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0995_ net70 net15 net98 net126 Inst_LUT4AB_ConfigMem.Inst_frame6_bit16.Q Inst_LUT4AB_ConfigMem.Inst_frame6_bit17.Q
+ VGND VGND VPWR VPWR _0139_ sky130_fd_sc_hd__mux4_2
X_1616_ net767 net719 VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_59_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1547_ net779 net709 VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7
+ sky130_fd_sc_hd__dlxtp_1
X_1478_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit7.Q _0522_ VGND VGND VPWR VPWR _0544_
+ sky130_fd_sc_hd__nand2_1
XFILLER_27_358 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_314 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_20_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout783 FrameData[22] VGND VGND VPWR VPWR net783 sky130_fd_sc_hd__clkbuf_4
Xfanout750 net52 VGND VGND VPWR VPWR net750 sky130_fd_sc_hd__buf_4
Xfanout794 net37 VGND VGND VPWR VPWR net794 sky130_fd_sc_hd__buf_4
Xfanout772 net773 VGND VGND VPWR VPWR net772 sky130_fd_sc_hd__buf_2
Xfanout761 net762 VGND VGND VPWR VPWR net761 sky130_fd_sc_hd__clkbuf_4
XFILLER_65_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_143 net216 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_154 net57 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_132 net786 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_110 net111 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_121 FrameStrobe[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0780_ net75 net103 net131 Inst_LUT4AB_switch_matrix.JN2BEG3 Inst_LUT4AB_ConfigMem.Inst_frame8_bit26.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame8_bit27.Q VGND VGND VPWR VPWR _0628_ sky130_fd_sc_hd__mux4_2
X_1401_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit6.Q _0500_ VGND VGND VPWR VPWR _0501_
+ sky130_fd_sc_hd__and2b_1
X_1263_ Inst_LUT4AB_switch_matrix.JS2BEG7 Inst_LUT4AB_ConfigMem.Inst_frame8_bit24.Q
+ _0386_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit25.Q VGND VGND VPWR VPWR _0387_ sky130_fd_sc_hd__o211a_1
X_1194_ Inst_LUT4AB_switch_matrix.JS2BEG6 Inst_LUT4AB_switch_matrix.JW2BEG6 Inst_LUT4AB_ConfigMem.Inst_frame8_bit22.Q
+ VGND VGND VPWR VPWR _0325_ sky130_fd_sc_hd__mux2_1
X_1332_ net627 _0652_ _0071_ _0099_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit17.Q Inst_LUT4AB_ConfigMem.Inst_frame11_bit18.Q
+ VGND VGND VPWR VPWR _0446_ sky130_fd_sc_hd__mux4_2
XFILLER_36_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput5 E1END[3] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_51_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0978_ _0109_ _0121_ VGND VGND VPWR VPWR _0123_ sky130_fd_sc_hd__and2_1
Xoutput375 net375 VGND VGND VPWR VPWR W6BEG[8] sky130_fd_sc_hd__buf_2
Xoutput331 net331 VGND VGND VPWR VPWR SS4BEG[12] sky130_fd_sc_hd__buf_2
Xoutput342 net342 VGND VGND VPWR VPWR SS4BEG[8] sky130_fd_sc_hd__buf_2
Xoutput320 net320 VGND VGND VPWR VPWR S4BEG[2] sky130_fd_sc_hd__buf_2
Xoutput353 net353 VGND VGND VPWR VPWR W2BEG[4] sky130_fd_sc_hd__buf_8
Xoutput364 net364 VGND VGND VPWR VPWR W2BEGb[7] sky130_fd_sc_hd__buf_2
Xoutput386 net386 VGND VGND VPWR VPWR WW4BEG[3] sky130_fd_sc_hd__buf_2
XFILLER_19_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_25_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_280 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1950_ net808 net688 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_33_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0901_ _0048_ _0046_ _0051_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit13.Q VGND VGND VPWR
+ VPWR Inst_LUT4AB_switch_matrix.E2BEG4 sky130_fd_sc_hd__o22a_4
X_1881_ net753 net681 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame6_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0832_ net639 net629 net624 net416 Inst_LUT4AB_ConfigMem.Inst_frame2_bit30.Q Inst_LUT4AB_ConfigMem.Inst_frame2_bit31.Q
+ VGND VGND VPWR VPWR _0676_ sky130_fd_sc_hd__mux4_1
X_0763_ net814 net93 net121 net133 Inst_LUT4AB_ConfigMem.Inst_frame3_bit6.Q Inst_LUT4AB_ConfigMem.Inst_frame3_bit7.Q
+ VGND VGND VPWR VPWR _0613_ sky130_fd_sc_hd__mux4_1
XFILLER_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1315_ _0427_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit1.Q _0429_ _0432_ VGND VGND VPWR
+ VPWR Inst_LUT4AB_switch_matrix.W6BEG1 sky130_fd_sc_hd__a22o_1
X_2295_ SS4END[4] VGND VGND VPWR VPWR net328 sky130_fd_sc_hd__clkbuf_2
X_1177_ Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 _0307_ _0308_ Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2
+ VGND VGND VPWR VPWR _0309_ sky130_fd_sc_hd__o22a_1
XFILLER_64_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1246_ net660 net657 net652 net637 Inst_LUT4AB_ConfigMem.Inst_frame1_bit22.Q Inst_LUT4AB_ConfigMem.Inst_frame1_bit23.Q
+ VGND VGND VPWR VPWR _0372_ sky130_fd_sc_hd__mux4_1
XANTENNA_32 net221 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_10 E6END[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_54 NN4END[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_43 N4END[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_21 EE4END[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_65 net324 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_331 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput161 Inst_LUT4AB_switch_matrix.E6BEG0 VGND VGND VPWR VPWR E6BEG[10] sky130_fd_sc_hd__buf_8
Xoutput150 net150 VGND VGND VPWR VPWR E2BEG[6] sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_30_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_76 _0053_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_87 _0662_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_98 net804 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_386 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput194 net194 VGND VGND VPWR VPWR FrameData_O[15] sky130_fd_sc_hd__buf_2
Xoutput183 net183 VGND VGND VPWR VPWR EE4BEG[5] sky130_fd_sc_hd__buf_2
Xoutput172 net172 VGND VGND VPWR VPWR EE4BEG[0] sky130_fd_sc_hd__buf_2
XFILLER_55_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1100_ _0232_ _0563_ _0236_ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.JN2BEG6
+ sky130_fd_sc_hd__o21a_4
XFILLER_53_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1031_ _0078_ _0077_ VGND VGND VPWR VPWR _0172_ sky130_fd_sc_hd__and2b_1
X_2080_ net804 net743 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame0_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1933_ net776 net683 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame5_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput96 S2END[7] VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__clkbuf_2
Xinput85 S1END[0] VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__buf_2
Xinput41 FrameData[21] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__buf_1
Xinput52 FrameData[8] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__buf_1
Xinput30 FrameData[11] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__dlymetal6s2s_1
X_1864_ net785 net676 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame7_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1795_ net35 net669 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0815_ _0657_ _0655_ _0660_ _0560_ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.JS2BEG1
+ sky130_fd_sc_hd__a22o_1
Xinput74 N2MID[5] VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__buf_2
Xinput63 N2END[2] VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__dlymetal6s2s_1
X_0746_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit31.Q VGND VGND VPWR VPWR _0597_ sky130_fd_sc_hd__inv_2
X_2278_ net104 VGND VGND VPWR VPWR net311 sky130_fd_sc_hd__buf_1
X_2347_ WW4END[7] VGND VGND VPWR VPWR net386 sky130_fd_sc_hd__clkbuf_2
X_1229_ net647 net633 net643 net414 Inst_LUT4AB_ConfigMem.Inst_frame3_bit23.Q Inst_LUT4AB_ConfigMem.Inst_frame3_bit22.Q
+ VGND VGND VPWR VPWR _0357_ sky130_fd_sc_hd__mux4_2
XFILLER_52_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_35_Left_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1580_ net777 net716 VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_44_Left_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2132_ E6END[7] VGND VGND VPWR VPWR net167 sky130_fd_sc_hd__buf_1
X_2201_ net725 VGND VGND VPWR VPWR net225 sky130_fd_sc_hd__clkbuf_1
XFILLER_3_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_53_Left_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1014_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit4.Q _0154_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit5.Q
+ VGND VGND VPWR VPWR _0157_ sky130_fd_sc_hd__a21o_1
XFILLER_34_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2063_ net769 net700 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_62_Left_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1847_ net758 net678 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame7_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_34_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1916_ net748 net683 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame5_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0729_ Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 VGND VGND VPWR VPWR
+ _0580_ sky130_fd_sc_hd__inv_1
X_1778_ net761 net739 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame10_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_71_Left_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_231 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_286 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1701_ net794 net730 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame12_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1632_ net803 net725 VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.c_out_mux
+ sky130_fd_sc_hd__dlxtp_1
X_1563_ net749 net713 VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4
+ sky130_fd_sc_hd__dlxtp_1
X_1494_ net760 net706 VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_69_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2115_ Inst_LUT4AB_switch_matrix.E2BEG4 VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__clkbuf_2
XFILLER_39_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2046_ net808 net701 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0994_ net14 net97 net125 Inst_LUT4AB_switch_matrix.JW2BEG5 Inst_LUT4AB_ConfigMem.Inst_frame7_bit16.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame7_bit17.Q VGND VGND VPWR VPWR _0138_ sky130_fd_sc_hd__mux4_2
X_1615_ net44 net719 VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.c_reset_value
+ sky130_fd_sc_hd__dlxtp_1
X_1477_ _0542_ _0543_ net482 _0541_ VGND VGND VPWR VPWR _0006_ sky130_fd_sc_hd__a2bb2o_1
X_1546_ net782 net709 VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_27_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2029_ net776 net695 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_10_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_20_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout784 FrameData[22] VGND VGND VPWR VPWR net784 sky130_fd_sc_hd__buf_4
XFILLER_49_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout762 net47 VGND VGND VPWR VPWR net762 sky130_fd_sc_hd__buf_4
Xfanout773 FrameData[27] VGND VGND VPWR VPWR net773 sky130_fd_sc_hd__clkbuf_4
Xfanout751 net752 VGND VGND VPWR VPWR net751 sky130_fd_sc_hd__clkbuf_4
Xfanout740 net741 VGND VGND VPWR VPWR net740 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout795 net796 VGND VGND VPWR VPWR net795 sky130_fd_sc_hd__clkbuf_4
XANTENNA_122 net223 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_111 net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_133 net787 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_155 net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_144 net375 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_100 net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_11_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1400_ net410 _0652_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit5.Q VGND VGND VPWR VPWR
+ _0500_ sky130_fd_sc_hd__mux2_1
X_1331_ _0445_ _0444_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit22.Q VGND VGND VPWR VPWR
+ Inst_LUT4AB_switch_matrix.WW4BEG2 sky130_fd_sc_hd__mux2_1
X_1193_ Inst_LUT4AB_switch_matrix.JN2BEG6 Inst_LUT4AB_switch_matrix.E2BEG6 Inst_LUT4AB_ConfigMem.Inst_frame8_bit22.Q
+ VGND VGND VPWR VPWR _0324_ sky130_fd_sc_hd__mux2_4
X_1262_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit24.Q _0378_ VGND VGND VPWR VPWR _0386_
+ sky130_fd_sc_hd__nand2_2
Xinput6 E2END[0] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_2
X_0977_ _0109_ _0121_ VGND VGND VPWR VPWR _0122_ sky130_fd_sc_hd__nand2b_1
Xoutput332 Inst_LUT4AB_switch_matrix.SS4BEG1 VGND VGND VPWR VPWR SS4BEG[13] sky130_fd_sc_hd__buf_6
Xoutput343 net343 VGND VGND VPWR VPWR SS4BEG[9] sky130_fd_sc_hd__buf_2
Xoutput321 net321 VGND VGND VPWR VPWR S4BEG[3] sky130_fd_sc_hd__buf_2
Xoutput310 net310 VGND VGND VPWR VPWR S2BEGb[6] sky130_fd_sc_hd__buf_2
Xoutput376 net376 VGND VGND VPWR VPWR W6BEG[9] sky130_fd_sc_hd__buf_2
X_1529_ net753 net707 VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8
+ sky130_fd_sc_hd__dlxtp_1
Xoutput354 net429 VGND VGND VPWR VPWR W2BEG[5] sky130_fd_sc_hd__buf_6
Xoutput387 net387 VGND VGND VPWR VPWR WW4BEG[4] sky130_fd_sc_hd__buf_2
Xoutput365 net365 VGND VGND VPWR VPWR W6BEG[0] sky130_fd_sc_hd__buf_2
XFILLER_67_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_25_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_33_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0900_ _0050_ _0049_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit12.Q VGND VGND VPWR VPWR
+ _0051_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_32_Right_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1880_ net755 net679 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame6_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0831_ net426 net634 net649 net644 Inst_LUT4AB_ConfigMem.Inst_frame2_bit31.Q Inst_LUT4AB_ConfigMem.Inst_frame2_bit30.Q
+ VGND VGND VPWR VPWR _0675_ sky130_fd_sc_hd__mux4_2
X_0762_ _0552_ _0611_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit9.Q VGND VGND VPWR VPWR
+ _0612_ sky130_fd_sc_hd__o21a_1
XFILLER_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_41_Right_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1314_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit0.Q _0431_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit1.Q
+ VGND VGND VPWR VPWR _0432_ sky130_fd_sc_hd__a21oi_1
X_2294_ Inst_LUT4AB_switch_matrix.S4BEG3 VGND VGND VPWR VPWR net318 sky130_fd_sc_hd__clkbuf_1
X_1176_ _0301_ _0302_ VGND VGND VPWR VPWR _0308_ sky130_fd_sc_hd__nand2b_1
Xclkbuf_1_1__f_UserCLK_regs clknet_0_UserCLK_regs VGND VGND VPWR VPWR clknet_1_1__leaf_UserCLK_regs
+ sky130_fd_sc_hd__clkbuf_16
XPHY_EDGE_ROW_50_Right_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1245_ net646 net631 net641 Inst_LUT4AB_switch_matrix.M_AB Inst_LUT4AB_ConfigMem.Inst_frame1_bit23.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame1_bit22.Q VGND VGND VPWR VPWR _0371_ sky130_fd_sc_hd__mux4_2
XANTENNA_33 net232 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_55 NN4END[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_44 N4END[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_11 net175 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_22 EE4END[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_88 net623 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_77 _0053_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_99 net2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_66 net325 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_398 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput195 net195 VGND VGND VPWR VPWR FrameData_O[16] sky130_fd_sc_hd__buf_2
Xoutput162 Inst_LUT4AB_switch_matrix.E6BEG1 VGND VGND VPWR VPWR E6BEG[11] sky130_fd_sc_hd__buf_6
Xoutput173 net173 VGND VGND VPWR VPWR EE4BEG[10] sky130_fd_sc_hd__buf_2
Xoutput184 net184 VGND VGND VPWR VPWR EE4BEG[6] sky130_fd_sc_hd__buf_2
Xoutput151 Inst_LUT4AB_switch_matrix.E2BEG7 VGND VGND VPWR VPWR E2BEG[7] sky130_fd_sc_hd__buf_8
Xoutput140 Inst_LUT4AB_switch_matrix.E1BEG0 VGND VGND VPWR VPWR E1BEG[0] sky130_fd_sc_hd__buf_8
XFILLER_47_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1030_ _0077_ _0078_ VGND VGND VPWR VPWR _0171_ sky130_fd_sc_hd__and2b_1
Xinput31 FrameData[12] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__clkbuf_2
XFILLER_61_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1863_ net787 net676 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame7_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_44_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput20 E2MID[6] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__clkbuf_2
X_1932_ net778 net683 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame5_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0814_ _0658_ _0659_ _0559_ VGND VGND VPWR VPWR _0660_ sky130_fd_sc_hd__mux2_1
XFILLER_14_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput97 S2MID[0] VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__clkbuf_2
Xinput86 S1END[1] VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__buf_2
Xinput42 FrameData[24] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__clkbuf_2
Xinput53 FrameData[9] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__buf_1
X_1794_ net799 net668 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0745_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit28.Q VGND VGND VPWR VPWR _0596_ sky130_fd_sc_hd__inv_1
Xinput64 N2END[3] VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__buf_2
Xinput75 N2MID[6] VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__buf_2
X_1228_ net661 net658 net653 net638 Inst_LUT4AB_ConfigMem.Inst_frame3_bit22.Q Inst_LUT4AB_ConfigMem.Inst_frame3_bit23.Q
+ VGND VGND VPWR VPWR _0356_ sky130_fd_sc_hd__mux4_1
X_2277_ net103 VGND VGND VPWR VPWR net310 sky130_fd_sc_hd__buf_1
X_2346_ WW4END[6] VGND VGND VPWR VPWR net385 sky130_fd_sc_hd__clkbuf_2
X_1159_ _0282_ _0291_ VGND VGND VPWR VPWR _0292_ sky130_fd_sc_hd__and2b_1
XFILLER_52_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_41_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2131_ E6END[6] VGND VGND VPWR VPWR net166 sky130_fd_sc_hd__buf_1
X_2200_ net727 VGND VGND VPWR VPWR net224 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_49_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2062_ net771 net700 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1013_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit4.Q _0155_ VGND VGND VPWR VPWR _0156_
+ sky130_fd_sc_hd__and2b_1
XFILLER_34_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1846_ net759 net676 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame7_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1915_ net750 net683 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame5_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1777_ net764 net739 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame10_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0728_ Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 VGND VGND VPWR VPWR
+ _0579_ sky130_fd_sc_hd__inv_1
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2329_ net130 VGND VGND VPWR VPWR net362 sky130_fd_sc_hd__clkbuf_2
XFILLER_27_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_243 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclone34 net663 VGND VGND VPWR VPWR net426 sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_3_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1631_ net805 net723 VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_69_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1700_ net795 net730 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame12_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1562_ net751 net713 VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3
+ sky130_fd_sc_hd__dlxtp_1
X_1493_ net766 net704 VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_69_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_316 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2045_ net810 net701 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_39_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2114_ Inst_LUT4AB_switch_matrix.E2BEG3 VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__buf_2
X_1829_ net794 net673 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame8_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_38_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0993_ _0571_ _0133_ _0136_ _0137_ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.JW2BEG5
+ sky130_fd_sc_hd__o22a_4
X_1614_ net772 net720 VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.c_I0mux
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_8_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1476_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit29.Q _0573_ _0522_ _0541_ VGND VGND VPWR
+ VPWR _0543_ sky130_fd_sc_hd__a31o_1
XFILLER_39_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1545_ net784 net709 VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5
+ sky130_fd_sc_hd__dlxtp_1
X_2028_ net778 net697 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_20_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout785 net786 VGND VGND VPWR VPWR net785 sky130_fd_sc_hd__buf_4
Xfanout752 net51 VGND VGND VPWR VPWR net752 sky130_fd_sc_hd__buf_4
XFILLER_45_135 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout796 net36 VGND VGND VPWR VPWR net796 sky130_fd_sc_hd__buf_4
Xfanout774 net776 VGND VGND VPWR VPWR net774 sky130_fd_sc_hd__buf_4
Xfanout741 net742 VGND VGND VPWR VPWR net741 sky130_fd_sc_hd__clkbuf_2
Xfanout730 net732 VGND VGND VPWR VPWR net730 sky130_fd_sc_hd__clkbuf_2
Xfanout763 net764 VGND VGND VPWR VPWR net763 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_71_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_145 net664 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_112 net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_101 net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_156 net768 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_123 net363 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_134 net788 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1261_ _0381_ _0584_ _0383_ _0385_ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.JS2BEG7
+ sky130_fd_sc_hd__o22a_1
X_1330_ net57 net113 net85 net430 Inst_LUT4AB_ConfigMem.Inst_frame11_bit21.Q Inst_LUT4AB_ConfigMem.Inst_frame11_bit20.Q
+ VGND VGND VPWR VPWR _0445_ sky130_fd_sc_hd__mux4_1
XFILLER_30_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1192_ _0323_ Inst_LH_LUT4c_frame_config_dffesr.LUT_flop Inst_LH_LUT4c_frame_config_dffesr.c_out_mux
+ VGND VGND VPWR VPWR H sky130_fd_sc_hd__mux2_4
Xinput7 E2END[1] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__dlymetal6s2s_1
X_0976_ _0119_ _0120_ _0111_ _0110_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit13.Q Inst_LUT4AB_ConfigMem.Inst_frame9_bit14.Q
+ VGND VGND VPWR VPWR _0121_ sky130_fd_sc_hd__mux4_2
Xoutput344 net344 VGND VGND VPWR VPWR UserCLKo sky130_fd_sc_hd__buf_1
Xoutput366 Inst_LUT4AB_switch_matrix.W6BEG0 VGND VGND VPWR VPWR W6BEG[10] sky130_fd_sc_hd__buf_8
Xoutput333 Inst_LUT4AB_switch_matrix.SS4BEG2 VGND VGND VPWR VPWR SS4BEG[14] sky130_fd_sc_hd__buf_8
Xoutput322 net322 VGND VGND VPWR VPWR S4BEG[4] sky130_fd_sc_hd__buf_2
Xoutput311 net311 VGND VGND VPWR VPWR S2BEGb[7] sky130_fd_sc_hd__buf_2
Xoutput300 net300 VGND VGND VPWR VPWR S2BEG[4] sky130_fd_sc_hd__buf_4
Xoutput355 net355 VGND VGND VPWR VPWR W2BEG[6] sky130_fd_sc_hd__buf_6
Xoutput377 net377 VGND VGND VPWR VPWR WW4BEG[0] sky130_fd_sc_hd__buf_2
X_1459_ _0035_ _0529_ VGND VGND VPWR VPWR _0530_ sky130_fd_sc_hd__nand2b_1
Xoutput388 net388 VGND VGND VPWR VPWR WW4BEG[5] sky130_fd_sc_hd__buf_2
X_1528_ net755 net707 VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_25_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_33_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0830_ net70 net15 net98 net126 Inst_LUT4AB_ConfigMem.Inst_frame6_bit0.Q Inst_LUT4AB_ConfigMem.Inst_frame6_bit1.Q
+ VGND VGND VPWR VPWR _0674_ sky130_fd_sc_hd__mux4_1
XFILLER_14_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0761_ net639 net629 net624 net406 Inst_LUT4AB_ConfigMem.Inst_frame3_bit6.Q Inst_LUT4AB_ConfigMem.Inst_frame3_bit7.Q
+ VGND VGND VPWR VPWR _0611_ sky130_fd_sc_hd__mux4_1
X_1244_ _0582_ _0366_ _0368_ _0370_ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.JN2BEG7
+ sky130_fd_sc_hd__o22a_1
XFILLER_56_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_39_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1313_ _0430_ VGND VGND VPWR VPWR _0431_ sky130_fd_sc_hd__inv_1
X_2293_ Inst_LUT4AB_switch_matrix.S4BEG2 VGND VGND VPWR VPWR net317 sky130_fd_sc_hd__buf_1
X_1175_ _0301_ _0302_ VGND VGND VPWR VPWR _0307_ sky130_fd_sc_hd__nand2_1
XFILLER_24_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_34 net235 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_56 NN4END[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_67 S4END[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_45 N4END[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_23 net188 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_12 net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_0959_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit16.Q _0105_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit17.Q
+ VGND VGND VPWR VPWR _0106_ sky130_fd_sc_hd__a21o_1
XANTENNA_78 _0063_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_89 net623 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput196 net196 VGND VGND VPWR VPWR FrameData_O[17] sky130_fd_sc_hd__buf_2
Xoutput174 net174 VGND VGND VPWR VPWR EE4BEG[11] sky130_fd_sc_hd__buf_2
Xoutput163 net163 VGND VGND VPWR VPWR E6BEG[1] sky130_fd_sc_hd__buf_2
Xoutput185 net185 VGND VGND VPWR VPWR EE4BEG[7] sky130_fd_sc_hd__buf_2
Xoutput152 net152 VGND VGND VPWR VPWR E2BEGb[0] sky130_fd_sc_hd__buf_2
Xoutput141 net141 VGND VGND VPWR VPWR E1BEG[1] sky130_fd_sc_hd__buf_4
XFILLER_55_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_44_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput43 FrameData[25] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__buf_1
Xinput32 FrameData[13] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__clkbuf_2
X_1862_ net791 net676 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame7_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1793_ net801 net668 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput10 E2END[4] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__buf_1
Xinput21 E2MID[7] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__clkbuf_2
X_1931_ net780 net683 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame5_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput54 FrameStrobe[10] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__clkbuf_2
X_0813_ net83 net26 net2 net814 Inst_LUT4AB_ConfigMem.Inst_frame3_bit31.Q Inst_LUT4AB_ConfigMem.Inst_frame3_bit30.Q
+ VGND VGND VPWR VPWR _0659_ sky130_fd_sc_hd__mux4_1
XFILLER_21_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput98 S2MID[1] VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__buf_2
Xinput87 S1END[2] VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__clkbuf_2
X_0744_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit16.Q VGND VGND VPWR VPWR _0595_ sky130_fd_sc_hd__inv_1
Xinput76 N2MID[7] VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__buf_2
Xinput65 N2END[4] VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__clkbuf_2
X_1227_ _0354_ _0355_ Inst_LUT4AB_ConfigMem.Inst_frame14_bit16.Q VGND VGND VPWR VPWR
+ Inst_LUT4AB_switch_matrix.M_AD sky130_fd_sc_hd__mux2_4
X_1158_ _0286_ _0290_ _0242_ VGND VGND VPWR VPWR _0291_ sky130_fd_sc_hd__mux2_1
X_2276_ net102 VGND VGND VPWR VPWR net309 sky130_fd_sc_hd__buf_1
X_2345_ WW4END[5] VGND VGND VPWR VPWR net384 sky130_fd_sc_hd__clkbuf_2
X_1089_ _0226_ _0224_ _0207_ VGND VGND VPWR VPWR _0227_ sky130_fd_sc_hd__mux2_1
XFILLER_52_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_288 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_70 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2130_ E6END[5] VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_49_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1012_ net64 net80 net3 net9 Inst_LUT4AB_ConfigMem.Inst_frame4_bit2.Q Inst_LUT4AB_ConfigMem.Inst_frame4_bit3.Q
+ VGND VGND VPWR VPWR _0155_ sky130_fd_sc_hd__mux4_1
XFILLER_19_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_263 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2061_ net774 net700 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1914_ net752 net684 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame5_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_22_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0727_ Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 VGND VGND VPWR VPWR
+ _0578_ sky130_fd_sc_hd__inv_1
X_1845_ net765 net676 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame7_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1776_ net767 net739 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame10_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_69_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2328_ net129 VGND VGND VPWR VPWR net361 sky130_fd_sc_hd__buf_1
XFILLER_25_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_9_Left_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1630_ net807 net723 VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_31_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1561_ net753 net713 VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_3_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1492_ net789 net704 VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_66_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2113_ Inst_LUT4AB_switch_matrix.E2BEG2 VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__clkbuf_2
X_2044_ net748 net699 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1828_ net796 net672 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame8_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1759_ net806 net739 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame10_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_9_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0992_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit16.Q _0134_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit17.Q
+ VGND VGND VPWR VPWR _0137_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_14_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1613_ net775 net719 VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.c_out_mux
+ sky130_fd_sc_hd__dlxtp_1
X_1544_ net785 net709 VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_8_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1475_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit29.Q _0522_ _0228_ VGND VGND VPWR VPWR
+ _0542_ sky130_fd_sc_hd__a21oi_1
XFILLER_39_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_65_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_59_Left_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2027_ net780 net697 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_50_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_68_Left_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout720 FrameStrobe[15] VGND VGND VPWR VPWR net720 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout742 net54 VGND VGND VPWR VPWR net742 sky130_fd_sc_hd__buf_2
Xfanout731 net732 VGND VGND VPWR VPWR net731 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_113 net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout797 net798 VGND VGND VPWR VPWR net797 sky130_fd_sc_hd__clkbuf_4
Xfanout786 net41 VGND VGND VPWR VPWR net786 sky130_fd_sc_hd__buf_4
XFILLER_45_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_102 net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout764 net46 VGND VGND VPWR VPWR net764 sky130_fd_sc_hd__buf_4
Xfanout775 net776 VGND VGND VPWR VPWR net775 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_28_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout753 net754 VGND VGND VPWR VPWR net753 sky130_fd_sc_hd__clkbuf_4
XANTENNA_124 net369 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_146 net786 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_135 net788 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_157 net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1191_ _0315_ _0310_ _0322_ _0311_ VGND VGND VPWR VPWR _0323_ sky130_fd_sc_hd__a22o_1
X_1260_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit24.Q _0384_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit25.Q
+ VGND VGND VPWR VPWR _0385_ sky130_fd_sc_hd__a21o_1
Xinput8 E2END[2] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__buf_2
XFILLER_24_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0975_ net72 net17 net100 net128 Inst_LUT4AB_ConfigMem.Inst_frame6_bit12.Q Inst_LUT4AB_ConfigMem.Inst_frame6_bit13.Q
+ VGND VGND VPWR VPWR _0120_ sky130_fd_sc_hd__mux4_2
Xoutput367 Inst_LUT4AB_switch_matrix.W6BEG1 VGND VGND VPWR VPWR W6BEG[11] sky130_fd_sc_hd__buf_6
X_1527_ net757 net707 VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6
+ sky130_fd_sc_hd__dlxtp_1
Xoutput334 net334 VGND VGND VPWR VPWR SS4BEG[15] sky130_fd_sc_hd__buf_6
Xoutput312 net312 VGND VGND VPWR VPWR S4BEG[0] sky130_fd_sc_hd__buf_2
Xoutput323 net323 VGND VGND VPWR VPWR S4BEG[5] sky130_fd_sc_hd__buf_2
Xoutput345 net345 VGND VGND VPWR VPWR W1BEG[0] sky130_fd_sc_hd__clkbuf_4
Xoutput301 net301 VGND VGND VPWR VPWR S2BEG[5] sky130_fd_sc_hd__buf_6
Xoutput356 Inst_LUT4AB_switch_matrix.JW2BEG7 VGND VGND VPWR VPWR W2BEG[7] sky130_fd_sc_hd__buf_6
Xoutput389 net389 VGND VGND VPWR VPWR WW4BEG[6] sky130_fd_sc_hd__buf_2
Xoutput378 net378 VGND VGND VPWR VPWR WW4BEG[10] sky130_fd_sc_hd__buf_2
X_1389_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit27.Q _0488_ _0491_ _0492_ VGND VGND
+ VPWR VPWR Inst_LUT4AB_switch_matrix.EE4BEG1 sky130_fd_sc_hd__o22a_4
X_1458_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit21.Q _0522_ VGND VGND VPWR VPWR _0529_
+ sky130_fd_sc_hd__nand2_1
XFILLER_50_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_33_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0760_ _0609_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit8.Q VGND VGND VPWR VPWR _0610_
+ sky130_fd_sc_hd__or2_4
XFILLER_14_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1174_ _0301_ _0302_ VGND VGND VPWR VPWR _0306_ sky130_fd_sc_hd__and2_1
X_1243_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit24.Q _0369_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit25.Q
+ VGND VGND VPWR VPWR _0370_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_39_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1312_ net650 net411 net646 net641 Inst_LUT4AB_ConfigMem.Inst_frame11_bit30.Q Inst_LUT4AB_ConfigMem.Inst_frame11_bit31.Q
+ VGND VGND VPWR VPWR _0430_ sky130_fd_sc_hd__mux4_1
XFILLER_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_22_Left_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_13 EE4END[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_57 NN4END[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_46 N4END[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_24 net191 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_35 Inst_LUT4AB_switch_matrix.JW2BEG6 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_0889_ net813 net92 net120 net134 Inst_LUT4AB_ConfigMem.Inst_frame3_bit2.Q Inst_LUT4AB_ConfigMem.Inst_frame3_bit3.Q
+ VGND VGND VPWR VPWR _0041_ sky130_fd_sc_hd__mux4_1
X_0958_ net87 net113 net95 net666 Inst_LUT4AB_ConfigMem.Inst_frame2_bit15.Q Inst_LUT4AB_ConfigMem.Inst_frame2_bit14.Q
+ VGND VGND VPWR VPWR _0105_ sky130_fd_sc_hd__mux4_1
XANTENNA_79 _0063_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_68 net331 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput197 net197 VGND VGND VPWR VPWR FrameData_O[18] sky130_fd_sc_hd__buf_2
Xoutput164 net164 VGND VGND VPWR VPWR E6BEG[2] sky130_fd_sc_hd__buf_2
Xoutput175 net175 VGND VGND VPWR VPWR EE4BEG[12] sky130_fd_sc_hd__buf_4
Xoutput186 net186 VGND VGND VPWR VPWR EE4BEG[8] sky130_fd_sc_hd__buf_2
Xoutput153 net153 VGND VGND VPWR VPWR E2BEGb[1] sky130_fd_sc_hd__buf_2
Xoutput142 Inst_LUT4AB_switch_matrix.E1BEG2 VGND VGND VPWR VPWR E1BEG[2] sky130_fd_sc_hd__buf_6
XFILLER_43_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_44_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1930_ net781 net685 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame5_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_36_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput88 S1END[3] VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__buf_2
Xinput44 FrameData[28] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__buf_2
Xinput33 FrameData[14] VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__clkbuf_2
X_1861_ net793 net677 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame7_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput22 E6END[0] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__dlymetal6s2s_1
X_1792_ net803 net668 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput11 E2END[5] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__clkbuf_2
Xinput66 N2END[5] VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__clkbuf_2
Xinput77 N4END[0] VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__clkbuf_2
Xinput55 FrameStrobe[19] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__clkbuf_2
X_0812_ net107 net111 net119 net133 Inst_LUT4AB_ConfigMem.Inst_frame3_bit30.Q Inst_LUT4AB_ConfigMem.Inst_frame3_bit31.Q
+ VGND VGND VPWR VPWR _0658_ sky130_fd_sc_hd__mux4_1
X_0743_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit29.Q VGND VGND VPWR VPWR _0594_ sky130_fd_sc_hd__inv_1
Xinput99 S2MID[2] VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__clkbuf_2
XFILLER_69_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2344_ WW4END[4] VGND VGND VPWR VPWR net377 sky130_fd_sc_hd__clkbuf_2
X_1226_ net623 _0354_ net412 VGND VGND VPWR VPWR _0355_ sky130_fd_sc_hd__mux2_4
X_1157_ _0287_ _0288_ _0289_ VGND VGND VPWR VPWR _0290_ sky130_fd_sc_hd__and3_1
XFILLER_37_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2275_ net101 VGND VGND VPWR VPWR net308 sky130_fd_sc_hd__clkbuf_2
X_1088_ Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 _0210_ _0214_ Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10
+ _0225_ VGND VGND VPWR VPWR _0226_ sky130_fd_sc_hd__a221o_1
XFILLER_20_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_41_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_49_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2060_ net778 net702 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1011_ net813 net92 net120 net136 Inst_LUT4AB_ConfigMem.Inst_frame4_bit2.Q Inst_LUT4AB_ConfigMem.Inst_frame4_bit3.Q
+ VGND VGND VPWR VPWR _0154_ sky130_fd_sc_hd__mux4_1
XFILLER_34_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1913_ net754 net684 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame5_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0726_ Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 VGND VGND VPWR VPWR
+ _0577_ sky130_fd_sc_hd__inv_1
X_1775_ net769 net742 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame10_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_31_Left_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1844_ net790 net675 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame7_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_57_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2327_ net128 VGND VGND VPWR VPWR net360 sky130_fd_sc_hd__clkbuf_2
XFILLER_40_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_40_Left_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2189_ FrameStrobe[2] VGND VGND VPWR VPWR net232 sky130_fd_sc_hd__clkbuf_2
X_1209_ Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 _0334_ _0336_ Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13
+ VGND VGND VPWR VPWR _0339_ sky130_fd_sc_hd__o22a_1
XFILLER_40_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_3_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1560_ net756 net712 VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_33_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2112_ Inst_LUT4AB_switch_matrix.E2BEG1 VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__buf_4
X_1491_ net811 net704 VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_52_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2043_ net750 net699 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1827_ net798 net674 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame8_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1689_ net50 net733 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame12_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0709_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit1.Q VGND VGND VPWR VPWR _0560_ sky130_fd_sc_hd__inv_1
XTAP_TAPCELL_ROW_9_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1758_ net807 net739 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame10_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_54_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0991_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit16.Q _0135_ VGND VGND VPWR VPWR _0136_
+ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_14_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1474_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit20.Q net621 VGND VGND VPWR VPWR _0541_
+ sky130_fd_sc_hd__and2_1
X_1612_ net777 net720 VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15
+ sky130_fd_sc_hd__dlxtp_1
X_1543_ net787 net709 VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_5_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2026_ net781 net697 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_50_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout721 net725 VGND VGND VPWR VPWR net721 sky130_fd_sc_hd__buf_2
Xfanout754 net50 VGND VGND VPWR VPWR net754 sky130_fd_sc_hd__buf_4
Xfanout765 net766 VGND VGND VPWR VPWR net765 sky130_fd_sc_hd__clkbuf_4
Xfanout776 FrameData[26] VGND VGND VPWR VPWR net776 sky130_fd_sc_hd__clkbuf_4
Xfanout710 net711 VGND VGND VPWR VPWR net710 sky130_fd_sc_hd__clkbuf_1
Xfanout732 net734 VGND VGND VPWR VPWR net732 sky130_fd_sc_hd__clkbuf_2
Xfanout743 net745 VGND VGND VPWR VPWR net743 sky130_fd_sc_hd__buf_2
Xfanout787 net788 VGND VGND VPWR VPWR net787 sky130_fd_sc_hd__clkbuf_4
XANTENNA_147 net787 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_136 net804 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout798 net35 VGND VGND VPWR VPWR net798 sky130_fd_sc_hd__buf_4
XANTENNA_158 net147 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_103 net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_114 net136 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_125 net371 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_310 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1190_ _0318_ _0321_ _0300_ VGND VGND VPWR VPWR _0322_ sky130_fd_sc_hd__mux2_1
Xinput9 E2END[3] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_2
XFILLER_44_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0974_ net71 net99 net16 Inst_LUT4AB_switch_matrix.E2BEG5 Inst_LUT4AB_ConfigMem.Inst_frame7_bit13.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame7_bit12.Q VGND VGND VPWR VPWR _0119_ sky130_fd_sc_hd__mux4_2
XFILLER_32_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput302 net302 VGND VGND VPWR VPWR S2BEG[6] sky130_fd_sc_hd__buf_4
Xoutput346 Inst_LUT4AB_switch_matrix.W1BEG1 VGND VGND VPWR VPWR W1BEG[1] sky130_fd_sc_hd__buf_8
Xoutput335 net335 VGND VGND VPWR VPWR SS4BEG[1] sky130_fd_sc_hd__buf_2
Xoutput313 net313 VGND VGND VPWR VPWR S4BEG[10] sky130_fd_sc_hd__buf_2
Xoutput324 net324 VGND VGND VPWR VPWR S4BEG[6] sky130_fd_sc_hd__buf_2
X_1457_ net480 _0528_ _0527_ VGND VGND VPWR VPWR _0001_ sky130_fd_sc_hd__mux2_1
Xoutput357 net357 VGND VGND VPWR VPWR W2BEGb[0] sky130_fd_sc_hd__buf_2
Xoutput368 net368 VGND VGND VPWR VPWR W6BEG[1] sky130_fd_sc_hd__buf_2
Xoutput379 net379 VGND VGND VPWR VPWR WW4BEG[11] sky130_fd_sc_hd__buf_2
X_1526_ net760 net707 VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5
+ sky130_fd_sc_hd__dlxtp_1
X_1388_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit26.Q _0489_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit27.Q
+ VGND VGND VPWR VPWR _0492_ sky130_fd_sc_hd__a21bo_1
XFILLER_35_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_310 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2009_ net754 net696 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_2_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1311_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit0.Q _0428_ VGND VGND VPWR VPWR _0429_
+ sky130_fd_sc_hd__or2_1
X_2291_ Inst_LUT4AB_switch_matrix.S4BEG0 VGND VGND VPWR VPWR net315 sky130_fd_sc_hd__clkbuf_2
X_1173_ Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 _0303_ _0304_ Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0
+ VGND VGND VPWR VPWR _0305_ sky130_fd_sc_hd__o22a_1
XFILLER_64_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1242_ net85 net113 net89 net666 Inst_LUT4AB_ConfigMem.Inst_frame4_bit23.Q Inst_LUT4AB_ConfigMem.Inst_frame4_bit22.Q
+ VGND VGND VPWR VPWR _0369_ sky130_fd_sc_hd__mux4_1
XFILLER_52_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_36 net257 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_47 N4END[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_25 net202 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_14 EE4END[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_58 NN4END[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_0888_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit4.Q _0039_ VGND VGND VPWR VPWR _0040_
+ sky130_fd_sc_hd__and2b_1
X_0957_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit16.Q _0103_ VGND VGND VPWR VPWR _0104_
+ sky130_fd_sc_hd__and2b_1
Xoutput143 Inst_LUT4AB_switch_matrix.E1BEG3 VGND VGND VPWR VPWR E1BEG[3] sky130_fd_sc_hd__buf_8
XANTENNA_69 net359 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput198 net198 VGND VGND VPWR VPWR FrameData_O[19] sky130_fd_sc_hd__buf_2
Xoutput165 net165 VGND VGND VPWR VPWR E6BEG[3] sky130_fd_sc_hd__buf_2
Xoutput176 Inst_LUT4AB_switch_matrix.EE4BEG1 VGND VGND VPWR VPWR EE4BEG[13] sky130_fd_sc_hd__buf_8
Xoutput187 net187 VGND VGND VPWR VPWR EE4BEG[9] sky130_fd_sc_hd__buf_2
Xoutput154 net154 VGND VGND VPWR VPWR E2BEGb[2] sky130_fd_sc_hd__buf_2
X_1509_ net793 net705 VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_23_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_44_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1860_ net795 net675 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame7_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_14_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput89 S2END[0] VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__buf_2
Xinput45 FrameData[29] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__clkbuf_2
Xinput34 FrameData[15] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__clkbuf_2
Xinput23 E6END[1] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__clkbuf_2
X_1791_ net805 net667 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput12 E2END[6] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__clkbuf_2
X_0811_ _0559_ _0656_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit1.Q VGND VGND VPWR VPWR
+ _0657_ sky130_fd_sc_hd__o21a_1
Xinput56 FrameStrobe[4] VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__buf_2
Xinput67 N2END[6] VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__buf_2
Xinput78 N4END[1] VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0742_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit28.Q VGND VGND VPWR VPWR _0593_ sky130_fd_sc_hd__inv_2
XFILLER_69_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2274_ net100 VGND VGND VPWR VPWR net307 sky130_fd_sc_hd__clkbuf_1
X_1225_ net652 net636 _0353_ VGND VGND VPWR VPWR _0354_ sky130_fd_sc_hd__mux2_4
X_1156_ Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 _0267_ _0268_ Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7
+ VGND VGND VPWR VPWR _0289_ sky130_fd_sc_hd__o22a_1
X_1087_ Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 _0212_ _0213_ Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12
+ VGND VGND VPWR VPWR _0225_ sky130_fd_sc_hd__a22o_1
XFILLER_37_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_35_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1989_ net794 net692 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_57_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_41_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_49_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1010_ _0151_ _0152_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit4.Q VGND VGND VPWR VPWR
+ _0153_ sky130_fd_sc_hd__mux2_4
XFILLER_14_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1843_ net812 net675 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame7_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1912_ net755 net684 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame5_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0725_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit21.Q VGND VGND VPWR VPWR _0576_ sky130_fd_sc_hd__inv_1
X_1774_ net771 net54 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame10_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2257_ Inst_LUT4AB_switch_matrix.NN4BEG2 VGND VGND VPWR VPWR net281 sky130_fd_sc_hd__clkbuf_1
X_1208_ _0191_ _0192_ _0183_ _0182_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit7.Q Inst_LUT4AB_ConfigMem.Inst_frame9_bit8.Q
+ VGND VGND VPWR VPWR _0338_ sky130_fd_sc_hd__mux4_2
X_2326_ net127 VGND VGND VPWR VPWR net359 sky130_fd_sc_hd__clkbuf_2
X_1139_ net646 net627 net642 net622 Inst_LUT4AB_ConfigMem.Inst_frame1_bit19.Q Inst_LUT4AB_ConfigMem.Inst_frame1_bit18.Q
+ VGND VGND VPWR VPWR _0273_ sky130_fd_sc_hd__mux4_1
XFILLER_65_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2188_ FrameStrobe[1] VGND VGND VPWR VPWR net231 sky130_fd_sc_hd__clkbuf_2
XFILLER_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1490_ net761 net55 VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_66_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2042_ net752 net699 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2111_ Inst_LUT4AB_switch_matrix.E2BEG0 VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__buf_4
XFILLER_47_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_227 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1826_ net799 net674 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame8_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1688_ net756 net733 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame12_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_39_Right_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0708_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit0.Q VGND VGND VPWR VPWR _0559_ sky130_fd_sc_hd__inv_2
X_1757_ net809 net739 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame10_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_68_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_48_Right_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_57_Right_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_66_Right_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1611_ net779 net718 VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14
+ sky130_fd_sc_hd__dlxtp_1
X_0990_ net59 net67 net816 net12 Inst_LUT4AB_ConfigMem.Inst_frame1_bit14.Q Inst_LUT4AB_ConfigMem.Inst_frame1_bit15.Q
+ VGND VGND VPWR VPWR _0135_ sky130_fd_sc_hd__mux4_1
XFILLER_8_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_14_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1473_ _0539_ _0540_ net483 _0538_ VGND VGND VPWR VPWR _0005_ sky130_fd_sc_hd__a2bb2o_1
X_1542_ net791 net709 VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_65_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2025_ net783 net697 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_39_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1809_ net764 net669 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_2_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout722 net725 VGND VGND VPWR VPWR net722 sky130_fd_sc_hd__clkbuf_2
Xfanout777 net778 VGND VGND VPWR VPWR net777 sky130_fd_sc_hd__clkbuf_4
Xfanout788 net40 VGND VGND VPWR VPWR net788 sky130_fd_sc_hd__buf_4
Xfanout733 net734 VGND VGND VPWR VPWR net733 sky130_fd_sc_hd__buf_2
Xfanout755 net756 VGND VGND VPWR VPWR net755 sky130_fd_sc_hd__clkbuf_4
Xfanout700 FrameStrobe[1] VGND VGND VPWR VPWR net700 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout766 FrameData[2] VGND VGND VPWR VPWR net766 sky130_fd_sc_hd__buf_4
Xfanout711 FrameStrobe[17] VGND VGND VPWR VPWR net711 sky130_fd_sc_hd__buf_1
Xfanout744 net745 VGND VGND VPWR VPWR net744 sky130_fd_sc_hd__clkbuf_2
Xfanout799 net800 VGND VGND VPWR VPWR net799 sky130_fd_sc_hd__clkbuf_4
XANTENNA_104 net44 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_115 net397 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_148 net2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_137 net809 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_126 net389 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0973_ _0114_ _0569_ _0116_ _0118_ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.E2BEG5
+ sky130_fd_sc_hd__o22a_4
Xoutput314 net314 VGND VGND VPWR VPWR S4BEG[11] sky130_fd_sc_hd__buf_2
Xoutput325 net325 VGND VGND VPWR VPWR S4BEG[7] sky130_fd_sc_hd__buf_2
Xoutput303 net303 VGND VGND VPWR VPWR S2BEG[7] sky130_fd_sc_hd__buf_8
X_1387_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit26.Q _0490_ VGND VGND VPWR VPWR _0491_
+ sky130_fd_sc_hd__and2b_1
X_1525_ net766 net708 VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4
+ sky130_fd_sc_hd__dlxtp_1
Xoutput347 Inst_LUT4AB_switch_matrix.W1BEG2 VGND VGND VPWR VPWR W1BEG[2] sky130_fd_sc_hd__buf_6
Xoutput336 net336 VGND VGND VPWR VPWR SS4BEG[2] sky130_fd_sc_hd__buf_2
X_1456_ Inst_LA_LUT4c_frame_config_dffesr.c_reset_value _0696_ _0526_ VGND VGND VPWR
+ VPWR _0528_ sky130_fd_sc_hd__mux2_1
Xoutput358 net358 VGND VGND VPWR VPWR W2BEGb[1] sky130_fd_sc_hd__buf_2
Xoutput369 net369 VGND VGND VPWR VPWR W6BEG[2] sky130_fd_sc_hd__buf_2
X_2008_ net755 net696 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_23_322 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2290_ S4END[15] VGND VGND VPWR VPWR net314 sky130_fd_sc_hd__clkbuf_2
X_1241_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit24.Q _0367_ VGND VGND VPWR VPWR _0368_
+ sky130_fd_sc_hd__and2b_1
XFILLER_44_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1310_ net4 net666 net660 net430 Inst_LUT4AB_ConfigMem.Inst_frame11_bit30.Q Inst_LUT4AB_ConfigMem.Inst_frame11_bit31.Q
+ VGND VGND VPWR VPWR _0428_ sky130_fd_sc_hd__mux4_1
X_1172_ _0301_ _0302_ VGND VGND VPWR VPWR _0304_ sky130_fd_sc_hd__or2_4
XFILLER_64_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_119 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_59 NN4END[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_48 NN4END[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_37 N4END[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_26 net213 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_0956_ net59 net67 net816 net12 Inst_LUT4AB_ConfigMem.Inst_frame2_bit14.Q Inst_LUT4AB_ConfigMem.Inst_frame2_bit15.Q
+ VGND VGND VPWR VPWR _0103_ sky130_fd_sc_hd__mux4_1
XFILLER_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_15 EE4END[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_22_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput166 net166 VGND VGND VPWR VPWR E6BEG[4] sky130_fd_sc_hd__buf_2
Xoutput177 net177 VGND VGND VPWR VPWR EE4BEG[14] sky130_fd_sc_hd__buf_4
X_0887_ net58 net80 net64 net9 Inst_LUT4AB_ConfigMem.Inst_frame3_bit3.Q Inst_LUT4AB_ConfigMem.Inst_frame3_bit2.Q
+ VGND VGND VPWR VPWR _0039_ sky130_fd_sc_hd__mux4_1
Xoutput155 net155 VGND VGND VPWR VPWR E2BEGb[3] sky130_fd_sc_hd__buf_2
Xoutput144 net144 VGND VGND VPWR VPWR E2BEG[0] sky130_fd_sc_hd__buf_6
Xoutput199 net199 VGND VGND VPWR VPWR FrameData_O[1] sky130_fd_sc_hd__buf_2
Xoutput188 net188 VGND VGND VPWR VPWR FrameData_O[0] sky130_fd_sc_hd__buf_2
X_1508_ net796 net703 VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6
+ sky130_fd_sc_hd__dlxtp_1
X_1439_ _0510_ _0511_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit30.Q VGND VGND VPWR VPWR
+ _0512_ sky130_fd_sc_hd__mux2_1
XFILLER_62_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1790_ net807 net667 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_44_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput13 E2END[7] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__clkbuf_2
X_0810_ net639 net629 net624 net622 Inst_LUT4AB_ConfigMem.Inst_frame3_bit30.Q Inst_LUT4AB_ConfigMem.Inst_frame3_bit31.Q
+ VGND VGND VPWR VPWR _0656_ sky130_fd_sc_hd__mux4_1
Xinput46 FrameData[30] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__buf_2
Xinput35 FrameData[16] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__clkbuf_2
Xinput24 EE4END[0] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__clkbuf_2
Xinput57 N1END[0] VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__clkbuf_4
Xinput79 N4END[2] VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__clkbuf_2
Xinput68 N2END[7] VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__buf_2
X_0741_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit29.Q VGND VGND VPWR VPWR _0592_ sky130_fd_sc_hd__inv_1
X_1224_ _0352_ net396 Inst_LUT4AB_ConfigMem.Inst_frame14_bit16.Q VGND VGND VPWR VPWR
+ _0353_ sky130_fd_sc_hd__mux2_4
X_2273_ net99 VGND VGND VPWR VPWR net306 sky130_fd_sc_hd__buf_1
X_1155_ Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 _0266_ _0254_ VGND
+ VGND VPWR VPWR _0288_ sky130_fd_sc_hd__or3b_1
X_1086_ Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 _0210_ _0212_ Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15
+ _0223_ VGND VGND VPWR VPWR _0224_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_35_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1988_ net795 net692 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0939_ _0086_ _0085_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit16.Q VGND VGND VPWR VPWR
+ _0087_ sky130_fd_sc_hd__mux2_2
XFILLER_43_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_41_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1773_ net774 net742 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame10_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1842_ net761 net674 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame8_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1911_ net757 net684 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame5_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0724_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit21.Q VGND VGND VPWR VPWR _0575_ sky130_fd_sc_hd__inv_1
XFILLER_72_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1207_ Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 _0075_ _0336_ Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12
+ _0335_ VGND VGND VPWR VPWR _0337_ sky130_fd_sc_hd__o221a_1
X_2187_ net746 VGND VGND VPWR VPWR net220 sky130_fd_sc_hd__clkbuf_2
XFILLER_25_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2325_ net126 VGND VGND VPWR VPWR net358 sky130_fd_sc_hd__clkbuf_2
X_1069_ Inst_LF_LUT4c_frame_config_dffesr.c_I0mux _0206_ _0205_ VGND VGND VPWR VPWR
+ _0207_ sky130_fd_sc_hd__o21a_1
XFILLER_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1138_ net62 net90 net27 net118 Inst_LUT4AB_ConfigMem.Inst_frame5_bit25.Q Inst_LUT4AB_ConfigMem.Inst_frame5_bit24.Q
+ VGND VGND VPWR VPWR _0272_ sky130_fd_sc_hd__mux4_2
Xclone38 net655 VGND VGND VPWR VPWR net430 sky130_fd_sc_hd__clkbuf_1
XFILLER_68_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2041_ net754 net699 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_17_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1825_ net801 net672 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame8_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_60_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0707_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit9.Q VGND VGND VPWR VPWR _0558_ sky130_fd_sc_hd__inv_1
X_1756_ net747 net739 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame10_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1687_ net758 net733 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame12_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_68_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2239_ Inst_LUT4AB_switch_matrix.N4BEG0 VGND VGND VPWR VPWR net263 sky130_fd_sc_hd__buf_4
XFILLER_21_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1610_ net782 net718 VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_14_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1472_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit19.Q _0572_ _0522_ _0538_ VGND VGND VPWR
+ VPWR _0540_ sky130_fd_sc_hd__a31o_1
X_1541_ net793 net709 VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_5_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2024_ net786 net698 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_65_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_28_Left_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1808_ net45 net668 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_49_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1739_ net780 net735 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame11_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
Xfanout723 net724 VGND VGND VPWR VPWR net723 sky130_fd_sc_hd__clkbuf_2
Xfanout778 net43 VGND VGND VPWR VPWR net778 sky130_fd_sc_hd__buf_4
Xfanout756 net49 VGND VGND VPWR VPWR net756 sky130_fd_sc_hd__clkbuf_4
Xfanout701 net702 VGND VGND VPWR VPWR net701 sky130_fd_sc_hd__clkbuf_2
Xfanout712 net714 VGND VGND VPWR VPWR net712 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_37_Left_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout745 net746 VGND VGND VPWR VPWR net745 sky130_fd_sc_hd__clkbuf_2
Xfanout734 FrameStrobe[12] VGND VGND VPWR VPWR net734 sky130_fd_sc_hd__clkbuf_2
Xfanout767 net768 VGND VGND VPWR VPWR net767 sky130_fd_sc_hd__clkbuf_4
Xfanout789 net790 VGND VGND VPWR VPWR net789 sky130_fd_sc_hd__buf_4
XFILLER_18_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_149 net57 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_116 net397 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_127 net753 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_46_Left_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_105 net48 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_138 net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_235 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0972_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit16.Q _0117_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit17.Q
+ VGND VGND VPWR VPWR _0118_ sky130_fd_sc_hd__a21o_1
XFILLER_32_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput348 Inst_LUT4AB_switch_matrix.W1BEG3 VGND VGND VPWR VPWR W1BEG[3] sky130_fd_sc_hd__buf_8
Xoutput337 net337 VGND VGND VPWR VPWR SS4BEG[3] sky130_fd_sc_hd__buf_2
Xoutput315 net315 VGND VGND VPWR VPWR S4BEG[12] sky130_fd_sc_hd__buf_4
Xoutput326 net326 VGND VGND VPWR VPWR S4BEG[8] sky130_fd_sc_hd__buf_2
Xoutput304 net304 VGND VGND VPWR VPWR S2BEGb[0] sky130_fd_sc_hd__buf_2
Xoutput359 net359 VGND VGND VPWR VPWR W2BEGb[2] sky130_fd_sc_hd__buf_2
X_1524_ net789 net707 VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3
+ sky130_fd_sc_hd__dlxtp_1
X_1386_ net410 _0652_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit25.Q VGND VGND VPWR VPWR
+ _0490_ sky130_fd_sc_hd__mux2_1
X_1455_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit2.Q net467 VGND VGND VPWR VPWR _0527_
+ sky130_fd_sc_hd__nand2_1
X_2007_ net757 net696 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_23_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1171_ _0302_ _0301_ VGND VGND VPWR VPWR _0303_ sky130_fd_sc_hd__nand2b_1
X_1240_ net57 net61 net2 net24 Inst_LUT4AB_ConfigMem.Inst_frame4_bit22.Q Inst_LUT4AB_ConfigMem.Inst_frame4_bit23.Q
+ VGND VGND VPWR VPWR _0367_ sky130_fd_sc_hd__mux4_1
XFILLER_2_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_47_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_16 EE4END[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_49 NN4END[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_38 N4END[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_27 net217 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_0886_ _0036_ _0037_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit4.Q VGND VGND VPWR VPWR
+ _0038_ sky130_fd_sc_hd__mux2_4
X_0955_ _0100_ _0101_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit16.Q VGND VGND VPWR VPWR
+ _0102_ sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_30_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput189 net189 VGND VGND VPWR VPWR FrameData_O[10] sky130_fd_sc_hd__buf_2
Xoutput167 net167 VGND VGND VPWR VPWR E6BEG[5] sky130_fd_sc_hd__buf_2
Xoutput178 Inst_LUT4AB_switch_matrix.EE4BEG3 VGND VGND VPWR VPWR EE4BEG[15] sky130_fd_sc_hd__buf_6
Xoutput156 net156 VGND VGND VPWR VPWR E2BEGb[4] sky130_fd_sc_hd__buf_2
Xoutput145 net145 VGND VGND VPWR VPWR E2BEG[1] sky130_fd_sc_hd__buf_4
X_1507_ net798 net703 VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5
+ sky130_fd_sc_hd__dlxtp_1
X_1369_ net647 net642 Inst_LUT4AB_ConfigMem.Inst_frame12_bit2.Q VGND VGND VPWR VPWR
+ _0476_ sky130_fd_sc_hd__mux2_1
XFILLER_55_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1438_ Inst_LUT4AB_switch_matrix.JS2BEG2 Inst_LUT4AB_switch_matrix.JW2BEG2 Inst_LUT4AB_ConfigMem.Inst_frame0_bit29.Q
+ VGND VGND VPWR VPWR _0511_ sky130_fd_sc_hd__mux2_1
XFILLER_11_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput36 FrameData[17] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_44_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput25 EE4END[1] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput14 E2MID[0] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__buf_1
X_0740_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit28.Q VGND VGND VPWR VPWR _0591_ sky130_fd_sc_hd__inv_2
XFILLER_14_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput47 FrameData[31] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__clkbuf_2
X_2341_ W6END[11] VGND VGND VPWR VPWR net376 sky130_fd_sc_hd__buf_4
Xinput58 N1END[1] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__clkbuf_4
Xinput69 N2MID[0] VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1154_ Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 _0254_ _0266_ VGND
+ VGND VPWR VPWR _0287_ sky130_fd_sc_hd__or3b_4
X_1223_ _0350_ _0351_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit21.Q VGND VGND VPWR VPWR
+ _0352_ sky130_fd_sc_hd__mux2_4
X_2272_ net98 VGND VGND VPWR VPWR net305 sky130_fd_sc_hd__clkbuf_1
X_1085_ Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 _0213_ _0214_ Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11
+ VGND VGND VPWR VPWR _0223_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_35_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1987_ net797 net692 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0938_ net662 net656 net653 net636 Inst_LUT4AB_ConfigMem.Inst_frame4_bit14.Q Inst_LUT4AB_ConfigMem.Inst_frame4_bit15.Q
+ VGND VGND VPWR VPWR _0086_ sky130_fd_sc_hd__mux4_1
X_0869_ _0016_ _0017_ VGND VGND VPWR VPWR _0022_ sky130_fd_sc_hd__nand2_1
XFILLER_51_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_57_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1910_ net759 net686 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame5_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_34_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0723_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit21.Q VGND VGND VPWR VPWR _0574_ sky130_fd_sc_hd__inv_1
X_1772_ net777 net742 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame10_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1841_ net763 net674 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame8_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2324_ net125 VGND VGND VPWR VPWR net357 sky130_fd_sc_hd__buf_1
XFILLER_69_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2255_ Inst_LUT4AB_switch_matrix.NN4BEG0 VGND VGND VPWR VPWR net279 sky130_fd_sc_hd__buf_1
X_1206_ _0054_ _0073_ VGND VGND VPWR VPWR _0336_ sky130_fd_sc_hd__nand2b_1
X_1137_ net81 net117 net22 Inst_LUT4AB_switch_matrix.JW2BEG4 Inst_LUT4AB_ConfigMem.Inst_frame0_bit25.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame0_bit24.Q VGND VGND VPWR VPWR _0271_ sky130_fd_sc_hd__mux4_2
X_2186_ net762 VGND VGND VPWR VPWR net212 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_63_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1068_ _0092_ _0093_ _0095_ _0094_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit21.Q Inst_LUT4AB_ConfigMem.Inst_frame9_bit22.Q
+ VGND VGND VPWR VPWR _0206_ sky130_fd_sc_hd__mux4_1
XFILLER_47_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2040_ net755 net700 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_62_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_17_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1686_ net760 net733 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame12_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1824_ net804 net672 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame8_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1755_ net749 net741 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame10_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0706_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit8.Q VGND VGND VPWR VPWR _0557_ sky130_fd_sc_hd__inv_1
X_2238_ N4END[15] VGND VGND VPWR VPWR net262 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_68_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2307_ Inst_LUT4AB_switch_matrix.SS4BEG0 VGND VGND VPWR VPWR net331 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_13_Left_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2169_ net801 VGND VGND VPWR VPWR net193 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_0_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1540_ net796 net709 VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0
+ sky130_fd_sc_hd__dlxtp_1
X_1471_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit19.Q _0522_ _0150_ VGND VGND VPWR VPWR
+ _0539_ sky130_fd_sc_hd__a21oi_1
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2023_ net788 net698 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_65_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1807_ net770 net667 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
Xfanout724 net725 VGND VGND VPWR VPWR net724 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout713 net714 VGND VGND VPWR VPWR net713 sky130_fd_sc_hd__buf_1
Xfanout702 FrameStrobe[1] VGND VGND VPWR VPWR net702 sky130_fd_sc_hd__clkbuf_2
X_1738_ net781 net736 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame11_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1669_ net793 net728 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame13_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
Xfanout779 net780 VGND VGND VPWR VPWR net779 sky130_fd_sc_hd__buf_4
XANTENNA_106 net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout768 net45 VGND VGND VPWR VPWR net768 sky130_fd_sc_hd__buf_4
Xfanout757 FrameData[4] VGND VGND VPWR VPWR net757 sky130_fd_sc_hd__clkbuf_4
Xfanout746 FrameStrobe[0] VGND VGND VPWR VPWR net746 sky130_fd_sc_hd__clkbuf_2
Xfanout735 net736 VGND VGND VPWR VPWR net735 sky130_fd_sc_hd__clkbuf_2
XANTENNA_117 net170 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_128 net754 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_139 net89 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_70_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0971_ net85 net87 net95 net666 Inst_LUT4AB_ConfigMem.Inst_frame3_bit14.Q Inst_LUT4AB_ConfigMem.Inst_frame3_bit15.Q
+ VGND VGND VPWR VPWR _0117_ sky130_fd_sc_hd__mux4_1
XFILLER_44_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1523_ net811 net708 VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2
+ sky130_fd_sc_hd__dlxtp_1
Xoutput338 net338 VGND VGND VPWR VPWR SS4BEG[4] sky130_fd_sc_hd__buf_2
Xoutput327 net327 VGND VGND VPWR VPWR S4BEG[9] sky130_fd_sc_hd__buf_2
Xoutput316 Inst_LUT4AB_switch_matrix.S4BEG1 VGND VGND VPWR VPWR S4BEG[13] sky130_fd_sc_hd__buf_4
Xoutput305 net305 VGND VGND VPWR VPWR S2BEGb[1] sky130_fd_sc_hd__buf_2
Xoutput349 net349 VGND VGND VPWR VPWR W2BEG[0] sky130_fd_sc_hd__buf_4
X_1454_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit11.Q _0522_ VGND VGND VPWR VPWR _0526_
+ sky130_fd_sc_hd__nand2_1
XFILLER_67_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1385_ _0071_ _0095_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit25.Q VGND VGND VPWR VPWR
+ _0489_ sky130_fd_sc_hd__mux2_4
X_2006_ net759 net696 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_16_Left_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1170_ _0264_ _0265_ _0256_ _0255_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit11.Q Inst_LUT4AB_ConfigMem.Inst_frame8_bit12.Q
+ VGND VGND VPWR VPWR _0302_ sky130_fd_sc_hd__mux4_2
XFILLER_64_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_140 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_17 EE4END[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_28 FrameStrobe[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_39 N4END[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_65_Left_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0885_ net642 net633 H net405 Inst_LUT4AB_ConfigMem.Inst_frame3_bit2.Q Inst_LUT4AB_ConfigMem.Inst_frame3_bit3.Q
+ VGND VGND VPWR VPWR _0037_ sky130_fd_sc_hd__mux4_1
X_0954_ net646 net631 net627 net622 Inst_LUT4AB_ConfigMem.Inst_frame2_bit14.Q Inst_LUT4AB_ConfigMem.Inst_frame2_bit15.Q
+ VGND VGND VPWR VPWR _0101_ sky130_fd_sc_hd__mux4_2
XFILLER_32_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_30_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput168 net168 VGND VGND VPWR VPWR E6BEG[6] sky130_fd_sc_hd__buf_2
Xoutput179 net179 VGND VGND VPWR VPWR EE4BEG[1] sky130_fd_sc_hd__buf_2
Xoutput157 net157 VGND VGND VPWR VPWR E2BEGb[5] sky130_fd_sc_hd__buf_2
Xoutput146 net146 VGND VGND VPWR VPWR E2BEG[2] sky130_fd_sc_hd__buf_6
X_1506_ net799 net705 VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4
+ sky130_fd_sc_hd__dlxtp_1
X_1437_ Inst_LUT4AB_switch_matrix.JN2BEG2 Inst_LUT4AB_switch_matrix.E2BEG2 Inst_LUT4AB_ConfigMem.Inst_frame0_bit29.Q
+ VGND VGND VPWR VPWR _0510_ sky130_fd_sc_hd__mux2_1
X_1368_ net815 net665 net661 net658 Inst_LUT4AB_ConfigMem.Inst_frame12_bit2.Q Inst_LUT4AB_ConfigMem.Inst_frame12_bit3.Q
+ VGND VGND VPWR VPWR _0475_ sky130_fd_sc_hd__mux4_1
XFILLER_70_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1299_ net654 net634 net649 net645 Inst_LUT4AB_ConfigMem.Inst_frame5_bit27.Q Inst_LUT4AB_ConfigMem.Inst_frame5_bit26.Q
+ VGND VGND VPWR VPWR _0418_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_44_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_1_Left_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput37 FrameData[18] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__buf_1
Xinput48 FrameData[3] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_52_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput26 EE4END[2] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__clkbuf_2
Xinput15 E2MID[1] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__buf_2
Xinput59 N1END[2] VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__buf_4
XFILLER_10_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2340_ W6END[10] VGND VGND VPWR VPWR net375 sky130_fd_sc_hd__buf_4
X_2271_ net97 VGND VGND VPWR VPWR net304 sky130_fd_sc_hd__buf_1
X_1153_ Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2
+ Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6
+ _0266_ _0254_ VGND VGND VPWR VPWR _0286_ sky130_fd_sc_hd__mux4_1
X_1084_ _0221_ _0217_ _0207_ VGND VGND VPWR VPWR _0222_ sky130_fd_sc_hd__mux2_4
X_1222_ Inst_LUT4AB_switch_matrix.JS2BEG5 Inst_LUT4AB_switch_matrix.JW2BEG5 Inst_LUT4AB_ConfigMem.Inst_frame8_bit20.Q
+ VGND VGND VPWR VPWR _0351_ sky130_fd_sc_hd__mux2_4
XFILLER_37_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1986_ net800 net692 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0937_ net646 net631 net627 net397 Inst_LUT4AB_ConfigMem.Inst_frame4_bit14.Q Inst_LUT4AB_ConfigMem.Inst_frame4_bit15.Q
+ VGND VGND VPWR VPWR _0085_ sky130_fd_sc_hd__mux4_1
X_0868_ _0016_ _0017_ VGND VGND VPWR VPWR _0021_ sky130_fd_sc_hd__and2_4
X_0799_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit8.Q _0645_ VGND VGND VPWR VPWR _0646_
+ sky130_fd_sc_hd__or2_4
XFILLER_51_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1840_ net767 net674 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame8_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0722_ Inst_LF_LUT4c_frame_config_dffesr.c_reset_value VGND VGND VPWR VPWR _0573_
+ sky130_fd_sc_hd__inv_1
X_1771_ net779 net742 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame10_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_8_66 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2254_ NN4END[15] VGND VGND VPWR VPWR net278 sky130_fd_sc_hd__buf_1
X_2185_ net764 VGND VGND VPWR VPWR net211 sky130_fd_sc_hd__buf_1
X_1136_ _0577_ _0578_ _0579_ _0580_ _0266_ _0254_ VGND VGND VPWR VPWR _0270_ sky130_fd_sc_hd__mux4_1
X_1067_ _0204_ _0126_ Inst_LF_LUT4c_frame_config_dffesr.c_I0mux VGND VGND VPWR VPWR
+ _0205_ sky130_fd_sc_hd__a21bo_1
X_1205_ Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 _0074_ _0334_ Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10
+ VGND VGND VPWR VPWR _0335_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_63_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclone18 H VGND VGND VPWR VPWR net410 sky130_fd_sc_hd__buf_6
XFILLER_33_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1969_ net763 net687 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_60_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1823_ net806 net671 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame8_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_15_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1685_ net765 net733 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame12_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1754_ net751 net741 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame10_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0705_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit1.Q VGND VGND VPWR VPWR _0556_ sky130_fd_sc_hd__inv_1
X_2306_ SS4END[15] VGND VGND VPWR VPWR net330 sky130_fd_sc_hd__clkbuf_2
X_2237_ N4END[14] VGND VGND VPWR VPWR net261 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_68_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2099_ clknet_1_1__leaf_UserCLK_regs _0000_ VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.LUT_flop
+ sky130_fd_sc_hd__dfxtp_1
X_2168_ net803 VGND VGND VPWR VPWR net192 sky130_fd_sc_hd__buf_1
X_1119_ _0252_ _0253_ _0244_ _0243_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit3.Q Inst_LUT4AB_ConfigMem.Inst_frame8_bit4.Q
+ VGND VGND VPWR VPWR _0254_ sky130_fd_sc_hd__mux4_2
XFILLER_54_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_51_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_35_Right_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1470_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit10.Q _0513_ VGND VGND VPWR VPWR _0538_
+ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_44_Right_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_73_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2022_ net792 net698 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_65_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_53_Right_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1806_ net772 net667 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
Xfanout725 FrameStrobe[14] VGND VGND VPWR VPWR net725 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_62_Right_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1599_ net31 net718 VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2
+ sky130_fd_sc_hd__dlxtp_1
Xfanout714 net715 VGND VGND VPWR VPWR net714 sky130_fd_sc_hd__buf_1
Xfanout758 FrameData[4] VGND VGND VPWR VPWR net758 sky130_fd_sc_hd__clkbuf_4
Xfanout736 net737 VGND VGND VPWR VPWR net736 sky130_fd_sc_hd__dlymetal6s2s_1
X_1737_ net783 net735 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame11_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
Xfanout703 net704 VGND VGND VPWR VPWR net703 sky130_fd_sc_hd__clkbuf_2
Xfanout747 net748 VGND VGND VPWR VPWR net747 sky130_fd_sc_hd__clkbuf_4
X_1668_ net795 net728 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame13_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
XANTENNA_129 net768 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_118 EE4END[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout769 net770 VGND VGND VPWR VPWR net769 sky130_fd_sc_hd__buf_4
XANTENNA_107 net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_71_Right_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_27_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_70_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0970_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit16.Q _0115_ VGND VGND VPWR VPWR _0116_
+ sky130_fd_sc_hd__and2b_1
X_1453_ net485 Inst_LUT4AB_ConfigMem.Inst_frame8_bit8.Q _0513_ _0524_ _0525_ VGND
+ VGND VPWR VPWR _0000_ sky130_fd_sc_hd__a32o_1
Xoutput339 net339 VGND VGND VPWR VPWR SS4BEG[5] sky130_fd_sc_hd__buf_2
Xoutput317 net317 VGND VGND VPWR VPWR S4BEG[14] sky130_fd_sc_hd__buf_2
Xoutput328 net328 VGND VGND VPWR VPWR SS4BEG[0] sky130_fd_sc_hd__buf_2
Xoutput306 net306 VGND VGND VPWR VPWR S2BEGb[2] sky130_fd_sc_hd__buf_2
X_1522_ net761 net706 VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_67_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1384_ net60 net815 net88 net661 Inst_LUT4AB_ConfigMem.Inst_frame13_bit25.Q Inst_LUT4AB_ConfigMem.Inst_frame13_bit26.Q
+ VGND VGND VPWR VPWR _0488_ sky130_fd_sc_hd__mux4_1
X_2005_ net766 net696 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_50_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_33_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrebuffer60 net453 VGND VGND VPWR VPWR net452 sky130_fd_sc_hd__buf_6
XFILLER_64_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_29 FrameStrobe[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_18 EE4END[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_0884_ net661 net658 net638 net648 Inst_LUT4AB_ConfigMem.Inst_frame3_bit2.Q Inst_LUT4AB_ConfigMem.Inst_frame3_bit3.Q
+ VGND VGND VPWR VPWR _0036_ sky130_fd_sc_hd__mux4_1
X_0953_ net660 net657 net652 net637 Inst_LUT4AB_ConfigMem.Inst_frame2_bit14.Q Inst_LUT4AB_ConfigMem.Inst_frame2_bit15.Q
+ VGND VGND VPWR VPWR _0100_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_30_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1367_ _0469_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit9.Q _0471_ _0474_ VGND VGND VPWR
+ VPWR Inst_LUT4AB_switch_matrix.E6BEG1 sky130_fd_sc_hd__a22o_1
Xoutput169 net169 VGND VGND VPWR VPWR E6BEG[7] sky130_fd_sc_hd__buf_2
Xoutput158 net158 VGND VGND VPWR VPWR E2BEGb[6] sky130_fd_sc_hd__buf_2
Xoutput147 net147 VGND VGND VPWR VPWR E2BEG[3] sky130_fd_sc_hd__buf_4
X_1505_ net801 net705 VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3
+ sky130_fd_sc_hd__dlxtp_1
X_1436_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit30.Q _0508_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit31.Q
+ _0507_ VGND VGND VPWR VPWR _0509_ sky130_fd_sc_hd__a211o_1
XFILLER_62_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_38_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1298_ _0412_ _0414_ _0417_ _0592_ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.E2BEG0
+ sky130_fd_sc_hd__a22o_1
XFILLER_62_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput38 FrameData[19] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__buf_1
Xinput49 FrameData[5] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput27 EE4END[3] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput16 E2MID[2] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__clkbuf_2
X_2270_ net400 VGND VGND VPWR VPWR net303 sky130_fd_sc_hd__buf_6
X_1221_ Inst_LUT4AB_switch_matrix.JN2BEG5 Inst_LUT4AB_switch_matrix.E2BEG5 Inst_LUT4AB_ConfigMem.Inst_frame8_bit20.Q
+ VGND VGND VPWR VPWR _0350_ sky130_fd_sc_hd__mux2_4
XFILLER_6_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1152_ _0242_ _0270_ _0284_ VGND VGND VPWR VPWR _0285_ sky130_fd_sc_hd__a21oi_2
X_1083_ _0219_ _0220_ VGND VGND VPWR VPWR _0221_ sky130_fd_sc_hd__or2_1
XFILLER_37_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_35_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1985_ net802 net692 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0936_ _0083_ _0080_ _0074_ _0076_ VGND VGND VPWR VPWR _0084_ sky130_fd_sc_hd__a31o_1
XFILLER_20_103 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0867_ Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 _0018_ _0019_ Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4
+ VGND VGND VPWR VPWR _0020_ sky130_fd_sc_hd__o22a_1
X_0798_ net659 net654 net649 net644 Inst_LUT4AB_ConfigMem.Inst_frame2_bit6.Q Inst_LUT4AB_ConfigMem.Inst_frame2_bit7.Q
+ VGND VGND VPWR VPWR _0645_ sky130_fd_sc_hd__mux4_2
X_1419_ net644 Inst_LUT4AB_switch_matrix.E2BEG3 _0192_ _0043_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit11.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame12_bit10.Q VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.S1BEG0
+ sky130_fd_sc_hd__mux4_2
XFILLER_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_40_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1770_ net782 net742 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame10_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0721_ Inst_LE_LUT4c_frame_config_dffesr.c_reset_value VGND VGND VPWR VPWR _0572_
+ sky130_fd_sc_hd__inv_1
XFILLER_6_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2253_ NN4END[14] VGND VGND VPWR VPWR net277 sky130_fd_sc_hd__buf_1
XFILLER_69_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2322_ Inst_LUT4AB_switch_matrix.JW2BEG6 VGND VGND VPWR VPWR net355 sky130_fd_sc_hd__buf_6
X_2184_ net767 VGND VGND VPWR VPWR net209 sky130_fd_sc_hd__clkbuf_1
X_1204_ _0073_ _0054_ VGND VGND VPWR VPWR _0334_ sky130_fd_sc_hd__nand2b_1
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1135_ _0268_ VGND VGND VPWR VPWR _0269_ sky130_fd_sc_hd__inv_2
X_1066_ _0083_ _0080_ _0074_ _0123_ _0076_ VGND VGND VPWR VPWR _0204_ sky130_fd_sc_hd__a311o_1
XFILLER_33_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0919_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit12.Q _0067_ VGND VGND VPWR VPWR _0068_
+ sky130_fd_sc_hd__and2b_1
Xclone19 D VGND VGND VPWR VPWR net411 sky130_fd_sc_hd__clkbuf_1
X_1899_ net779 net680 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame6_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1968_ net768 net687 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_17_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1822_ net807 net671 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame8_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_30_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1753_ net753 net740 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame10_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1684_ net789 net733 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame12_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0704_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit0.Q VGND VGND VPWR VPWR _0555_ sky130_fd_sc_hd__inv_1
X_2305_ SS4END[14] VGND VGND VPWR VPWR net329 sky130_fd_sc_hd__clkbuf_2
X_2236_ N4END[13] VGND VGND VPWR VPWR net275 sky130_fd_sc_hd__buf_1
X_2167_ net805 VGND VGND VPWR VPWR net191 sky130_fd_sc_hd__buf_1
XFILLER_72_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_68_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1049_ net86 net94 net88 net114 Inst_LUT4AB_ConfigMem.Inst_frame1_bit11.Q Inst_LUT4AB_ConfigMem.Inst_frame1_bit10.Q
+ VGND VGND VPWR VPWR _0189_ sky130_fd_sc_hd__mux4_1
X_1118_ net74 net19 net102 net130 Inst_LUT4AB_ConfigMem.Inst_frame6_bit22.Q Inst_LUT4AB_ConfigMem.Inst_frame6_bit23.Q
+ VGND VGND VPWR VPWR _0253_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_0_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2098_ net762 net744 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame0_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_21_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_8_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2021_ net794 net698 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_65_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1805_ net774 net668 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1736_ net786 net735 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame11_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1598_ net807 net717 VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1
+ sky130_fd_sc_hd__dlxtp_1
Xfanout726 net727 VGND VGND VPWR VPWR net726 sky130_fd_sc_hd__clkbuf_2
Xfanout748 net53 VGND VGND VPWR VPWR net748 sky130_fd_sc_hd__buf_4
Xfanout759 net760 VGND VGND VPWR VPWR net759 sky130_fd_sc_hd__clkbuf_4
Xfanout715 net716 VGND VGND VPWR VPWR net715 sky130_fd_sc_hd__buf_1
Xfanout737 net738 VGND VGND VPWR VPWR net737 sky130_fd_sc_hd__buf_2
X_1667_ net797 net728 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame13_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
Xfanout704 FrameStrobe[18] VGND VGND VPWR VPWR net704 sky130_fd_sc_hd__clkbuf_2
XANTENNA_119 net211 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_108 net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2219_ net69 VGND VGND VPWR VPWR net252 sky130_fd_sc_hd__buf_1
XFILLER_41_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_348 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput307 net307 VGND VGND VPWR VPWR S2BEGb[3] sky130_fd_sc_hd__buf_2
X_1452_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit8.Q _0513_ _0523_ Inst_LH_LUT4c_frame_config_dffesr.c_reset_value
+ VGND VGND VPWR VPWR _0525_ sky130_fd_sc_hd__o2bb2a_4
X_1383_ _0487_ _0486_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit30.Q VGND VGND VPWR VPWR
+ Inst_LUT4AB_switch_matrix.EE4BEG2 sky130_fd_sc_hd__mux2_1
Xoutput318 net318 VGND VGND VPWR VPWR S4BEG[15] sky130_fd_sc_hd__buf_2
Xoutput329 net329 VGND VGND VPWR VPWR SS4BEG[10] sky130_fd_sc_hd__buf_2
X_1521_ net763 net706 VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_27_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2004_ net790 net695 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_33_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1719_ net757 net738 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame11_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
Xrebuffer61 net454 VGND VGND VPWR VPWR net453 sky130_fd_sc_hd__buf_6
XFILLER_41_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_226 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0952_ net66 net11 net110 net122 Inst_LUT4AB_ConfigMem.Inst_frame5_bit14.Q Inst_LUT4AB_ConfigMem.Inst_frame5_bit15.Q
+ VGND VGND VPWR VPWR _0099_ sky130_fd_sc_hd__mux4_2
XANTENNA_19 EE4END[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput159 net159 VGND VGND VPWR VPWR E2BEGb[7] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_30_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput148 net148 VGND VGND VPWR VPWR E2BEG[4] sky130_fd_sc_hd__buf_2
X_0883_ _0035_ Inst_LB_LUT4c_frame_config_dffesr.LUT_flop Inst_LB_LUT4c_frame_config_dffesr.c_out_mux
+ VGND VGND VPWR VPWR B sky130_fd_sc_hd__mux2_4
X_1504_ net804 net705 VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2
+ sky130_fd_sc_hd__dlxtp_1
X_1366_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit8.Q _0473_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit9.Q
+ VGND VGND VPWR VPWR _0474_ sky130_fd_sc_hd__a21oi_1
X_1435_ _0192_ _0139_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit29.Q VGND VGND VPWR VPWR
+ _0508_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_38_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1297_ _0415_ _0416_ _0591_ VGND VGND VPWR VPWR _0417_ sky130_fd_sc_hd__mux2_1
XFILLER_23_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput39 FrameData[1] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__clkbuf_2
Xinput28 FrameData[0] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput17 E2MID[3] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__buf_2
XFILLER_6_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1151_ _0283_ _0242_ _0282_ VGND VGND VPWR VPWR _0284_ sky130_fd_sc_hd__o21ai_2
X_1220_ _0349_ Inst_LD_LUT4c_frame_config_dffesr.LUT_flop Inst_LD_LUT4c_frame_config_dffesr.c_out_mux
+ VGND VGND VPWR VPWR D sky130_fd_sc_hd__mux2_4
XFILLER_35_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1082_ Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 _0213_ _0214_ Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2
+ VGND VGND VPWR VPWR _0220_ sky130_fd_sc_hd__a22o_1
XFILLER_45_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1984_ net803 net692 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_43_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0935_ _0011_ _0012_ _0023_ _0021_ _0081_ VGND VGND VPWR VPWR _0083_ sky130_fd_sc_hd__a311o_1
X_0866_ _0017_ _0016_ VGND VGND VPWR VPWR _0019_ sky130_fd_sc_hd__nand2b_1
XFILLER_20_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0797_ Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12
+ _0643_ VGND VGND VPWR VPWR _0644_ sky130_fd_sc_hd__mux2_4
XFILLER_68_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_259 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1349_ net626 _0652_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit29.Q VGND VGND VPWR VPWR
+ _0459_ sky130_fd_sc_hd__mux2_1
X_1418_ net424 _0093_ Inst_LUT4AB_switch_matrix.E2BEG0 _0098_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit12.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame12_bit13.Q VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.S1BEG1
+ sky130_fd_sc_hd__mux4_1
XFILLER_73_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0720_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit17.Q VGND VGND VPWR VPWR _0571_ sky130_fd_sc_hd__inv_1
XTAP_TAPCELL_ROW_40_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2252_ NN4END[13] VGND VGND VPWR VPWR net291 sky130_fd_sc_hd__buf_1
X_1134_ _0254_ _0266_ VGND VGND VPWR VPWR _0268_ sky130_fd_sc_hd__nand2_1
X_1203_ Inst_LD_LUT4c_frame_config_dffesr.c_I0mux _0080_ _0083_ _0332_ VGND VGND VPWR
+ VPWR _0333_ sky130_fd_sc_hd__a31o_1
X_2183_ net769 VGND VGND VPWR VPWR net208 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_63_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1065_ _0203_ Inst_LC_LUT4c_frame_config_dffesr.LUT_flop Inst_LC_LUT4c_frame_config_dffesr.c_out_mux
+ VGND VGND VPWR VPWR C sky130_fd_sc_hd__mux2_4
X_0918_ net58 net66 net3 net11 Inst_LUT4AB_ConfigMem.Inst_frame2_bit10.Q Inst_LUT4AB_ConfigMem.Inst_frame2_bit11.Q
+ VGND VGND VPWR VPWR _0067_ sky130_fd_sc_hd__mux4_1
X_1898_ net782 net681 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame6_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0849_ Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2
+ _0643_ VGND VGND VPWR VPWR _0692_ sky130_fd_sc_hd__mux2_1
X_1967_ net770 net687 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_68_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_54_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_17_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1821_ net809 net671 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame8_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1683_ net28 net734 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame12_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_30_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0703_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit5.Q VGND VGND VPWR VPWR _0554_ sky130_fd_sc_hd__inv_2
X_1752_ net755 net740 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame10_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2304_ SS4END[13] VGND VGND VPWR VPWR net343 sky130_fd_sc_hd__clkbuf_2
X_2166_ net807 VGND VGND VPWR VPWR net190 sky130_fd_sc_hd__buf_1
X_2235_ N4END[12] VGND VGND VPWR VPWR net274 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_68_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1117_ net18 net129 net101 Inst_LUT4AB_switch_matrix.JS2BEG6 Inst_LUT4AB_ConfigMem.Inst_frame7_bit23.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame7_bit22.Q VGND VGND VPWR VPWR _0252_ sky130_fd_sc_hd__mux4_2
XFILLER_38_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2097_ net764 net744 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame0_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_51_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1048_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit12.Q _0187_ VGND VGND VPWR VPWR _0188_
+ sky130_fd_sc_hd__and2b_1
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2020_ net796 net697 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_35_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1804_ net777 net668 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1735_ net788 net735 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame11_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1666_ net799 net728 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame13_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1597_ net809 net718 VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0
+ sky130_fd_sc_hd__dlxtp_1
Xfanout727 net729 VGND VGND VPWR VPWR net727 sky130_fd_sc_hd__clkbuf_2
Xfanout716 FrameStrobe[16] VGND VGND VPWR VPWR net716 sky130_fd_sc_hd__clkbuf_2
Xfanout738 FrameStrobe[11] VGND VGND VPWR VPWR net738 sky130_fd_sc_hd__clkbuf_2
Xfanout749 net750 VGND VGND VPWR VPWR net749 sky130_fd_sc_hd__clkbuf_4
Xfanout705 net706 VGND VGND VPWR VPWR net705 sky130_fd_sc_hd__clkbuf_2
X_2149_ EE4END[14] VGND VGND VPWR VPWR net173 sky130_fd_sc_hd__buf_1
X_2218_ Inst_LUT4AB_switch_matrix.JN2BEG7 VGND VGND VPWR VPWR net251 sky130_fd_sc_hd__clkbuf_1
XFILLER_41_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_109 net111 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput319 net319 VGND VGND VPWR VPWR S4BEG[1] sky130_fd_sc_hd__buf_2
Xoutput308 net308 VGND VGND VPWR VPWR S2BEGb[4] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_10_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1520_ net767 net704 VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.c_reset_value
+ sky130_fd_sc_hd__dlxtp_1
X_1451_ _0323_ _0523_ VGND VGND VPWR VPWR _0524_ sky130_fd_sc_hd__nand2b_1
X_1382_ net57 net85 net2 net658 Inst_LUT4AB_ConfigMem.Inst_frame13_bit29.Q Inst_LUT4AB_ConfigMem.Inst_frame13_bit28.Q
+ VGND VGND VPWR VPWR _0487_ sky130_fd_sc_hd__mux4_1
XFILLER_4_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2003_ net812 net695 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_50_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_33_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1649_ net764 net722 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame14_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1718_ net48 net738 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame11_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
Xrebuffer62 net398 VGND VGND VPWR VPWR net454 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_41_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_30_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0882_ _0014_ _0027_ _0034_ VGND VGND VPWR VPWR _0035_ sky130_fd_sc_hd__o21a_1
X_0951_ net78 net110 net121 Inst_LUT4AB_switch_matrix.JS2BEG3 Inst_LUT4AB_ConfigMem.Inst_frame0_bit14.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame0_bit15.Q VGND VGND VPWR VPWR _0098_ sky130_fd_sc_hd__mux4_2
XPHY_EDGE_ROW_34_Left_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput149 net149 VGND VGND VPWR VPWR E2BEG[5] sky130_fd_sc_hd__buf_4
X_1503_ net806 net703 VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1
+ sky130_fd_sc_hd__dlxtp_1
X_1365_ _0472_ VGND VGND VPWR VPWR _0473_ sky130_fd_sc_hd__inv_1
XTAP_TAPCELL_ROW_38_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1296_ net60 net62 net78 net25 Inst_LUT4AB_ConfigMem.Inst_frame4_bit26.Q Inst_LUT4AB_ConfigMem.Inst_frame4_bit27.Q
+ VGND VGND VPWR VPWR _0416_ sky130_fd_sc_hd__mux4_1
X_1434_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit30.Q _0506_ VGND VGND VPWR VPWR _0507_
+ sky130_fd_sc_hd__and2b_1
XFILLER_63_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_46_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_43_Left_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_52_Left_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_61_Left_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_32 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput18 E2MID[4] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_70_Left_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput29 FrameData[10] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1150_ Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10
+ Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14
+ _0266_ _0254_ VGND VGND VPWR VPWR _0283_ sky130_fd_sc_hd__mux4_1
X_1081_ Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 _0210_ _0212_ Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6
+ VGND VGND VPWR VPWR _0219_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_43_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1983_ net805 net692 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0865_ _0016_ _0017_ VGND VGND VPWR VPWR _0018_ sky130_fd_sc_hd__nand2b_1
X_0934_ _0012_ _0011_ _0023_ _0021_ VGND VGND VPWR VPWR _0082_ sky130_fd_sc_hd__a31o_1
X_0796_ _0551_ net1 _0642_ VGND VGND VPWR VPWR _0643_ sky130_fd_sc_hd__o21ai_4
X_1417_ net399 Inst_LUT4AB_switch_matrix.E2BEG1 net664 _0271_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit15.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame12_bit14.Q VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.S1BEG2
+ sky130_fd_sc_hd__mux4_2
XFILLER_68_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1279_ net60 net7 net62 net813 Inst_LUT4AB_ConfigMem.Inst_frame2_bit27.Q Inst_LUT4AB_ConfigMem.Inst_frame2_bit26.Q
+ VGND VGND VPWR VPWR _0401_ sky130_fd_sc_hd__mux4_1
X_1348_ _0071_ _0130_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit29.Q VGND VGND VPWR VPWR
+ _0458_ sky130_fd_sc_hd__mux2_4
XFILLER_22_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_5_Left_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2251_ NN4END[12] VGND VGND VPWR VPWR net290 sky130_fd_sc_hd__buf_1
X_2320_ Inst_LUT4AB_switch_matrix.JW2BEG4 VGND VGND VPWR VPWR net353 sky130_fd_sc_hd__buf_6
XFILLER_65_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1133_ _0266_ _0254_ VGND VGND VPWR VPWR _0267_ sky130_fd_sc_hd__or2_4
X_1202_ Inst_LD_LUT4c_frame_config_dffesr.c_I0mux _0331_ VGND VGND VPWR VPWR _0332_
+ sky130_fd_sc_hd__and2b_1
X_1064_ _0202_ _0197_ _0193_ VGND VGND VPWR VPWR _0203_ sky130_fd_sc_hd__mux2_4
X_2182_ net771 VGND VGND VPWR VPWR net207 sky130_fd_sc_hd__clkbuf_2
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1966_ net773 net687 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_18_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0917_ _0064_ _0065_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit12.Q VGND VGND VPWR VPWR
+ _0066_ sky130_fd_sc_hd__mux2_4
X_1897_ net784 net682 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame6_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0779_ _0623_ _0548_ _0625_ _0627_ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.JN2BEG3
+ sky130_fd_sc_hd__o22a_4
X_0848_ _0690_ _0689_ _0620_ VGND VGND VPWR VPWR _0691_ sky130_fd_sc_hd__mux2_1
XFILLER_0_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_78 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1820_ net747 net671 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame8_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1682_ net762 net729 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame13_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0702_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit9.Q VGND VGND VPWR VPWR _0553_ sky130_fd_sc_hd__inv_1
X_1751_ net757 net740 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame10_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2303_ SS4END[12] VGND VGND VPWR VPWR net342 sky130_fd_sc_hd__clkbuf_2
X_2234_ N4END[11] VGND VGND VPWR VPWR net273 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_68_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1116_ _0575_ _0247_ _0249_ _0251_ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.JS2BEG6
+ sky130_fd_sc_hd__o22a_4
X_2165_ net809 VGND VGND VPWR VPWR net189 sky130_fd_sc_hd__buf_1
X_1047_ net58 net66 net3 net11 Inst_LUT4AB_ConfigMem.Inst_frame1_bit10.Q Inst_LUT4AB_ConfigMem.Inst_frame1_bit11.Q
+ VGND VGND VPWR VPWR _0187_ sky130_fd_sc_hd__mux4_1
XFILLER_38_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2096_ net767 net744 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame0_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1949_ net810 net688 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_51_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_8_Left_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_73_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1803_ net42 net667 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_13_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1596_ net747 net717 VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.c_reset_value
+ sky130_fd_sc_hd__dlxtp_1
X_1734_ net792 net736 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame11_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1665_ net801 net728 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame13_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
Xfanout706 FrameStrobe[18] VGND VGND VPWR VPWR net706 sky130_fd_sc_hd__buf_1
X_2217_ Inst_LUT4AB_switch_matrix.JN2BEG6 VGND VGND VPWR VPWR net250 sky130_fd_sc_hd__buf_1
Xfanout717 net720 VGND VGND VPWR VPWR net717 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_31_Right_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout728 FrameStrobe[13] VGND VGND VPWR VPWR net728 sky130_fd_sc_hd__buf_2
Xfanout739 net741 VGND VGND VPWR VPWR net739 sky130_fd_sc_hd__buf_2
XFILLER_53_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2079_ net806 net743 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame0_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2148_ EE4END[13] VGND VGND VPWR VPWR net187 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_40_Right_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1450_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit17.Q _0522_ VGND VGND VPWR VPWR _0523_
+ sky130_fd_sc_hd__nand2_1
XFILLER_4_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput309 net309 VGND VGND VPWR VPWR S2BEGb[5] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_10_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1381_ net653 _0120_ net664 _0159_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit28.Q Inst_LUT4AB_ConfigMem.Inst_frame13_bit29.Q
+ VGND VGND VPWR VPWR _0486_ sky130_fd_sc_hd__mux4_1
XFILLER_35_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2002_ net761 net691 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_33_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1579_ net779 net716 VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1
+ sky130_fd_sc_hd__dlxtp_1
X_1648_ net768 net722 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame14_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1717_ net766 net738 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame11_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
Xrebuffer41 net454 VGND VGND VPWR VPWR net433 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_41_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_103 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0950_ _0096_ _0084_ Inst_LE_LUT4c_frame_config_dffesr.c_I0mux VGND VGND VPWR VPWR
+ _0097_ sky130_fd_sc_hd__mux2_4
X_0881_ _0030_ _0033_ _0014_ VGND VGND VPWR VPWR _0034_ sky130_fd_sc_hd__or3b_1
XFILLER_20_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput139 net139 VGND VGND VPWR VPWR Co sky130_fd_sc_hd__buf_6
X_1502_ net807 net703 VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0
+ sky130_fd_sc_hd__dlxtp_1
X_1433_ _0280_ _0674_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit29.Q VGND VGND VPWR VPWR
+ _0506_ sky130_fd_sc_hd__mux2_4
X_1364_ net653 net638 net647 net642 Inst_LUT4AB_ConfigMem.Inst_frame12_bit6.Q Inst_LUT4AB_ConfigMem.Inst_frame12_bit7.Q
+ VGND VGND VPWR VPWR _0472_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_38_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1295_ net813 net118 net90 net134 Inst_LUT4AB_ConfigMem.Inst_frame4_bit27.Q Inst_LUT4AB_ConfigMem.Inst_frame4_bit26.Q
+ VGND VGND VPWR VPWR _0415_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_46_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput19 E2MID[5] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__clkbuf_2
XFILLER_10_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_158 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1080_ _0138_ _0139_ _0130_ _0129_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit27.Q Inst_LUT4AB_ConfigMem.Inst_frame9_bit28.Q
+ VGND VGND VPWR VPWR _0218_ sky130_fd_sc_hd__mux4_2
XFILLER_60_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1982_ net808 net692 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_52_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0933_ _0077_ _0078_ VGND VGND VPWR VPWR _0081_ sky130_fd_sc_hd__and2_1
X_0864_ _0616_ _0617_ _0606_ _0605_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit15.Q Inst_LUT4AB_ConfigMem.Inst_frame10_bit16.Q
+ VGND VGND VPWR VPWR _0017_ sky130_fd_sc_hd__mux4_2
X_0795_ _0641_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit4.Q _0631_ Inst_LA_LUT4c_frame_config_dffesr.c_I0mux
+ VGND VGND VPWR VPWR _0642_ sky130_fd_sc_hd__a211o_1
XPHY_EDGE_ROW_21_Left_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1347_ net60 net815 net665 net663 Inst_LUT4AB_ConfigMem.Inst_frame12_bit29.Q Inst_LUT4AB_ConfigMem.Inst_frame12_bit30.Q
+ VGND VGND VPWR VPWR _0457_ sky130_fd_sc_hd__mux4_1
X_1416_ net626 _0653_ Inst_LUT4AB_switch_matrix.E2BEG2 _0639_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit16.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame12_bit17.Q VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.S1BEG3
+ sky130_fd_sc_hd__mux4_2
X_1278_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit28.Q _0399_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit29.Q
+ VGND VGND VPWR VPWR _0400_ sky130_fd_sc_hd__o21a_1
XFILLER_3_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_57_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_69_Right_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_286 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2250_ NN4END[11] VGND VGND VPWR VPWR net289 sky130_fd_sc_hd__buf_1
X_1201_ _0329_ _0330_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit2.Q VGND VGND VPWR VPWR
+ _0331_ sky130_fd_sc_hd__mux2_1
X_1132_ _0264_ _0265_ _0256_ _0255_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit1.Q Inst_LUT4AB_ConfigMem.Inst_frame8_bit2.Q
+ VGND VGND VPWR VPWR _0266_ sky130_fd_sc_hd__mux4_2
X_2181_ net775 VGND VGND VPWR VPWR net206 sky130_fd_sc_hd__clkbuf_1
X_1063_ _0201_ _0199_ _0170_ VGND VGND VPWR VPWR _0202_ sky130_fd_sc_hd__mux2_1
X_0916_ net641 net631 net410 net427 Inst_LUT4AB_ConfigMem.Inst_frame2_bit10.Q Inst_LUT4AB_ConfigMem.Inst_frame2_bit11.Q
+ VGND VGND VPWR VPWR _0065_ sky130_fd_sc_hd__mux4_2
X_1965_ net776 net687 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0778_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit8.Q _0626_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit9.Q
+ VGND VGND VPWR VPWR _0627_ sky130_fd_sc_hd__a21o_1
X_0847_ Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6
+ _0643_ VGND VGND VPWR VPWR _0690_ sky130_fd_sc_hd__mux2_1
X_1896_ net786 net679 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame6_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_71_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_3_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1750_ net760 net742 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame10_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1681_ net764 net729 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame13_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0701_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit8.Q VGND VGND VPWR VPWR _0552_ sky130_fd_sc_hd__inv_2
X_2302_ SS4END[11] VGND VGND VPWR VPWR net341 sky130_fd_sc_hd__clkbuf_2
X_2164_ net747 VGND VGND VPWR VPWR net219 sky130_fd_sc_hd__buf_1
X_2233_ N4END[10] VGND VGND VPWR VPWR net272 sky130_fd_sc_hd__clkbuf_1
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1115_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit20.Q _0250_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit21.Q
+ VGND VGND VPWR VPWR _0251_ sky130_fd_sc_hd__a21o_1
XFILLER_53_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_51_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1046_ _0184_ _0185_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit12.Q VGND VGND VPWR VPWR
+ _0186_ sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_0_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2095_ net769 net744 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame0_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1948_ net748 net687 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1879_ net757 net679 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame6_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_16_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_8_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1802_ net782 net667 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1733_ net794 net736 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame11_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_13_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout718 net719 VGND VGND VPWR VPWR net718 sky130_fd_sc_hd__clkbuf_2
X_1595_ net749 net717 VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.c_I0mux
+ sky130_fd_sc_hd__dlxtp_1
X_1664_ net803 net726 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame13_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
Xfanout707 net708 VGND VGND VPWR VPWR net707 sky130_fd_sc_hd__clkbuf_2
Xfanout729 FrameStrobe[13] VGND VGND VPWR VPWR net729 sky130_fd_sc_hd__clkbuf_2
XFILLER_38_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2147_ EE4END[12] VGND VGND VPWR VPWR net186 sky130_fd_sc_hd__clkbuf_1
X_2078_ net30 net746 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame0_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_34_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1029_ _0169_ _0082_ Inst_LC_LUT4c_frame_config_dffesr.c_I0mux VGND VGND VPWR VPWR
+ _0170_ sky130_fd_sc_hd__mux2_4
XFILLER_30_68 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1380_ _0484_ _0485_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit1.Q VGND VGND VPWR VPWR
+ Inst_LUT4AB_switch_matrix.EE4BEG3 sky130_fd_sc_hd__mux2_4
XFILLER_4_230 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2001_ net763 net691 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_35_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1716_ net789 net738 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame11_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1578_ net782 net716 VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0
+ sky130_fd_sc_hd__dlxtp_1
X_1647_ net770 net722 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame14_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
Xrebuffer20 net428 VGND VGND VPWR VPWR net412 sky130_fd_sc_hd__buf_6
XFILLER_14_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_115 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0880_ Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 _0023_ _0031_ _0032_
+ VGND VGND VPWR VPWR _0033_ sky130_fd_sc_hd__o211a_1
X_1432_ _0267_ _0294_ _0304_ _0306_ VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__a31o_1
X_1363_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit8.Q _0470_ VGND VGND VPWR VPWR _0471_
+ sky130_fd_sc_hd__or2_1
X_1501_ net809 net703 VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.c_reset_value
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_38_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1294_ _0591_ _0413_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit29.Q VGND VGND VPWR VPWR
+ _0414_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_46_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_56 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1981_ net810 net693 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0932_ _0079_ VGND VGND VPWR VPWR _0080_ sky130_fd_sc_hd__inv_2
X_0863_ _0652_ _0653_ _0662_ _0661_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit17.Q Inst_LUT4AB_ConfigMem.Inst_frame10_bit18.Q
+ VGND VGND VPWR VPWR _0016_ sky130_fd_sc_hd__mux4_2
X_0794_ _0639_ _0640_ _0549_ VGND VGND VPWR VPWR _0641_ sky130_fd_sc_hd__mux2_4
XFILLER_68_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1346_ _0456_ _0455_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit2.Q VGND VGND VPWR VPWR
+ Inst_LUT4AB_switch_matrix.SS4BEG2 sky130_fd_sc_hd__mux2_4
X_1415_ net813 net106 net91 net663 Inst_LUT4AB_ConfigMem.Inst_frame12_bit19.Q Inst_LUT4AB_ConfigMem.Inst_frame12_bit18.Q
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.S4BEG0 sky130_fd_sc_hd__mux4_1
X_1277_ net654 net634 net649 net644 Inst_LUT4AB_ConfigMem.Inst_frame2_bit27.Q Inst_LUT4AB_ConfigMem.Inst_frame2_bit26.Q
+ VGND VGND VPWR VPWR _0399_ sky130_fd_sc_hd__mux4_1
XFILLER_3_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_57_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2180_ net777 VGND VGND VPWR VPWR net205 sky130_fd_sc_hd__buf_1
X_1200_ _0159_ _0158_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit1.Q VGND VGND VPWR VPWR
+ _0330_ sky130_fd_sc_hd__mux2_1
XFILLER_65_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1062_ Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 _0079_ _0081_ Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6
+ _0200_ VGND VGND VPWR VPWR _0201_ sky130_fd_sc_hd__a221o_1
X_1131_ net72 net17 net100 net128 Inst_LUT4AB_ConfigMem.Inst_frame6_bit20.Q Inst_LUT4AB_ConfigMem.Inst_frame6_bit21.Q
+ VGND VGND VPWR VPWR _0265_ sky130_fd_sc_hd__mux4_2
X_1964_ net778 net689 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0915_ net661 net658 C net637 Inst_LUT4AB_ConfigMem.Inst_frame2_bit10.Q Inst_LUT4AB_ConfigMem.Inst_frame2_bit11.Q
+ VGND VGND VPWR VPWR _0064_ sky130_fd_sc_hd__mux4_1
X_1895_ net788 net679 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame6_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_21_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0777_ net814 net93 net121 net133 Inst_LUT4AB_ConfigMem.Inst_frame4_bit6.Q Inst_LUT4AB_ConfigMem.Inst_frame4_bit7.Q
+ VGND VGND VPWR VPWR _0626_ sky130_fd_sc_hd__mux4_1
X_0846_ Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4
+ _0643_ VGND VGND VPWR VPWR _0689_ sky130_fd_sc_hd__mux2_1
XFILLER_68_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclone5 net409 net401 Inst_LUT4AB_ConfigMem.Inst_frame14_bit16.Q VGND VGND VPWR VPWR
+ net397 sky130_fd_sc_hd__mux2_4
X_1329_ net650 _0120_ net664 _0063_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit20.Q Inst_LUT4AB_ConfigMem.Inst_frame11_bit21.Q
+ VGND VGND VPWR VPWR _0444_ sky130_fd_sc_hd__mux4_1
XFILLER_17_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_62_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_49_Left_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput290 net290 VGND VGND VPWR VPWR NN4BEG[8] sky130_fd_sc_hd__buf_2
XFILLER_58_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_58_Left_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_67_Left_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0700_ Inst_LA_LUT4c_frame_config_dffesr.c_I0mux VGND VGND VPWR VPWR _0551_ sky130_fd_sc_hd__inv_2
X_2301_ SS4END[10] VGND VGND VPWR VPWR net340 sky130_fd_sc_hd__clkbuf_2
X_1680_ net767 net729 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame13_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1114_ net88 net114 net96 net665 Inst_LUT4AB_ConfigMem.Inst_frame2_bit19.Q Inst_LUT4AB_ConfigMem.Inst_frame2_bit18.Q
+ VGND VGND VPWR VPWR _0250_ sky130_fd_sc_hd__mux4_1
X_2163_ net749 VGND VGND VPWR VPWR net218 sky130_fd_sc_hd__buf_1
X_2232_ N4END[9] VGND VGND VPWR VPWR net271 sky130_fd_sc_hd__clkbuf_1
XFILLER_65_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_51_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1045_ net641 net631 net627 net402 Inst_LUT4AB_ConfigMem.Inst_frame1_bit10.Q Inst_LUT4AB_ConfigMem.Inst_frame1_bit11.Q
+ VGND VGND VPWR VPWR _0185_ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_16_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2094_ net771 net744 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame0_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_21_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1878_ net759 net681 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame6_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0829_ net69 net14 net97 Inst_LUT4AB_switch_matrix.JW2BEG3 Inst_LUT4AB_ConfigMem.Inst_frame7_bit0.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame7_bit1.Q VGND VGND VPWR VPWR _0673_ sky130_fd_sc_hd__mux4_2
X_1947_ net750 net687 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_9_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_206 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_73_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1663_ net805 net726 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame13_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1801_ net784 net667 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1732_ net795 net736 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame11_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_13_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout719 net720 VGND VGND VPWR VPWR net719 sky130_fd_sc_hd__clkbuf_2
X_1594_ net751 net717 VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.c_out_mux
+ sky130_fd_sc_hd__dlxtp_1
Xfanout708 net711 VGND VGND VPWR VPWR net708 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2215_ Inst_LUT4AB_switch_matrix.JN2BEG4 VGND VGND VPWR VPWR net248 sky130_fd_sc_hd__buf_4
XFILLER_53_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2077_ net29 net746 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame0_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2146_ EE4END[11] VGND VGND VPWR VPWR net185 sky130_fd_sc_hd__clkbuf_1
X_1028_ _0167_ _0168_ _0159_ _0158_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit23.Q Inst_LUT4AB_ConfigMem.Inst_frame10_bit24.Q
+ VGND VGND VPWR VPWR _0169_ sky130_fd_sc_hd__mux4_1
XFILLER_14_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_70_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_102 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2000_ net768 net691 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1715_ net811 net738 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame11_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1646_ net773 net721 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame14_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1577_ net784 net714 VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.c_reset_value
+ sky130_fd_sc_hd__dlxtp_1
X_2129_ E6END[4] VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__buf_1
Xrebuffer10 Inst_LUT4AB_switch_matrix.M_AD VGND VGND VPWR VPWR net402 sky130_fd_sc_hd__buf_6
Xrebuffer54 net447 VGND VGND VPWR VPWR net446 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_24_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1500_ net747 net705 VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.c_I0mux
+ sky130_fd_sc_hd__dlxtp_1
X_1362_ net816 net666 net661 net658 Inst_LUT4AB_ConfigMem.Inst_frame12_bit6.Q Inst_LUT4AB_ConfigMem.Inst_frame12_bit7.Q
+ VGND VGND VPWR VPWR _0470_ sky130_fd_sc_hd__mux4_1
X_1431_ net650 Inst_LUT4AB_switch_matrix.JW2BEG3 _0192_ _0043_ Inst_LUT4AB_ConfigMem.Inst_frame14_bit19.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame14_bit18.Q VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.N1BEG0
+ sky130_fd_sc_hd__mux4_1
X_1293_ net639 net629 net624 net622 Inst_LUT4AB_ConfigMem.Inst_frame4_bit26.Q Inst_LUT4AB_ConfigMem.Inst_frame4_bit27.Q
+ VGND VGND VPWR VPWR _0413_ sky130_fd_sc_hd__mux4_1
XFILLER_55_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_46_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1629_ net809 net724 VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_36_68 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_30_Left_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0931_ _0077_ _0078_ VGND VGND VPWR VPWR _0079_ sky130_fd_sc_hd__nor2_2
X_1980_ net748 net691 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_13_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0862_ _0673_ _0674_ _0683_ _0682_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit19.Q Inst_LUT4AB_ConfigMem.Inst_frame10_bit20.Q
+ VGND VGND VPWR VPWR _0015_ sky130_fd_sc_hd__mux4_2
X_0793_ net67 net112 net12 net123 Inst_LUT4AB_ConfigMem.Inst_frame6_bit27.Q Inst_LUT4AB_ConfigMem.Inst_frame6_bit26.Q
+ VGND VGND VPWR VPWR _0640_ sky130_fd_sc_hd__mux4_2
XFILLER_68_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1345_ net57 net113 net2 net655 Inst_LUT4AB_ConfigMem.Inst_frame11_bit1.Q Inst_LUT4AB_ConfigMem.Inst_frame11_bit0.Q
+ VGND VGND VPWR VPWR _0456_ sky130_fd_sc_hd__mux4_1
X_1276_ _0587_ _0397_ VGND VGND VPWR VPWR _0398_ sky130_fd_sc_hd__or2_1
X_1414_ net814 net107 net92 net655 Inst_LUT4AB_ConfigMem.Inst_frame12_bit21.Q Inst_LUT4AB_ConfigMem.Inst_frame12_bit20.Q
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.S4BEG1 sky130_fd_sc_hd__mux4_1
XFILLER_51_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_57_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1130_ net71 net127 net99 Inst_LUT4AB_switch_matrix.E2BEG6 Inst_LUT4AB_ConfigMem.Inst_frame7_bit21.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame7_bit20.Q VGND VGND VPWR VPWR _0264_ sky130_fd_sc_hd__mux4_2
XFILLER_2_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1061_ Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 _0171_ _0172_ Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2
+ VGND VGND VPWR VPWR _0200_ sky130_fd_sc_hd__a22o_1
X_1963_ net780 net689 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1894_ net791 net681 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame6_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0914_ net65 net10 net111 net121 Inst_LUT4AB_ConfigMem.Inst_frame5_bit6.Q Inst_LUT4AB_ConfigMem.Inst_frame5_bit7.Q
+ VGND VGND VPWR VPWR _0063_ sky130_fd_sc_hd__mux4_2
X_0845_ _0687_ _0665_ _0663_ VGND VGND VPWR VPWR _0688_ sky130_fd_sc_hd__mux2_1
X_0776_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit8.Q _0624_ VGND VGND VPWR VPWR _0625_
+ sky130_fd_sc_hd__and2b_1
XFILLER_68_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1259_ net85 net113 net89 net115 Inst_LUT4AB_ConfigMem.Inst_frame2_bit23.Q Inst_LUT4AB_ConfigMem.Inst_frame2_bit22.Q
+ VGND VGND VPWR VPWR _0384_ sky130_fd_sc_hd__mux4_1
Xclone6 net417 _0396_ Inst_LUT4AB_ConfigMem.Inst_frame14_bit17.Q VGND VGND VPWR VPWR
+ net398 sky130_fd_sc_hd__mux2_4
X_1328_ _0442_ _0443_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit25.Q VGND VGND VPWR VPWR
+ Inst_LUT4AB_switch_matrix.WW4BEG3 sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_62_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput291 net291 VGND VGND VPWR VPWR NN4BEG[9] sky130_fd_sc_hd__buf_2
Xoutput280 Inst_LUT4AB_switch_matrix.NN4BEG1 VGND VGND VPWR VPWR NN4BEG[13] sky130_fd_sc_hd__buf_6
XFILLER_58_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_2_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2300_ SS4END[9] VGND VGND VPWR VPWR net339 sky130_fd_sc_hd__clkbuf_2
X_2231_ N4END[8] VGND VGND VPWR VPWR net270 sky130_fd_sc_hd__clkbuf_1
X_1113_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit20.Q _0248_ VGND VGND VPWR VPWR _0249_
+ sky130_fd_sc_hd__and2b_1
X_2162_ net751 VGND VGND VPWR VPWR net217 sky130_fd_sc_hd__buf_1
XFILLER_53_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1044_ net660 net656 net652 net636 Inst_LUT4AB_ConfigMem.Inst_frame1_bit10.Q Inst_LUT4AB_ConfigMem.Inst_frame1_bit11.Q
+ VGND VGND VPWR VPWR _0184_ sky130_fd_sc_hd__mux4_1
X_2093_ net774 net744 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_61_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1877_ net766 net681 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame6_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1946_ net752 net56 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0759_ net659 net654 net649 net644 Inst_LUT4AB_ConfigMem.Inst_frame3_bit6.Q Inst_LUT4AB_ConfigMem.Inst_frame3_bit7.Q
+ VGND VGND VPWR VPWR _0609_ sky130_fd_sc_hd__mux4_2
X_0828_ _0668_ _0561_ _0670_ _0672_ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.JW2BEG3
+ sky130_fd_sc_hd__o22a_4
XFILLER_28_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_73_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1800_ net785 net667 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_43_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1731_ net798 net737 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame11_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1662_ net808 net726 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame13_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1593_ net753 net717 VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15
+ sky130_fd_sc_hd__dlxtp_1
X_2214_ Inst_LUT4AB_switch_matrix.JN2BEG3 VGND VGND VPWR VPWR net247 sky130_fd_sc_hd__buf_6
Xfanout709 net711 VGND VGND VPWR VPWR net709 sky130_fd_sc_hd__clkbuf_2
XFILLER_53_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2145_ EE4END[10] VGND VGND VPWR VPWR net184 sky130_fd_sc_hd__clkbuf_1
X_1027_ net76 net21 net104 net132 Inst_LUT4AB_ConfigMem.Inst_frame6_bit2.Q Inst_LUT4AB_ConfigMem.Inst_frame6_bit3.Q
+ VGND VGND VPWR VPWR _0168_ sky130_fd_sc_hd__mux4_1
XFILLER_26_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2076_ net747 net744 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame0_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1929_ net783 net685 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame5_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_39_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_70_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_114 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_27_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold90 Inst_LF_LUT4c_frame_config_dffesr.LUT_flop VGND VGND VPWR VPWR net482 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_35_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1576_ net785 net714 VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.c_I0mux
+ sky130_fd_sc_hd__dlxtp_1
X_1714_ net762 net731 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame12_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1645_ net776 net721 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame14_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
Xrebuffer11 net402 VGND VGND VPWR VPWR net403 sky130_fd_sc_hd__buf_6
X_2128_ E6END[3] VGND VGND VPWR VPWR net163 sky130_fd_sc_hd__buf_1
Xrebuffer33 Inst_LUT4AB_switch_matrix.M_AD VGND VGND VPWR VPWR net425 sky130_fd_sc_hd__clkbuf_2
Xrebuffer22 Inst_LUT4AB_switch_matrix.M_AH VGND VGND VPWR VPWR net414 sky130_fd_sc_hd__buf_6
Xrebuffer55 net448 VGND VGND VPWR VPWR net447 sky130_fd_sc_hd__buf_6
X_2059_ net780 net702 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_24_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_25 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1430_ net637 _0093_ Inst_LUT4AB_switch_matrix.JW2BEG0 _0098_ Inst_LUT4AB_ConfigMem.Inst_frame14_bit20.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame14_bit21.Q VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.N1BEG1
+ sky130_fd_sc_hd__mux4_1
X_1361_ _0468_ _0467_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit8.Q VGND VGND VPWR VPWR
+ _0469_ sky130_fd_sc_hd__mux2_4
XFILLER_48_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1292_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit28.Q _0411_ VGND VGND VPWR VPWR _0412_
+ sky130_fd_sc_hd__or2_1
XFILLER_63_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1628_ net747 net724 VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12
+ sky130_fd_sc_hd__dlxtp_1
X_1559_ net758 net712 VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_46_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_223 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0930_ _0071_ _0072_ _0063_ _0062_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit27.Q Inst_LUT4AB_ConfigMem.Inst_frame10_bit28.Q
+ VGND VGND VPWR VPWR _0078_ sky130_fd_sc_hd__mux4_2
XFILLER_9_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0861_ _0012_ _0011_ Inst_LB_LUT4c_frame_config_dffesr.c_I0mux _0013_ VGND VGND VPWR
+ VPWR _0014_ sky130_fd_sc_hd__a31o_1
X_0792_ net84 net135 net108 Inst_LUT4AB_switch_matrix.JN2BEG1 Inst_LUT4AB_ConfigMem.Inst_frame1_bit27.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame1_bit26.Q VGND VGND VPWR VPWR _0639_ sky130_fd_sc_hd__mux4_2
XFILLER_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1413_ net89 net134 net108 net651 Inst_LUT4AB_ConfigMem.Inst_frame12_bit23.Q Inst_LUT4AB_ConfigMem.Inst_frame12_bit22.Q
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.S4BEG2 sky130_fd_sc_hd__mux4_1
XFILLER_36_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1344_ net651 _0120_ net664 _0183_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit0.Q Inst_LUT4AB_ConfigMem.Inst_frame11_bit1.Q
+ VGND VGND VPWR VPWR _0455_ sky130_fd_sc_hd__mux4_1
XFILLER_3_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1275_ net639 net629 net624 net397 Inst_LUT4AB_ConfigMem.Inst_frame2_bit26.Q Inst_LUT4AB_ConfigMem.Inst_frame2_bit27.Q
+ VGND VGND VPWR VPWR _0397_ sky130_fd_sc_hd__mux4_1
XFILLER_59_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_29_Right_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_38_Right_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_47_Right_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_25_Left_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1060_ Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 _0081_ _0172_ Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3
+ _0198_ VGND VGND VPWR VPWR _0199_ sky130_fd_sc_hd__a221o_1
X_1962_ net781 net689 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_56_Right_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1893_ net793 net681 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame6_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0913_ net82 net25 net106 Inst_LUT4AB_switch_matrix.JS2BEG2 Inst_LUT4AB_ConfigMem.Inst_frame0_bit6.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame0_bit7.Q VGND VGND VPWR VPWR _0062_ sky130_fd_sc_hd__mux4_2
X_0844_ _0686_ _0685_ _0620_ VGND VGND VPWR VPWR _0687_ sky130_fd_sc_hd__mux2_1
X_0775_ net65 net816 net77 net10 Inst_LUT4AB_ConfigMem.Inst_frame4_bit7.Q Inst_LUT4AB_ConfigMem.Inst_frame4_bit6.Q
+ VGND VGND VPWR VPWR _0624_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_65_Right_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1189_ Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 _0304_ _0319_ _0320_
+ VGND VGND VPWR VPWR _0321_ sky130_fd_sc_hd__o211a_1
XFILLER_68_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1258_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit24.Q _0382_ VGND VGND VPWR VPWR _0383_
+ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_54_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1327_ net645 net431 _0252_ _0662_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit23.Q Inst_LUT4AB_ConfigMem.Inst_frame11_bit24.Q
+ VGND VGND VPWR VPWR _0443_ sky130_fd_sc_hd__mux4_1
Xclone7 G VGND VGND VPWR VPWR net399 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_19_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput270 net270 VGND VGND VPWR VPWR N4BEG[4] sky130_fd_sc_hd__buf_2
XFILLER_3_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput281 net281 VGND VGND VPWR VPWR NN4BEG[14] sky130_fd_sc_hd__clkbuf_4
XFILLER_59_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput292 Inst_LUT4AB_switch_matrix.S1BEG0 VGND VGND VPWR VPWR S1BEG[0] sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_2_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2230_ N4END[7] VGND VGND VPWR VPWR net269 sky130_fd_sc_hd__clkbuf_1
X_1112_ net60 net68 net5 net13 Inst_LUT4AB_ConfigMem.Inst_frame2_bit18.Q Inst_LUT4AB_ConfigMem.Inst_frame2_bit19.Q
+ VGND VGND VPWR VPWR _0248_ sky130_fd_sc_hd__mux4_1
X_2161_ net753 VGND VGND VPWR VPWR net216 sky130_fd_sc_hd__buf_1
X_2092_ net778 net743 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame0_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1043_ net61 net89 net25 net117 Inst_LUT4AB_ConfigMem.Inst_frame5_bit9.Q Inst_LUT4AB_ConfigMem.Inst_frame5_bit8.Q
+ VGND VGND VPWR VPWR _0183_ sky130_fd_sc_hd__mux4_2
XFILLER_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1945_ net754 net56 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_16_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1876_ net789 net680 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame6_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0758_ _0554_ _0605_ _0607_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit6.Q VGND VGND VPWR
+ VPWR _0608_ sky130_fd_sc_hd__o211a_1
X_0827_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit8.Q _0671_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit9.Q
+ VGND VGND VPWR VPWR _0672_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_67_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_73_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1661_ net810 net727 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame13_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1730_ net800 net737 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame11_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1592_ net756 net717 VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_7_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2144_ EE4END[9] VGND VGND VPWR VPWR net183 sky130_fd_sc_hd__clkbuf_1
XFILLER_38_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2213_ Inst_LUT4AB_switch_matrix.JN2BEG2 VGND VGND VPWR VPWR net246 sky130_fd_sc_hd__buf_8
XFILLER_53_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1026_ net20 net131 net103 Inst_LUT4AB_switch_matrix.JN2BEG4 Inst_LUT4AB_ConfigMem.Inst_frame7_bit3.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame7_bit2.Q VGND VGND VPWR VPWR _0167_ sky130_fd_sc_hd__mux4_1
XFILLER_38_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2075_ net749 net744 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame0_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1928_ net41 net686 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame5_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1859_ net797 net675 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame7_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_12_Left_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_70_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold91 Inst_LE_LUT4c_frame_config_dffesr.LUT_flop VGND VGND VPWR VPWR net483 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_43_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1713_ net763 net731 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame12_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_16_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1575_ net787 net714 VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.c_out_mux
+ sky130_fd_sc_hd__dlxtp_1
X_1644_ net778 net721 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame14_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2127_ E6END[2] VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__clkbuf_1
Xrebuffer12 net425 VGND VGND VPWR VPWR net404 sky130_fd_sc_hd__buf_6
Xrebuffer23 net414 VGND VGND VPWR VPWR net415 sky130_fd_sc_hd__buf_6
XFILLER_58_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer56 net449 VGND VGND VPWR VPWR net448 sky130_fd_sc_hd__buf_6
X_1009_ net643 net633 net628 net415 Inst_LUT4AB_ConfigMem.Inst_frame4_bit2.Q Inst_LUT4AB_ConfigMem.Inst_frame4_bit3.Q
+ VGND VGND VPWR VPWR _0152_ sky130_fd_sc_hd__mux4_2
X_2058_ net781 net702 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_24_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1360_ net413 net410 net397 net432 Inst_LUT4AB_ConfigMem.Inst_frame12_bit6.Q Inst_LUT4AB_ConfigMem.Inst_frame12_bit7.Q
+ VGND VGND VPWR VPWR _0468_ sky130_fd_sc_hd__mux4_1
X_1291_ net654 net411 net649 net645 Inst_LUT4AB_ConfigMem.Inst_frame4_bit27.Q Inst_LUT4AB_ConfigMem.Inst_frame4_bit26.Q
+ VGND VGND VPWR VPWR _0411_ sky130_fd_sc_hd__mux4_1
XFILLER_63_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1627_ net749 net724 VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11
+ sky130_fd_sc_hd__dlxtp_1
X_1558_ net760 net715 VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.c_reset_value
+ sky130_fd_sc_hd__dlxtp_1
X_1489_ net763 net55 VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_14_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_210 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_235 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0791_ _0637_ _0638_ _0550_ _0634_ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.JN2BEG1
+ sky130_fd_sc_hd__o2bb2a_4
X_0860_ Inst_LB_LUT4c_frame_config_dffesr.c_I0mux _0010_ VGND VGND VPWR VPWR _0013_
+ sky130_fd_sc_hd__and2b_1
XFILLER_68_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1343_ _0454_ _0453_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit5.Q VGND VGND VPWR VPWR
+ Inst_LUT4AB_switch_matrix.SS4BEG3 sky130_fd_sc_hd__mux2_4
XFILLER_5_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1412_ net90 net105 net133 net635 Inst_LUT4AB_ConfigMem.Inst_frame12_bit24.Q Inst_LUT4AB_ConfigMem.Inst_frame12_bit25.Q
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.S4BEG3 sky130_fd_sc_hd__mux4_1
X_1274_ net660 net656 net407 VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.M_AB sky130_fd_sc_hd__mux2_4
XFILLER_51_246 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0989_ net85 net87 net95 net666 Inst_LUT4AB_ConfigMem.Inst_frame1_bit14.Q Inst_LUT4AB_ConfigMem.Inst_frame1_bit15.Q
+ VGND VGND VPWR VPWR _0134_ sky130_fd_sc_hd__mux4_1
XFILLER_3_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_0_Left_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout690 net56 VGND VGND VPWR VPWR net690 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_5_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1961_ net783 net689 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0912_ _0058_ _0056_ _0061_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit5.Q VGND VGND VPWR
+ VPWR Inst_LUT4AB_switch_matrix.JS2BEG2 sky130_fd_sc_hd__o22a_4
X_1892_ net796 net680 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame6_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0774_ _0621_ _0622_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit8.Q VGND VGND VPWR VPWR
+ _0623_ sky130_fd_sc_hd__mux2_4
X_0843_ Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10
+ _0643_ VGND VGND VPWR VPWR _0686_ sky130_fd_sc_hd__mux2_1
X_1326_ net58 net86 net114 net411 Inst_LUT4AB_ConfigMem.Inst_frame11_bit23.Q Inst_LUT4AB_ConfigMem.Inst_frame11_bit24.Q
+ VGND VGND VPWR VPWR _0442_ sky130_fd_sc_hd__mux4_1
X_1188_ Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 _0303_ VGND VGND
+ VPWR VPWR _0320_ sky130_fd_sc_hd__or2_1
X_1257_ net57 net61 net2 net6 Inst_LUT4AB_ConfigMem.Inst_frame2_bit22.Q Inst_LUT4AB_ConfigMem.Inst_frame2_bit23.Q
+ VGND VGND VPWR VPWR _0382_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_54_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput282 Inst_LUT4AB_switch_matrix.NN4BEG3 VGND VGND VPWR VPWR NN4BEG[15] sky130_fd_sc_hd__buf_8
Xoutput271 net271 VGND VGND VPWR VPWR N4BEG[5] sky130_fd_sc_hd__buf_2
Xoutput260 net260 VGND VGND VPWR VPWR N4BEG[0] sky130_fd_sc_hd__buf_2
Xoutput293 Inst_LUT4AB_switch_matrix.S1BEG1 VGND VGND VPWR VPWR S1BEG[1] sky130_fd_sc_hd__buf_6
XPHY_EDGE_ROW_27_Left_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_36_Left_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2160_ net756 VGND VGND VPWR VPWR net215 sky130_fd_sc_hd__clkbuf_1
XFILLER_65_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1111_ _0245_ _0246_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit20.Q VGND VGND VPWR VPWR
+ _0247_ sky130_fd_sc_hd__mux2_2
XFILLER_61_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2091_ net780 net743 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame0_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1042_ net77 net133 net109 Inst_LUT4AB_switch_matrix.JW2BEG2 Inst_LUT4AB_ConfigMem.Inst_frame0_bit9.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame0_bit8.Q VGND VGND VPWR VPWR _0182_ sky130_fd_sc_hd__mux4_2
X_1944_ net756 net690 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1875_ net811 net680 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame6_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0757_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit5.Q _0606_ VGND VGND VPWR VPWR _0607_
+ sky130_fd_sc_hd__or2_1
X_0826_ net93 net121 net105 net137 Inst_LUT4AB_ConfigMem.Inst_frame1_bit7.Q Inst_LUT4AB_ConfigMem.Inst_frame1_bit6.Q
+ VGND VGND VPWR VPWR _0671_ sky130_fd_sc_hd__mux4_1
X_2289_ S4END[14] VGND VGND VPWR VPWR net313 sky130_fd_sc_hd__clkbuf_2
X_1309_ _0426_ _0425_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit0.Q VGND VGND VPWR VPWR
+ _0427_ sky130_fd_sc_hd__mux2_4
X_2358_ Inst_LUT4AB_switch_matrix.WW4BEG2 VGND VGND VPWR VPWR net382 sky130_fd_sc_hd__clkbuf_1
XFILLER_44_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_271 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_92 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1660_ net748 net726 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame13_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_50_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1591_ net758 net717 VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13
+ sky130_fd_sc_hd__dlxtp_1
X_2143_ EE4END[8] VGND VGND VPWR VPWR net182 sky130_fd_sc_hd__clkbuf_1
X_2212_ Inst_LUT4AB_switch_matrix.JN2BEG1 VGND VGND VPWR VPWR net245 sky130_fd_sc_hd__buf_8
X_1025_ _0161_ _0163_ _0166_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit13.Q VGND VGND VPWR
+ VPWR Inst_LUT4AB_switch_matrix.JN2BEG4 sky130_fd_sc_hd__o22a_4
X_2074_ net752 net745 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame0_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_19_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1927_ net40 net686 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame5_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1858_ net800 net677 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame7_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0809_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit0.Q _0654_ VGND VGND VPWR VPWR _0655_
+ sky130_fd_sc_hd__or2_1
X_1789_ net809 net668 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_55_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_70_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold92 Inst_LD_LUT4c_frame_config_dffesr.LUT_flop VGND VGND VPWR VPWR net484 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_43_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1 net141 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1643_ net780 net721 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame14_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1712_ net767 net731 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame12_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1574_ net791 net712 VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer13 net404 VGND VGND VPWR VPWR net405 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer24 Inst_LUT4AB_switch_matrix.M_AH VGND VGND VPWR VPWR net416 sky130_fd_sc_hd__buf_6
XFILLER_54_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer35 net433 VGND VGND VPWR VPWR net427 sky130_fd_sc_hd__buf_6
Xrebuffer57 net450 VGND VGND VPWR VPWR net449 sky130_fd_sc_hd__buf_6
X_2057_ net783 net702 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2126_ net21 VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__buf_1
XFILLER_26_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1008_ net661 net658 net638 net647 Inst_LUT4AB_ConfigMem.Inst_frame4_bit2.Q Inst_LUT4AB_ConfigMem.Inst_frame4_bit3.Q
+ VGND VGND VPWR VPWR _0151_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_32_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1290_ _0407_ _0406_ _0410_ _0590_ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.JS2BEG0
+ sky130_fd_sc_hd__a22o_4
X_1626_ net751 net723 VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10
+ sky130_fd_sc_hd__dlxtp_1
X_1557_ net765 net715 VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.c_I0mux
+ sky130_fd_sc_hd__dlxtp_1
X_1488_ net767 net55 VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_37_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_43_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrebuffer4 _0327_ VGND VGND VPWR VPWR net396 sky130_fd_sc_hd__buf_6
XFILLER_42_70 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0790_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit0.Q _0635_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit1.Q
+ VGND VGND VPWR VPWR _0638_ sky130_fd_sc_hd__a21oi_1
X_1273_ _0395_ _0396_ Inst_LUT4AB_ConfigMem.Inst_frame14_bit17.Q VGND VGND VPWR VPWR
+ Inst_LUT4AB_switch_matrix.M_AH sky130_fd_sc_hd__mux2_4
X_1342_ net58 net3 net114 net635 Inst_LUT4AB_ConfigMem.Inst_frame11_bit3.Q Inst_LUT4AB_ConfigMem.Inst_frame11_bit4.Q
+ VGND VGND VPWR VPWR _0454_ sky130_fd_sc_hd__mux4_1
X_1411_ net639 Inst_LUT4AB_switch_matrix.JS2BEG3 _0192_ _0043_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit7.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame11_bit6.Q VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.W1BEG0
+ sky130_fd_sc_hd__mux4_1
X_0988_ _0131_ _0132_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit16.Q VGND VGND VPWR VPWR
+ _0133_ sky130_fd_sc_hd__mux2_4
X_1609_ net784 net718 VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_67_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout691 net694 VGND VGND VPWR VPWR net691 sky130_fd_sc_hd__clkbuf_2
Xfanout680 FrameStrobe[6] VGND VGND VPWR VPWR net680 sky130_fd_sc_hd__buf_1
XFILLER_18_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1960_ net786 net689 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_33_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0911_ _0060_ _0059_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit4.Q VGND VGND VPWR VPWR
+ _0061_ sky130_fd_sc_hd__mux2_1
X_0842_ Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8
+ _0643_ VGND VGND VPWR VPWR _0685_ sky130_fd_sc_hd__mux2_1
X_1891_ net798 net680 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame6_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_21_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0773_ net640 net630 net625 net622 Inst_LUT4AB_ConfigMem.Inst_frame4_bit6.Q Inst_LUT4AB_ConfigMem.Inst_frame4_bit7.Q
+ VGND VGND VPWR VPWR _0622_ sky130_fd_sc_hd__mux4_1
X_1256_ _0380_ _0379_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit24.Q VGND VGND VPWR VPWR
+ _0381_ sky130_fd_sc_hd__mux2_4
XFILLER_56_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1325_ _0438_ _0441_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit29.Q VGND VGND VPWR VPWR
+ Inst_LUT4AB_switch_matrix.W6BEG0 sky130_fd_sc_hd__mux2_4
X_1187_ Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 _0307_ _0308_ Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11
+ VGND VGND VPWR VPWR _0319_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_19_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput283 net283 VGND VGND VPWR VPWR NN4BEG[1] sky130_fd_sc_hd__buf_2
Xoutput250 net250 VGND VGND VPWR VPWR N2BEG[6] sky130_fd_sc_hd__buf_6
Xoutput261 net261 VGND VGND VPWR VPWR N4BEG[10] sky130_fd_sc_hd__buf_2
Xoutput272 net272 VGND VGND VPWR VPWR N4BEG[6] sky130_fd_sc_hd__buf_2
XFILLER_59_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput294 Inst_LUT4AB_switch_matrix.S1BEG2 VGND VGND VPWR VPWR S1BEG[2] sky130_fd_sc_hd__buf_6
XFILLER_62_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_2_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1110_ net646 net627 net642 net623 Inst_LUT4AB_ConfigMem.Inst_frame2_bit19.Q Inst_LUT4AB_ConfigMem.Inst_frame2_bit18.Q
+ VGND VGND VPWR VPWR _0246_ sky130_fd_sc_hd__mux4_1
XFILLER_38_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2090_ net781 net746 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame0_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_31_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1041_ _0177_ _0178_ _0181_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit5.Q VGND VGND VPWR
+ VPWR Inst_LUT4AB_switch_matrix.JW2BEG2 sky130_fd_sc_hd__o22a_4
X_1943_ net758 net690 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1874_ net762 net676 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame7_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0825_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit8.Q _0669_ VGND VGND VPWR VPWR _0670_
+ sky130_fd_sc_hd__and2b_1
Xclkbuf_0_UserCLK UserCLK VGND VGND VPWR VPWR clknet_0_UserCLK sky130_fd_sc_hd__clkbuf_16
X_0756_ net81 net91 net8 net119 Inst_LUT4AB_ConfigMem.Inst_frame6_bit29.Q Inst_LUT4AB_ConfigMem.Inst_frame6_bit28.Q
+ VGND VGND VPWR VPWR _0606_ sky130_fd_sc_hd__mux4_2
X_2288_ S4END[13] VGND VGND VPWR VPWR net327 sky130_fd_sc_hd__clkbuf_2
X_1239_ _0364_ _0365_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit24.Q VGND VGND VPWR VPWR
+ _0366_ sky130_fd_sc_hd__mux2_1
X_1308_ net631 net627 net397 net432 Inst_LUT4AB_ConfigMem.Inst_frame11_bit30.Q Inst_LUT4AB_ConfigMem.Inst_frame11_bit31.Q
+ VGND VGND VPWR VPWR _0426_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_50_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_71 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1590_ net760 net717 VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12
+ sky130_fd_sc_hd__dlxtp_1
X_1024_ _0164_ _0165_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit12.Q VGND VGND VPWR VPWR
+ _0166_ sky130_fd_sc_hd__mux2_1
X_2142_ EE4END[7] VGND VGND VPWR VPWR net181 sky130_fd_sc_hd__clkbuf_1
X_2073_ net754 net745 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame0_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_26_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2211_ Inst_LUT4AB_switch_matrix.JN2BEG0 VGND VGND VPWR VPWR net244 sky130_fd_sc_hd__buf_4
X_1926_ net792 net685 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame5_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1788_ net747 net669 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1857_ net802 net677 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame7_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0808_ net426 net634 net649 net644 Inst_LUT4AB_ConfigMem.Inst_frame3_bit31.Q Inst_LUT4AB_ConfigMem.Inst_frame3_bit30.Q
+ VGND VGND VPWR VPWR _0654_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_55_Left_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0739_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit29.Q VGND VGND VPWR VPWR _0590_ sky130_fd_sc_hd__inv_1
XPHY_EDGE_ROW_64_Left_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_73_Left_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold93 Inst_LH_LUT4c_frame_config_dffesr.LUT_flop VGND VGND VPWR VPWR net485 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_43_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_180 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_2 net152 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1642_ net781 net721 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame14_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_31_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1711_ net769 net734 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame12_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1573_ net793 net712 VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14
+ sky130_fd_sc_hd__dlxtp_1
Xrebuffer25 _0395_ VGND VGND VPWR VPWR net417 sky130_fd_sc_hd__buf_6
X_2056_ net786 net701 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_66_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrebuffer36 _0352_ VGND VGND VPWR VPWR net428 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer58 net451 VGND VGND VPWR VPWR net450 sky130_fd_sc_hd__buf_6
X_2125_ net20 VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__buf_1
Xrebuffer14 net446 VGND VGND VPWR VPWR net406 sky130_fd_sc_hd__buf_6
X_1007_ _0150_ Inst_LE_LUT4c_frame_config_dffesr.LUT_flop Inst_LE_LUT4c_frame_config_dffesr.c_out_mux
+ VGND VGND VPWR VPWR E sky130_fd_sc_hd__mux2_4
XFILLER_41_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1909_ net765 net686 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame5_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_32_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1625_ net753 net723 VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9
+ sky130_fd_sc_hd__dlxtp_1
X_1556_ net789 net715 VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.c_out_mux
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_54_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1487_ net769 net55 VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4
+ sky130_fd_sc_hd__dlxtp_1
X_2039_ net757 net700 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2108_ Inst_LUT4AB_switch_matrix.E1BEG1 VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__buf_4
XFILLER_10_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_43_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1410_ net629 _0093_ Inst_LUT4AB_switch_matrix.JS2BEG0 _0098_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit8.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame11_bit9.Q VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.W1BEG1
+ sky130_fd_sc_hd__mux4_2
X_1272_ _0355_ _0394_ _0390_ VGND VGND VPWR VPWR _0396_ sky130_fd_sc_hd__mux2_4
XFILLER_68_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1341_ net648 net431 _0252_ _0683_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit3.Q Inst_LUT4AB_ConfigMem.Inst_frame11_bit4.Q
+ VGND VGND VPWR VPWR _0453_ sky130_fd_sc_hd__mux4_1
X_0987_ net647 net632 net628 net398 Inst_LUT4AB_ConfigMem.Inst_frame1_bit14.Q Inst_LUT4AB_ConfigMem.Inst_frame1_bit15.Q
+ VGND VGND VPWR VPWR _0132_ sky130_fd_sc_hd__mux4_2
XFILLER_59_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1608_ net785 net718 VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11
+ sky130_fd_sc_hd__dlxtp_1
X_1539_ net798 net711 VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.c_reset_value
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_27_267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout692 net693 VGND VGND VPWR VPWR net692 sky130_fd_sc_hd__clkbuf_2
Xfanout670 FrameStrobe[9] VGND VGND VPWR VPWR net670 sky130_fd_sc_hd__buf_2
Xfanout681 net682 VGND VGND VPWR VPWR net681 sky130_fd_sc_hd__clkbuf_2
XFILLER_2_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_5_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1890_ net34 net681 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame6_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0910_ net84 net3 net9 net813 Inst_LUT4AB_ConfigMem.Inst_frame2_bit2.Q Inst_LUT4AB_ConfigMem.Inst_frame2_bit3.Q
+ VGND VGND VPWR VPWR _0060_ sky130_fd_sc_hd__mux4_1
X_0772_ net659 net655 net650 net645 Inst_LUT4AB_ConfigMem.Inst_frame4_bit6.Q Inst_LUT4AB_ConfigMem.Inst_frame4_bit7.Q
+ VGND VGND VPWR VPWR _0621_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0841_ _0673_ _0674_ _0683_ _0682_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit9.Q Inst_LUT4AB_ConfigMem.Inst_frame10_bit10.Q
+ VGND VGND VPWR VPWR _0684_ sky130_fd_sc_hd__mux4_2
XFILLER_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1186_ Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 _0304_ _0316_ _0317_
+ VGND VGND VPWR VPWR _0318_ sky130_fd_sc_hd__o211a_1
X_1255_ net660 net657 net652 net637 Inst_LUT4AB_ConfigMem.Inst_frame2_bit22.Q Inst_LUT4AB_ConfigMem.Inst_frame2_bit23.Q
+ VGND VGND VPWR VPWR _0380_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_34_Right_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1324_ _0440_ _0439_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit28.Q VGND VGND VPWR VPWR
+ _0441_ sky130_fd_sc_hd__mux2_4
XPHY_EDGE_ROW_43_Right_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput284 net284 VGND VGND VPWR VPWR NN4BEG[2] sky130_fd_sc_hd__buf_2
Xoutput262 net262 VGND VGND VPWR VPWR N4BEG[11] sky130_fd_sc_hd__buf_2
Xoutput251 net251 VGND VGND VPWR VPWR N2BEG[7] sky130_fd_sc_hd__buf_2
Xoutput240 net240 VGND VGND VPWR VPWR N1BEG[0] sky130_fd_sc_hd__clkbuf_4
Xoutput273 net273 VGND VGND VPWR VPWR N4BEG[7] sky130_fd_sc_hd__buf_2
XFILLER_59_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_52_Right_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput295 Inst_LUT4AB_switch_matrix.S1BEG3 VGND VGND VPWR VPWR S1BEG[3] sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_53_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_61_Right_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_70_Right_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_70 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1040_ _0180_ _0179_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit4.Q VGND VGND VPWR VPWR
+ _0181_ sky130_fd_sc_hd__mux2_1
XFILLER_64_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1942_ net759 net690 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1873_ net46 net676 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame7_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0824_ net59 net10 net65 net814 Inst_LUT4AB_ConfigMem.Inst_frame1_bit7.Q Inst_LUT4AB_ConfigMem.Inst_frame1_bit6.Q
+ VGND VGND VPWR VPWR _0669_ sky130_fd_sc_hd__mux4_1
X_0755_ net26 net107 net124 Inst_LUT4AB_switch_matrix.E2BEG1 Inst_LUT4AB_ConfigMem.Inst_frame1_bit28.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame1_bit29.Q VGND VGND VPWR VPWR _0605_ sky130_fd_sc_hd__mux4_1
X_2356_ Inst_LUT4AB_switch_matrix.WW4BEG0 VGND VGND VPWR VPWR net380 sky130_fd_sc_hd__clkbuf_2
XFILLER_28_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2287_ S4END[12] VGND VGND VPWR VPWR net326 sky130_fd_sc_hd__clkbuf_2
X_1169_ _0252_ _0253_ _0244_ _0243_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit13.Q Inst_LUT4AB_ConfigMem.Inst_frame8_bit14.Q
+ VGND VGND VPWR VPWR _0301_ sky130_fd_sc_hd__mux4_2
X_1238_ net646 net631 net641 net432 Inst_LUT4AB_ConfigMem.Inst_frame4_bit23.Q Inst_LUT4AB_ConfigMem.Inst_frame4_bit22.Q
+ VGND VGND VPWR VPWR _0365_ sky130_fd_sc_hd__mux4_1
XFILLER_52_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1307_ _0652_ _0071_ _0107_ _0252_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit30.Q Inst_LUT4AB_ConfigMem.Inst_frame11_bit31.Q
+ VGND VGND VPWR VPWR _0425_ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_50_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2210_ Inst_LUT4AB_switch_matrix.N1BEG3 VGND VGND VPWR VPWR net243 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_64_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1023_ net86 net94 net114 net665 Inst_LUT4AB_ConfigMem.Inst_frame4_bit10.Q Inst_LUT4AB_ConfigMem.Inst_frame4_bit11.Q
+ VGND VGND VPWR VPWR _0165_ sky130_fd_sc_hd__mux4_1
X_2141_ EE4END[6] VGND VGND VPWR VPWR net180 sky130_fd_sc_hd__clkbuf_1
X_2072_ net755 net743 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame0_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1925_ net794 net685 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame5_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_34_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1856_ net803 net676 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame7_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0807_ net74 net19 net102 net130 Inst_LUT4AB_ConfigMem.Inst_frame7_bit30.Q Inst_LUT4AB_ConfigMem.Inst_frame7_bit31.Q
+ VGND VGND VPWR VPWR _0653_ sky130_fd_sc_hd__mux4_2
X_1787_ net749 net670 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0738_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit28.Q VGND VGND VPWR VPWR _0589_ sky130_fd_sc_hd__inv_1
XFILLER_69_284 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2339_ W6END[9] VGND VGND VPWR VPWR net374 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold94 Inst_LC_LUT4c_frame_config_dffesr.LUT_flop VGND VGND VPWR VPWR net486 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_16_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1572_ net796 net712 VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13
+ sky130_fd_sc_hd__dlxtp_1
XANTENNA_3 net155 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1710_ net771 net731 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame12_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1641_ net783 net721 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame14_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2124_ net19 VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__clkbuf_1
X_2055_ net788 net701 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
Xrebuffer59 net452 VGND VGND VPWR VPWR net451 sky130_fd_sc_hd__buf_6
Xrebuffer37 Inst_LUT4AB_switch_matrix.JW2BEG5 VGND VGND VPWR VPWR net429 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer15 _0327_ VGND VGND VPWR VPWR net407 sky130_fd_sc_hd__buf_6
X_1006_ _0149_ _0144_ _0140_ VGND VGND VPWR VPWR _0150_ sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_32_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1908_ net790 net684 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame5_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1839_ net769 net674 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame8_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_1_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1624_ net756 net723 VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8
+ sky130_fd_sc_hd__dlxtp_1
X_1555_ net811 net715 VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_27_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1486_ net771 net55 VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3
+ sky130_fd_sc_hd__dlxtp_1
X_2038_ net759 net699 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_6_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_43_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1340_ _0595_ _0448_ _0452_ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.WW4BEG0
+ sky130_fd_sc_hd__o21a_1
X_1271_ _0393_ _0394_ Inst_LUT4AB_ConfigMem.Inst_frame14_bit16.Q VGND VGND VPWR VPWR
+ _0395_ sky130_fd_sc_hd__mux2_4
X_0986_ net660 net656 net652 net636 Inst_LUT4AB_ConfigMem.Inst_frame1_bit14.Q Inst_LUT4AB_ConfigMem.Inst_frame1_bit15.Q
+ VGND VGND VPWR VPWR _0131_ sky130_fd_sc_hd__mux4_1
X_1607_ net787 net718 VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_59_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1469_ net484 Inst_LUT4AB_ConfigMem.Inst_frame9_bit0.Q net467 _0536_ _0537_ VGND
+ VGND VPWR VPWR _0004_ sky130_fd_sc_hd__a32o_1
X_1538_ net799 net708 VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.c_I0mux
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_67_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_19_Left_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout671 net672 VGND VGND VPWR VPWR net671 sky130_fd_sc_hd__clkbuf_2
Xfanout660 net662 VGND VGND VPWR VPWR net660 sky130_fd_sc_hd__buf_2
Xfanout693 net694 VGND VGND VPWR VPWR net693 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_5_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout682 FrameStrobe[6] VGND VGND VPWR VPWR net682 sky130_fd_sc_hd__clkbuf_4
XFILLER_73_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_56_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0840_ net61 net89 net6 net138 Inst_LUT4AB_ConfigMem.Inst_frame5_bit1.Q Inst_LUT4AB_ConfigMem.Inst_frame5_bit0.Q
+ VGND VGND VPWR VPWR _0683_ sky130_fd_sc_hd__mux4_2
X_0771_ _0608_ _0619_ VGND VGND VPWR VPWR _0620_ sky130_fd_sc_hd__nor2_1
XFILLER_68_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1323_ net399 net625 net623 net406 Inst_LUT4AB_ConfigMem.Inst_frame11_bit26.Q Inst_LUT4AB_ConfigMem.Inst_frame11_bit27.Q
+ VGND VGND VPWR VPWR _0440_ sky130_fd_sc_hd__mux4_2
XFILLER_5_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1185_ Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 _0308_ VGND VGND
+ VPWR VPWR _0317_ sky130_fd_sc_hd__or2_1
X_1254_ net646 net631 net641 Inst_LUT4AB_switch_matrix.M_AD Inst_LUT4AB_ConfigMem.Inst_frame2_bit23.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame2_bit22.Q VGND VGND VPWR VPWR _0379_ sky130_fd_sc_hd__mux4_2
XFILLER_24_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_238 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput241 net241 VGND VGND VPWR VPWR N1BEG[1] sky130_fd_sc_hd__buf_4
Xoutput230 net230 VGND VGND VPWR VPWR FrameStrobe_O[19] sky130_fd_sc_hd__buf_2
Xoutput252 net252 VGND VGND VPWR VPWR N2BEGb[0] sky130_fd_sc_hd__buf_2
X_0969_ net59 net67 net816 net12 Inst_LUT4AB_ConfigMem.Inst_frame3_bit14.Q Inst_LUT4AB_ConfigMem.Inst_frame3_bit15.Q
+ VGND VGND VPWR VPWR _0115_ sky130_fd_sc_hd__mux4_1
XFILLER_3_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput263 net263 VGND VGND VPWR VPWR N4BEG[12] sky130_fd_sc_hd__buf_4
Xoutput274 net274 VGND VGND VPWR VPWR N4BEG[8] sky130_fd_sc_hd__buf_2
Xoutput285 net285 VGND VGND VPWR VPWR NN4BEG[3] sky130_fd_sc_hd__buf_2
XFILLER_58_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput296 net296 VGND VGND VPWR VPWR S2BEG[0] sky130_fd_sc_hd__buf_8
XFILLER_70_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_190 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_4_Left_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1941_ net765 net690 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1872_ net768 net675 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame7_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0754_ _0601_ _0599_ _0604_ _0556_ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.E2BEG1
+ sky130_fd_sc_hd__a22o_1
X_0823_ _0666_ _0667_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit8.Q VGND VGND VPWR VPWR
+ _0668_ sky130_fd_sc_hd__mux2_4
X_2286_ S4END[11] VGND VGND VPWR VPWR net325 sky130_fd_sc_hd__clkbuf_2
XFILLER_56_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1306_ _0419_ _0421_ _0424_ _0594_ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.JN2BEG0
+ sky130_fd_sc_hd__a22o_1
X_2355_ WW4END[15] VGND VGND VPWR VPWR net379 sky130_fd_sc_hd__clkbuf_2
X_1099_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit20.Q _0233_ _0235_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit21.Q
+ VGND VGND VPWR VPWR _0236_ sky130_fd_sc_hd__a211o_1
X_1168_ _0294_ _0267_ Inst_LH_LUT4c_frame_config_dffesr.c_I0mux _0299_ VGND VGND VPWR
+ VPWR _0300_ sky130_fd_sc_hd__a31o_1
X_1237_ net662 net656 net652 net636 Inst_LUT4AB_ConfigMem.Inst_frame4_bit22.Q Inst_LUT4AB_ConfigMem.Inst_frame4_bit23.Q
+ VGND VGND VPWR VPWR _0364_ sky130_fd_sc_hd__mux4_1
XFILLER_44_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2140_ EE4END[5] VGND VGND VPWR VPWR net179 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_64_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1022_ net58 net66 net3 net11 Inst_LUT4AB_ConfigMem.Inst_frame4_bit10.Q Inst_LUT4AB_ConfigMem.Inst_frame4_bit11.Q
+ VGND VGND VPWR VPWR _0164_ sky130_fd_sc_hd__mux4_1
XFILLER_38_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2071_ net757 net743 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame0_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_19_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1855_ net805 net676 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame7_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1924_ net795 net683 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame5_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1786_ net751 net670 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0806_ net73 net18 net129 Inst_LUT4AB_switch_matrix.JS2BEG3 Inst_LUT4AB_ConfigMem.Inst_frame8_bit30.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame8_bit31.Q VGND VGND VPWR VPWR _0652_ sky130_fd_sc_hd__mux4_2
X_0737_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit29.Q VGND VGND VPWR VPWR _0588_ sky130_fd_sc_hd__inv_1
XFILLER_72_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2269_ Inst_LUT4AB_switch_matrix.JS2BEG6 VGND VGND VPWR VPWR net302 sky130_fd_sc_hd__buf_4
X_2338_ W6END[8] VGND VGND VPWR VPWR net373 sky130_fd_sc_hd__clkbuf_2
XFILLER_40_325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold95 Inst_LB_LUT4c_frame_config_dffesr.LUT_flop VGND VGND VPWR VPWR net487 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_16_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_7_Left_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1571_ net798 net713 VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12
+ sky130_fd_sc_hd__dlxtp_1
XANTENNA_4 net156 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1640_ net786 net721 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame14_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
Xrebuffer16 Inst_LUT4AB_switch_matrix.JS2BEG5 VGND VGND VPWR VPWR net408 sky130_fd_sc_hd__clkbuf_2
X_2123_ net18 VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__clkbuf_2
X_2054_ net792 net701 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1005_ _0146_ _0148_ _0097_ VGND VGND VPWR VPWR _0149_ sky130_fd_sc_hd__mux2_1
XFILLER_22_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1838_ net771 net674 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame8_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1907_ net812 net684 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame5_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_66_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1769_ net784 net739 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame10_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_23_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput130 W2MID[5] VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__clkbuf_2
XFILLER_72_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1623_ net758 net723 VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7
+ sky130_fd_sc_hd__dlxtp_1
X_1554_ net762 net710 VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14
+ sky130_fd_sc_hd__dlxtp_1
X_1485_ net774 net55 VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2
+ sky130_fd_sc_hd__dlxtp_1
.ends

