module N_IO (A_I_top,
    A_O_top,
    A_T_top,
    A_config_C_bit0,
    A_config_C_bit1,
    A_config_C_bit2,
    A_config_C_bit3,
    B_I_top,
    B_O_top,
    B_T_top,
    B_config_C_bit0,
    B_config_C_bit1,
    B_config_C_bit2,
    B_config_C_bit3,
    Ci,
    UserCLK,
    UserCLKo,
    VPWR,
    VGND,
    FrameData,
    FrameData_O,
    FrameStrobe,
    FrameStrobe_O,
    N1END,
    N2END,
    N2MID,
    N4END,
    NN4END,
    S1BEG,
    S2BEG,
    S2BEGb,
    S4BEG,
    SS4BEG);
 output A_I_top;
 input A_O_top;
 output A_T_top;
 output A_config_C_bit0;
 output A_config_C_bit1;
 output A_config_C_bit2;
 output A_config_C_bit3;
 output B_I_top;
 input B_O_top;
 output B_T_top;
 output B_config_C_bit0;
 output B_config_C_bit1;
 output B_config_C_bit2;
 output B_config_C_bit3;
 input Ci;
 input UserCLK;
 output UserCLKo;
 inout VPWR;
 inout VGND;
 input [31:0] FrameData;
 output [31:0] FrameData_O;
 input [19:0] FrameStrobe;
 output [19:0] FrameStrobe_O;
 input [3:0] N1END;
 input [7:0] N2END;
 input [7:0] N2MID;
 input [15:0] N4END;
 input [15:0] NN4END;
 output [3:0] S1BEG;
 output [7:0] S2BEG;
 output [7:0] S2BEGb;
 output [15:0] S4BEG;
 output [15:0] SS4BEG;

 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire \Inst_A_IO_1_bidirectional_frame_config_pass.Q ;
 wire \Inst_B_IO_1_bidirectional_frame_config_pass.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame0_bit0.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame0_bit1.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame0_bit10.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame0_bit11.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame0_bit12.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame0_bit13.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame0_bit14.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame0_bit15.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame0_bit16.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame0_bit17.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame0_bit18.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame0_bit19.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame0_bit2.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame0_bit20.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame0_bit21.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame0_bit22.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame0_bit23.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame0_bit24.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame0_bit25.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame0_bit26.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame0_bit27.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame0_bit28.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame0_bit29.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame0_bit3.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame0_bit30.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame0_bit31.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame0_bit4.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame0_bit5.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame0_bit6.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame0_bit7.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame0_bit8.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame0_bit9.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame1_bit0.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame1_bit1.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame1_bit10.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame1_bit11.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame1_bit12.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame1_bit13.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame1_bit14.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame1_bit15.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame1_bit16.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame1_bit17.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame1_bit18.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame1_bit19.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame1_bit2.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame1_bit20.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame1_bit21.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame1_bit22.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame1_bit23.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame1_bit24.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame1_bit25.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame1_bit26.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame1_bit27.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame1_bit28.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame1_bit29.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame1_bit3.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame1_bit30.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame1_bit31.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame1_bit4.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame1_bit5.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame1_bit6.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame1_bit7.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame1_bit8.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame1_bit9.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame2_bit0.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame2_bit1.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame2_bit10.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame2_bit11.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame2_bit12.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame2_bit13.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame2_bit14.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame2_bit15.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame2_bit16.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame2_bit17.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame2_bit18.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame2_bit19.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame2_bit2.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame2_bit20.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame2_bit21.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame2_bit22.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame2_bit23.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame2_bit24.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame2_bit25.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame2_bit26.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame2_bit27.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame2_bit28.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame2_bit29.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame2_bit3.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame2_bit30.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame2_bit31.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame2_bit4.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame2_bit5.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame2_bit6.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame2_bit7.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame2_bit8.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame2_bit9.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame3_bit14.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame3_bit15.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame3_bit16.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame3_bit17.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame3_bit18.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame3_bit19.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame3_bit20.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame3_bit21.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame3_bit22.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame3_bit23.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame3_bit24.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame3_bit25.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame3_bit26.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame3_bit27.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame3_bit28.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame3_bit29.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame3_bit30.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame3_bit31.Q ;
 wire \Inst_N_IO_switch_matrix.S1BEG0 ;
 wire \Inst_N_IO_switch_matrix.S1BEG1 ;
 wire \Inst_N_IO_switch_matrix.S1BEG2 ;
 wire \Inst_N_IO_switch_matrix.S1BEG3 ;
 wire \Inst_N_IO_switch_matrix.S2BEG0 ;
 wire \Inst_N_IO_switch_matrix.S2BEG1 ;
 wire \Inst_N_IO_switch_matrix.S2BEG2 ;
 wire \Inst_N_IO_switch_matrix.S2BEG3 ;
 wire \Inst_N_IO_switch_matrix.S2BEG4 ;
 wire \Inst_N_IO_switch_matrix.S2BEG5 ;
 wire \Inst_N_IO_switch_matrix.S2BEG6 ;
 wire \Inst_N_IO_switch_matrix.S2BEG7 ;
 wire \Inst_N_IO_switch_matrix.S2BEGb0 ;
 wire \Inst_N_IO_switch_matrix.S2BEGb1 ;
 wire \Inst_N_IO_switch_matrix.S2BEGb2 ;
 wire \Inst_N_IO_switch_matrix.S2BEGb3 ;
 wire \Inst_N_IO_switch_matrix.S2BEGb4 ;
 wire \Inst_N_IO_switch_matrix.S2BEGb5 ;
 wire \Inst_N_IO_switch_matrix.S2BEGb6 ;
 wire \Inst_N_IO_switch_matrix.S2BEGb7 ;
 wire \Inst_N_IO_switch_matrix.S4BEG0 ;
 wire \Inst_N_IO_switch_matrix.S4BEG1 ;
 wire \Inst_N_IO_switch_matrix.S4BEG10 ;
 wire \Inst_N_IO_switch_matrix.S4BEG11 ;
 wire \Inst_N_IO_switch_matrix.S4BEG12 ;
 wire \Inst_N_IO_switch_matrix.S4BEG13 ;
 wire \Inst_N_IO_switch_matrix.S4BEG14 ;
 wire \Inst_N_IO_switch_matrix.S4BEG15 ;
 wire \Inst_N_IO_switch_matrix.S4BEG2 ;
 wire \Inst_N_IO_switch_matrix.S4BEG3 ;
 wire \Inst_N_IO_switch_matrix.S4BEG4 ;
 wire \Inst_N_IO_switch_matrix.S4BEG5 ;
 wire \Inst_N_IO_switch_matrix.S4BEG6 ;
 wire \Inst_N_IO_switch_matrix.S4BEG7 ;
 wire \Inst_N_IO_switch_matrix.S4BEG8 ;
 wire \Inst_N_IO_switch_matrix.S4BEG9 ;
 wire \Inst_N_IO_switch_matrix.SS4BEG0 ;
 wire \Inst_N_IO_switch_matrix.SS4BEG1 ;
 wire \Inst_N_IO_switch_matrix.SS4BEG10 ;
 wire \Inst_N_IO_switch_matrix.SS4BEG11 ;
 wire \Inst_N_IO_switch_matrix.SS4BEG12 ;
 wire \Inst_N_IO_switch_matrix.SS4BEG13 ;
 wire \Inst_N_IO_switch_matrix.SS4BEG14 ;
 wire \Inst_N_IO_switch_matrix.SS4BEG15 ;
 wire \Inst_N_IO_switch_matrix.SS4BEG2 ;
 wire \Inst_N_IO_switch_matrix.SS4BEG3 ;
 wire \Inst_N_IO_switch_matrix.SS4BEG4 ;
 wire \Inst_N_IO_switch_matrix.SS4BEG5 ;
 wire \Inst_N_IO_switch_matrix.SS4BEG6 ;
 wire \Inst_N_IO_switch_matrix.SS4BEG7 ;
 wire \Inst_N_IO_switch_matrix.SS4BEG8 ;
 wire \Inst_N_IO_switch_matrix.SS4BEG9 ;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire net229;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net228;

 sg13g2_mux4_1 _049_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame2_bit23.Q ),
    .A0(net58),
    .A1(net101),
    .A2(net97),
    .A3(net1),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame2_bit22.Q ),
    .X(\Inst_N_IO_switch_matrix.S4BEG2 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _050_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame2_bit20.Q ),
    .A0(net39),
    .A1(net61),
    .A2(net100),
    .A3(net2),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame2_bit21.Q ),
    .X(\Inst_N_IO_switch_matrix.S4BEG1 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _051_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame2_bit18.Q ),
    .A0(net38),
    .A1(net62),
    .A2(net101),
    .A3(net1),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame2_bit19.Q ),
    .X(\Inst_N_IO_switch_matrix.S4BEG0 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _052_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame2_bit16.Q ),
    .A0(net40),
    .A1(net56),
    .A2(net95),
    .A3(net109),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame2_bit17.Q ),
    .X(\Inst_N_IO_switch_matrix.S2BEGb7 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _053_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame2_bit14.Q ),
    .A0(net41),
    .A1(net63),
    .A2(net102),
    .A3(net110),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame2_bit15.Q ),
    .X(\Inst_N_IO_switch_matrix.S2BEGb6 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _054_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame2_bit12.Q ),
    .A0(net42),
    .A1(net64),
    .A2(net103),
    .A3(net96),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame2_bit13.Q ),
    .X(\Inst_N_IO_switch_matrix.S2BEGb5 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _055_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame2_bit10.Q ),
    .A0(net43),
    .A1(net65),
    .A2(net104),
    .A3(net97),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame2_bit11.Q ),
    .X(\Inst_N_IO_switch_matrix.S2BEGb4 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _056_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame2_bit8.Q ),
    .A0(net44),
    .A1(net66),
    .A2(net105),
    .A3(net98),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame2_bit9.Q ),
    .X(\Inst_N_IO_switch_matrix.S2BEGb3 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _057_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame2_bit6.Q ),
    .A0(net45),
    .A1(net67),
    .A2(net106),
    .A3(net99),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame2_bit7.Q ),
    .X(\Inst_N_IO_switch_matrix.S2BEGb2 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _058_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame2_bit4.Q ),
    .A0(net46),
    .A1(net68),
    .A2(net107),
    .A3(net100),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame2_bit5.Q ),
    .X(\Inst_N_IO_switch_matrix.S2BEGb1 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _059_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame2_bit2.Q ),
    .A0(net47),
    .A1(net92),
    .A2(net108),
    .A3(net101),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame2_bit3.Q ),
    .X(\Inst_N_IO_switch_matrix.S2BEGb0 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _060_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame2_bit0.Q ),
    .A0(net48),
    .A1(net56),
    .A2(net95),
    .A3(net109),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame2_bit1.Q ),
    .X(\Inst_N_IO_switch_matrix.S2BEG7 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _061_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame3_bit30.Q ),
    .A0(net49),
    .A1(net63),
    .A2(net102),
    .A3(net110),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame3_bit31.Q ),
    .X(\Inst_N_IO_switch_matrix.S2BEG6 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _062_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame3_bit28.Q ),
    .A0(net50),
    .A1(net64),
    .A2(net103),
    .A3(net96),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame3_bit29.Q ),
    .X(\Inst_N_IO_switch_matrix.S2BEG5 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _063_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame3_bit26.Q ),
    .A0(net51),
    .A1(net65),
    .A2(net104),
    .A3(net97),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame3_bit27.Q ),
    .X(\Inst_N_IO_switch_matrix.S2BEG4 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _064_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame3_bit24.Q ),
    .A0(net52),
    .A1(net66),
    .A2(net105),
    .A3(net98),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame3_bit25.Q ),
    .X(\Inst_N_IO_switch_matrix.S2BEG3 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _065_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame3_bit22.Q ),
    .A0(net53),
    .A1(net67),
    .A2(net106),
    .A3(net99),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame3_bit23.Q ),
    .X(\Inst_N_IO_switch_matrix.S2BEG2 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _066_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame3_bit20.Q ),
    .A0(net54),
    .A1(net68),
    .A2(net107),
    .A3(net100),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame3_bit21.Q ),
    .X(\Inst_N_IO_switch_matrix.S2BEG1 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _067_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame3_bit18.Q ),
    .A0(net55),
    .A1(net92),
    .A2(net108),
    .A3(net101),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame3_bit19.Q ),
    .X(\Inst_N_IO_switch_matrix.S2BEG0 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _068_ (.A0(net36),
    .A1(\Inst_B_IO_1_bidirectional_frame_config_pass.Q ),
    .S(\Inst_N_IO_ConfigMem.Inst_frame3_bit17.Q ),
    .X(\Inst_N_IO_switch_matrix.S1BEG3 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _069_ (.A0(net37),
    .A1(net2),
    .S(\Inst_N_IO_ConfigMem.Inst_frame3_bit16.Q ),
    .X(\Inst_N_IO_switch_matrix.S1BEG2 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _070_ (.A0(net38),
    .A1(\Inst_A_IO_1_bidirectional_frame_config_pass.Q ),
    .S(\Inst_N_IO_ConfigMem.Inst_frame3_bit15.Q ),
    .X(\Inst_N_IO_switch_matrix.S1BEG1 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _071_ (.A0(net39),
    .A1(net1),
    .S(\Inst_N_IO_ConfigMem.Inst_frame3_bit14.Q ),
    .X(\Inst_N_IO_switch_matrix.S1BEG0 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _072_ (.Y(_032_),
    .B(\Inst_N_IO_ConfigMem.Inst_frame0_bit24.Q ),
    .A_N(net43),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _073_ (.B1(_032_),
    .VDD(VPWR),
    .Y(_033_),
    .VSS(VGND),
    .A1(net55),
    .A2(\Inst_N_IO_ConfigMem.Inst_frame0_bit24.Q ));
 sg13g2_nand3_1 _074_ (.B(\Inst_N_IO_ConfigMem.Inst_frame0_bit23.Q ),
    .C(_001_),
    .A(net41),
    .Y(_034_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _075_ (.B1(_034_),
    .VDD(VPWR),
    .Y(_035_),
    .VSS(VGND),
    .A1(\Inst_N_IO_ConfigMem.Inst_frame0_bit23.Q ),
    .A2(_033_));
 sg13g2_nand3b_1 _076_ (.B(_001_),
    .C(net40),
    .Y(_036_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(\Inst_N_IO_ConfigMem.Inst_frame0_bit23.Q ));
 sg13g2_o21ai_1 _077_ (.B1(\Inst_N_IO_ConfigMem.Inst_frame0_bit23.Q ),
    .VDD(VPWR),
    .Y(_037_),
    .VSS(VGND),
    .A1(net42),
    .A2(\Inst_N_IO_ConfigMem.Inst_frame0_bit24.Q ));
 sg13g2_nand2_1 _078_ (.Y(_038_),
    .A(net44),
    .B(\Inst_N_IO_ConfigMem.Inst_frame0_bit24.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _079_ (.B(_036_),
    .C(_037_),
    .A(\Inst_N_IO_ConfigMem.Inst_frame0_bit22.Q ),
    .Y(_039_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_038_));
 sg13g2_o21ai_1 _080_ (.B1(_039_),
    .VDD(VPWR),
    .Y(net112),
    .VSS(VGND),
    .A1(\Inst_N_IO_ConfigMem.Inst_frame0_bit22.Q ),
    .A2(_035_));
 sg13g2_nand2b_1 _081_ (.Y(_040_),
    .B(net45),
    .A_N(\Inst_N_IO_ConfigMem.Inst_frame0_bit30.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _082_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame0_bit29.Q ),
    .A0(net54),
    .A1(net55),
    .A2(net40),
    .A3(net44),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame0_bit30.Q ),
    .X(_041_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _083_ (.B1(\Inst_N_IO_ConfigMem.Inst_frame0_bit29.Q ),
    .VDD(VPWR),
    .Y(_042_),
    .VSS(VGND),
    .A1(net46),
    .A2(\Inst_N_IO_ConfigMem.Inst_frame0_bit30.Q ));
 sg13g2_o21ai_1 _084_ (.B1(\Inst_N_IO_ConfigMem.Inst_frame0_bit31.Q ),
    .VDD(VPWR),
    .Y(_043_),
    .VSS(VGND),
    .A1(\Inst_N_IO_ConfigMem.Inst_frame0_bit29.Q ),
    .A2(_040_));
 sg13g2_nand2b_1 _085_ (.Y(_044_),
    .B(_042_),
    .A_N(_043_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _086_ (.B1(_044_),
    .VDD(VPWR),
    .Y(net118),
    .VSS(VGND),
    .A1(\Inst_N_IO_ConfigMem.Inst_frame0_bit31.Q ),
    .A2(_041_));
 sg13g2_inv_1 _087_ (.VDD(VPWR),
    .Y(_000_),
    .A(net41),
    .VSS(VGND));
 sg13g2_inv_1 _088_ (.VDD(VPWR),
    .Y(_001_),
    .A(\Inst_N_IO_ConfigMem.Inst_frame0_bit24.Q ),
    .VSS(VGND));
 sg13g2_mux2_1 _089_ (.A0(net42),
    .A1(net43),
    .S(net69),
    .X(_002_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _090_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_003_),
    .B(net40),
    .A(net69));
 sg13g2_a21oi_1 _091_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net69),
    .A2(_000_),
    .Y(_004_),
    .B1(\Inst_N_IO_ConfigMem.Inst_frame0_bit26.Q ));
 sg13g2_a221oi_1 _092_ (.VSS(VGND),
    .VDD(VPWR),
    .B2(_004_),
    .C1(\Inst_N_IO_ConfigMem.Inst_frame0_bit27.Q ),
    .B1(_003_),
    .A1(\Inst_N_IO_ConfigMem.Inst_frame0_bit26.Q ),
    .Y(_005_),
    .A2(_002_));
 sg13g2_nand2_1 _093_ (.Y(_006_),
    .A(net69),
    .B(net45),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _094_ (.Y(_007_),
    .B(net44),
    .A_N(net69),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _095_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_006_),
    .A2(_007_),
    .Y(_008_),
    .B1(\Inst_N_IO_ConfigMem.Inst_frame0_bit26.Q ));
 sg13g2_nor2b_1 _096_ (.A(net47),
    .B_N(\Inst_N_IO_ConfigMem.Inst_frame0_bit25.Q ),
    .Y(_009_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _097_ (.B1(\Inst_N_IO_ConfigMem.Inst_frame0_bit26.Q ),
    .VDD(VPWR),
    .Y(_010_),
    .VSS(VGND),
    .A1(net69),
    .A2(net46));
 sg13g2_o21ai_1 _098_ (.B1(\Inst_N_IO_ConfigMem.Inst_frame0_bit27.Q ),
    .VDD(VPWR),
    .Y(_011_),
    .VSS(VGND),
    .A1(_009_),
    .A2(_010_));
 sg13g2_o21ai_1 _099_ (.B1(\Inst_N_IO_ConfigMem.Inst_frame0_bit28.Q ),
    .VDD(VPWR),
    .Y(_012_),
    .VSS(VGND),
    .A1(_008_),
    .A2(_011_));
 sg13g2_mux4_1 _100_ (.S0(net69),
    .A0(net52),
    .A1(net53),
    .A2(net54),
    .A3(net55),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame0_bit26.Q ),
    .X(_013_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _101_ (.S0(net69),
    .A0(net48),
    .A1(net49),
    .A2(net50),
    .A3(net51),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame0_bit26.Q ),
    .X(_014_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _102_ (.A0(_014_),
    .A1(_013_),
    .S(\Inst_N_IO_ConfigMem.Inst_frame0_bit27.Q ),
    .X(_015_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _103_ (.Y(_016_),
    .B(_015_),
    .A_N(\Inst_N_IO_ConfigMem.Inst_frame0_bit28.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _104_ (.B1(_016_),
    .VDD(VPWR),
    .Y(net117),
    .VSS(VGND),
    .A1(_005_),
    .A2(_012_));
 sg13g2_mux2_1 _105_ (.A0(net42),
    .A1(net43),
    .S(net70),
    .X(_017_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _106_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_018_),
    .B(net70),
    .A(net40));
 sg13g2_a21oi_1 _107_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_000_),
    .A2(net70),
    .Y(_019_),
    .B1(\Inst_N_IO_ConfigMem.Inst_frame0_bit19.Q ));
 sg13g2_a221oi_1 _108_ (.VSS(VGND),
    .VDD(VPWR),
    .B2(_019_),
    .C1(\Inst_N_IO_ConfigMem.Inst_frame0_bit20.Q ),
    .B1(_018_),
    .A1(\Inst_N_IO_ConfigMem.Inst_frame0_bit19.Q ),
    .Y(_020_),
    .A2(_017_));
 sg13g2_nand2_1 _109_ (.Y(_021_),
    .A(net45),
    .B(net70),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _110_ (.Y(_022_),
    .B(net44),
    .A_N(net70),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _111_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_021_),
    .A2(_022_),
    .Y(_023_),
    .B1(\Inst_N_IO_ConfigMem.Inst_frame0_bit19.Q ));
 sg13g2_nor2b_1 _112_ (.A(net47),
    .B_N(net70),
    .Y(_024_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _113_ (.B1(\Inst_N_IO_ConfigMem.Inst_frame0_bit19.Q ),
    .VDD(VPWR),
    .Y(_025_),
    .VSS(VGND),
    .A1(net46),
    .A2(net70));
 sg13g2_o21ai_1 _114_ (.B1(\Inst_N_IO_ConfigMem.Inst_frame0_bit20.Q ),
    .VDD(VPWR),
    .Y(_026_),
    .VSS(VGND),
    .A1(_024_),
    .A2(_025_));
 sg13g2_o21ai_1 _115_ (.B1(\Inst_N_IO_ConfigMem.Inst_frame0_bit21.Q ),
    .VDD(VPWR),
    .Y(_027_),
    .VSS(VGND),
    .A1(_023_),
    .A2(_026_));
 sg13g2_mux4_1 _116_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame0_bit18.Q ),
    .A0(net48),
    .A1(net49),
    .A2(net50),
    .A3(net51),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame0_bit19.Q ),
    .X(_028_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _117_ (.S0(net70),
    .A0(net52),
    .A1(net53),
    .A2(net54),
    .A3(net55),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame0_bit19.Q ),
    .X(_029_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _118_ (.A0(_028_),
    .A1(_029_),
    .S(\Inst_N_IO_ConfigMem.Inst_frame0_bit20.Q ),
    .X(_030_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _119_ (.Y(_031_),
    .B(_030_),
    .A_N(\Inst_N_IO_ConfigMem.Inst_frame0_bit21.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _120_ (.B1(_031_),
    .VDD(VPWR),
    .Y(net111),
    .VSS(VGND),
    .A1(_020_),
    .A2(_027_));
 sg13g2_mux4_1 _121_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame0_bit17.Q ),
    .A0(net49),
    .A1(net53),
    .A2(net51),
    .A3(net55),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame0_bit16.Q ),
    .X(\Inst_N_IO_switch_matrix.SS4BEG15 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _122_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame0_bit15.Q ),
    .A0(net48),
    .A1(net52),
    .A2(net50),
    .A3(net54),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame0_bit14.Q ),
    .X(\Inst_N_IO_switch_matrix.SS4BEG14 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _123_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame0_bit12.Q ),
    .A0(net92),
    .A1(net94),
    .A2(net58),
    .A3(\Inst_B_IO_1_bidirectional_frame_config_pass.Q ),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame0_bit13.Q ),
    .X(\Inst_N_IO_switch_matrix.SS4BEG13 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _124_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame0_bit10.Q ),
    .A0(net63),
    .A1(net65),
    .A2(net67),
    .A3(\Inst_A_IO_1_bidirectional_frame_config_pass.Q ),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame0_bit11.Q ),
    .X(\Inst_N_IO_switch_matrix.SS4BEG12 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _125_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame0_bit8.Q ),
    .A0(net68),
    .A1(net93),
    .A2(net57),
    .A3(net2),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame0_bit9.Q ),
    .X(\Inst_N_IO_switch_matrix.SS4BEG11 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _126_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame0_bit6.Q ),
    .A0(net56),
    .A1(net64),
    .A2(net66),
    .A3(net1),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame0_bit7.Q ),
    .X(\Inst_N_IO_switch_matrix.SS4BEG10 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _127_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame0_bit4.Q ),
    .A0(net63),
    .A1(net65),
    .A2(net67),
    .A3(net92),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame0_bit5.Q ),
    .X(\Inst_N_IO_switch_matrix.SS4BEG9 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _128_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame0_bit3.Q ),
    .A0(net66),
    .A1(net93),
    .A2(net68),
    .A3(net57),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame0_bit2.Q ),
    .X(\Inst_N_IO_switch_matrix.SS4BEG8 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _129_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame0_bit1.Q ),
    .A0(net49),
    .A1(net53),
    .A2(net51),
    .A3(net55),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame0_bit0.Q ),
    .X(\Inst_N_IO_switch_matrix.SS4BEG7 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _130_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame1_bit31.Q ),
    .A0(net48),
    .A1(net52),
    .A2(net50),
    .A3(net54),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame1_bit30.Q ),
    .X(\Inst_N_IO_switch_matrix.SS4BEG6 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _131_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame1_bit28.Q ),
    .A0(net41),
    .A1(net43),
    .A2(net45),
    .A3(net47),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame1_bit29.Q ),
    .X(\Inst_N_IO_switch_matrix.SS4BEG5 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _132_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame1_bit26.Q ),
    .A0(net40),
    .A1(net42),
    .A2(net44),
    .A3(net46),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame1_bit27.Q ),
    .X(\Inst_N_IO_switch_matrix.SS4BEG4 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _133_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame1_bit24.Q ),
    .A0(net92),
    .A1(net94),
    .A2(net58),
    .A3(\Inst_B_IO_1_bidirectional_frame_config_pass.Q ),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame1_bit25.Q ),
    .X(\Inst_N_IO_switch_matrix.SS4BEG3 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _134_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame1_bit22.Q ),
    .A0(net63),
    .A1(net65),
    .A2(net67),
    .A3(\Inst_A_IO_1_bidirectional_frame_config_pass.Q ),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame1_bit23.Q ),
    .X(\Inst_N_IO_switch_matrix.SS4BEG2 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _135_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame1_bit20.Q ),
    .A0(net68),
    .A1(net93),
    .A2(net57),
    .A3(net2),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame1_bit21.Q ),
    .X(\Inst_N_IO_switch_matrix.SS4BEG1 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _136_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame1_bit18.Q ),
    .A0(net56),
    .A1(net64),
    .A2(net66),
    .A3(net1),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame1_bit19.Q ),
    .X(\Inst_N_IO_switch_matrix.SS4BEG0 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _137_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame1_bit16.Q ),
    .A0(net56),
    .A1(net95),
    .A2(net98),
    .A3(\Inst_B_IO_1_bidirectional_frame_config_pass.Q ),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame1_bit17.Q ),
    .X(\Inst_N_IO_switch_matrix.S4BEG15 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _138_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame1_bit14.Q ),
    .A0(net63),
    .A1(net102),
    .A2(net99),
    .A3(\Inst_A_IO_1_bidirectional_frame_config_pass.Q ),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame1_bit15.Q ),
    .X(\Inst_N_IO_switch_matrix.S4BEG14 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _139_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame1_bit13.Q ),
    .A0(net36),
    .A1(net105),
    .A2(net66),
    .A3(\Inst_B_IO_1_bidirectional_frame_config_pass.Q ),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame1_bit12.Q ),
    .X(\Inst_N_IO_switch_matrix.S4BEG13 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _140_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame1_bit11.Q ),
    .A0(net37),
    .A1(net106),
    .A2(net67),
    .A3(\Inst_A_IO_1_bidirectional_frame_config_pass.Q ),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame1_bit10.Q ),
    .X(\Inst_N_IO_switch_matrix.S4BEG12 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _141_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame1_bit9.Q ),
    .A0(net93),
    .A1(net98),
    .A2(net109),
    .A3(\Inst_B_IO_1_bidirectional_frame_config_pass.Q ),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame1_bit8.Q ),
    .X(\Inst_N_IO_switch_matrix.S4BEG11 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _142_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame1_bit7.Q ),
    .A0(net94),
    .A1(net99),
    .A2(net110),
    .A3(\Inst_A_IO_1_bidirectional_frame_config_pass.Q ),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame1_bit6.Q ),
    .X(\Inst_N_IO_switch_matrix.S4BEG10 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _143_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame1_bit4.Q ),
    .A0(net36),
    .A1(net59),
    .A2(net98),
    .A3(\Inst_B_IO_1_bidirectional_frame_config_pass.Q ),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame1_bit5.Q ),
    .X(\Inst_N_IO_switch_matrix.S4BEG9 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _144_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame1_bit2.Q ),
    .A0(net37),
    .A1(net60),
    .A2(net99),
    .A3(\Inst_A_IO_1_bidirectional_frame_config_pass.Q ),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame1_bit3.Q ),
    .X(\Inst_N_IO_switch_matrix.S4BEG8 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _145_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame1_bit0.Q ),
    .A0(net64),
    .A1(net103),
    .A2(net100),
    .A3(net2),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame1_bit1.Q ),
    .X(\Inst_N_IO_switch_matrix.S4BEG7 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _146_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame2_bit30.Q ),
    .A0(net65),
    .A1(net104),
    .A2(net101),
    .A3(net1),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame2_bit31.Q ),
    .X(\Inst_N_IO_switch_matrix.S4BEG6 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _147_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame2_bit29.Q ),
    .A0(net39),
    .A1(net107),
    .A2(net68),
    .A3(net2),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame2_bit28.Q ),
    .X(\Inst_N_IO_switch_matrix.S4BEG5 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _148_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame2_bit27.Q ),
    .A0(net38),
    .A1(net108),
    .A2(net92),
    .A3(net1),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame2_bit26.Q ),
    .X(\Inst_N_IO_switch_matrix.S4BEG4 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _149_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame2_bit25.Q ),
    .A0(net57),
    .A1(net100),
    .A2(net96),
    .A3(net2),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame2_bit24.Q ),
    .X(\Inst_N_IO_switch_matrix.S4BEG3 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _150_ (.D(net31),
    .GATE(net74),
    .Q(net113),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _151_ (.D(net32),
    .GATE(net71),
    .Q(net114),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _152_ (.D(net33),
    .GATE(net71),
    .Q(net115),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _153_ (.D(net34),
    .GATE(net71),
    .Q(net116),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _154_ (.D(net4),
    .GATE(net74),
    .Q(net119),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _155_ (.D(net5),
    .GATE(net74),
    .Q(net120),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _156_ (.D(net6),
    .GATE(net72),
    .Q(net121),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _157_ (.D(net7),
    .GATE(net73),
    .Q(net122),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _158_ (.D(net8),
    .GATE(net71),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame3_bit14.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _159_ (.D(net9),
    .GATE(net75),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame3_bit15.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _160_ (.D(net10),
    .GATE(net71),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame3_bit16.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _161_ (.D(net11),
    .GATE(net75),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame3_bit17.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _162_ (.D(net12),
    .GATE(net71),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame3_bit18.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _163_ (.D(net13),
    .GATE(net73),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame3_bit19.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _164_ (.D(net15),
    .GATE(net71),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame3_bit20.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _165_ (.D(net16),
    .GATE(net71),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame3_bit21.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _166_ (.D(net17),
    .GATE(net73),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame3_bit22.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _167_ (.D(net18),
    .GATE(net75),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame3_bit23.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _168_ (.D(net19),
    .GATE(net72),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame3_bit24.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _169_ (.D(net20),
    .GATE(net73),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame3_bit25.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _170_ (.D(net21),
    .GATE(net72),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame3_bit26.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _171_ (.D(net22),
    .GATE(net72),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame3_bit27.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _172_ (.D(net23),
    .GATE(net72),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame3_bit28.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _173_ (.D(net24),
    .GATE(net72),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame3_bit29.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _174_ (.D(net26),
    .GATE(net72),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame3_bit30.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _175_ (.D(net27),
    .GATE(net72),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame3_bit31.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _176_ (.D(net3),
    .GATE(net76),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame2_bit0.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _177_ (.D(net14),
    .GATE(net77),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame2_bit1.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _178_ (.D(net25),
    .GATE(net76),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame2_bit2.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _179_ (.D(net28),
    .GATE(net76),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame2_bit3.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _180_ (.D(net29),
    .GATE(net76),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame2_bit4.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _181_ (.D(net30),
    .GATE(net76),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame2_bit5.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _182_ (.D(net31),
    .GATE(net79),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame2_bit6.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _183_ (.D(net32),
    .GATE(net79),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame2_bit7.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _184_ (.D(net33),
    .GATE(net79),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame2_bit8.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _185_ (.D(net34),
    .GATE(net80),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame2_bit9.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _186_ (.D(net4),
    .GATE(net78),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame2_bit10.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _187_ (.D(net5),
    .GATE(net78),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame2_bit11.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _188_ (.D(net6),
    .GATE(net76),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame2_bit12.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _189_ (.D(net7),
    .GATE(net77),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame2_bit13.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _190_ (.D(net8),
    .GATE(net76),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame2_bit14.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _191_ (.D(net9),
    .GATE(net76),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame2_bit15.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _192_ (.D(net10),
    .GATE(net81),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame2_bit16.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _193_ (.D(net11),
    .GATE(net81),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame2_bit17.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _194_ (.D(net12),
    .GATE(net81),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame2_bit18.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _195_ (.D(net13),
    .GATE(net81),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame2_bit19.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _196_ (.D(net15),
    .GATE(net77),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame2_bit20.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _197_ (.D(net16),
    .GATE(net77),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame2_bit21.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _198_ (.D(net17),
    .GATE(net80),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame2_bit22.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _199_ (.D(net18),
    .GATE(net79),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame2_bit23.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _200_ (.D(net19),
    .GATE(net79),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame2_bit24.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _201_ (.D(net20),
    .GATE(net78),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame2_bit25.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _202_ (.D(net21),
    .GATE(net80),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame2_bit26.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _203_ (.D(net22),
    .GATE(net80),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame2_bit27.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _204_ (.D(net23),
    .GATE(net79),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame2_bit28.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _205_ (.D(net24),
    .GATE(net78),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame2_bit29.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _206_ (.D(net26),
    .GATE(net80),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame2_bit30.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _207_ (.D(net27),
    .GATE(net79),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame2_bit31.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _208_ (.D(net3),
    .GATE(net82),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame1_bit0.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _209_ (.D(net14),
    .GATE(net35),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame1_bit1.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _210_ (.D(net25),
    .GATE(net83),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame1_bit2.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _211_ (.D(net28),
    .GATE(net83),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame1_bit3.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _212_ (.D(net29),
    .GATE(net83),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame1_bit4.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _213_ (.D(net30),
    .GATE(net85),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame1_bit5.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _214_ (.D(net31),
    .GATE(net83),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame1_bit6.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _215_ (.D(net32),
    .GATE(net84),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame1_bit7.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _216_ (.D(net33),
    .GATE(net85),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame1_bit8.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _217_ (.D(net34),
    .GATE(net85),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame1_bit9.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _218_ (.D(net4),
    .GATE(net84),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame1_bit10.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _219_ (.D(net5),
    .GATE(net84),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame1_bit11.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _220_ (.D(net6),
    .GATE(net84),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame1_bit12.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _221_ (.D(net7),
    .GATE(net84),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame1_bit13.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _222_ (.D(net8),
    .GATE(net83),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame1_bit14.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _223_ (.D(net9),
    .GATE(net83),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame1_bit15.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _224_ (.D(net10),
    .GATE(net83),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame1_bit16.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _225_ (.D(net11),
    .GATE(net85),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame1_bit17.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _226_ (.D(net12),
    .GATE(net83),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame1_bit18.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _227_ (.D(net13),
    .GATE(net85),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame1_bit19.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _228_ (.D(net15),
    .GATE(net85),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame1_bit20.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _229_ (.D(net16),
    .GATE(net85),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame1_bit21.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _230_ (.D(net17),
    .GATE(net86),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame1_bit22.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _231_ (.D(net18),
    .GATE(net86),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame1_bit23.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _232_ (.D(net19),
    .GATE(net86),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame1_bit24.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _233_ (.D(net20),
    .GATE(net85),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame1_bit25.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _234_ (.D(net21),
    .GATE(net82),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame1_bit26.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _235_ (.D(net22),
    .GATE(net82),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame1_bit27.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _236_ (.D(net23),
    .GATE(net82),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame1_bit28.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _237_ (.D(net24),
    .GATE(net82),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame1_bit29.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _238_ (.D(net26),
    .GATE(net82),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame1_bit30.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _239_ (.D(net27),
    .GATE(net82),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame1_bit31.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _240_ (.D(net3),
    .GATE(net88),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame0_bit0.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _241_ (.D(net14),
    .GATE(net88),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame0_bit1.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _242_ (.D(net25),
    .GATE(net90),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame0_bit2.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _243_ (.D(net28),
    .GATE(net90),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame0_bit3.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _244_ (.D(net29),
    .GATE(net90),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame0_bit4.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _245_ (.D(net30),
    .GATE(net90),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame0_bit5.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _246_ (.D(net31),
    .GATE(net91),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame0_bit6.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _247_ (.D(net32),
    .GATE(net91),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame0_bit7.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _248_ (.D(net33),
    .GATE(net90),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame0_bit8.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _249_ (.D(net34),
    .GATE(net90),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame0_bit9.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _250_ (.D(net4),
    .GATE(net90),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame0_bit10.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _251_ (.D(net5),
    .GATE(net90),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame0_bit11.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _252_ (.D(net6),
    .GATE(net91),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame0_bit12.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _253_ (.D(net7),
    .GATE(net91),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame0_bit13.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _254_ (.D(net8),
    .GATE(net89),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame0_bit14.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _255_ (.D(net9),
    .GATE(net88),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame0_bit15.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _256_ (.D(net10),
    .GATE(net89),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame0_bit16.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _257_ (.D(net11),
    .GATE(net88),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame0_bit17.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _258_ (.D(net12),
    .GATE(net88),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame0_bit18.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _259_ (.D(net13),
    .GATE(net88),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame0_bit19.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _260_ (.D(net15),
    .GATE(net88),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame0_bit20.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _261_ (.D(net16),
    .GATE(net88),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame0_bit21.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _262_ (.D(net17),
    .GATE(net87),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame0_bit22.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _263_ (.D(net18),
    .GATE(net87),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame0_bit23.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _264_ (.D(net19),
    .GATE(net87),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame0_bit24.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _265_ (.D(net20),
    .GATE(net87),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame0_bit25.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _266_ (.D(net21),
    .GATE(net87),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame0_bit26.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _267_ (.D(net22),
    .GATE(net87),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame0_bit27.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _268_ (.D(net23),
    .GATE(net89),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame0_bit28.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _269_ (.D(net24),
    .GATE(net89),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame0_bit29.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _270_ (.D(net26),
    .GATE(net87),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame0_bit30.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _271_ (.D(net27),
    .GATE(net87),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame0_bit31.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dfrbp_1 _272_ (.CLK(UserCLK),
    .RESET_B(net228),
    .D(net1),
    .Q_N(_046_),
    .Q(\Inst_A_IO_1_bidirectional_frame_config_pass.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dfrbp_1 _273_ (.CLK(UserCLK),
    .RESET_B(net229),
    .D(net2),
    .Q_N(_045_),
    .Q(\Inst_B_IO_1_bidirectional_frame_config_pass.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_tiehi _273__206 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net229));
 sg13g2_fill_2 FILLER_0_12 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _276_ (.A(net3),
    .X(net123),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _277_ (.A(net14),
    .X(net134),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _278_ (.A(net25),
    .X(net145),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _279_ (.A(net28),
    .X(net148),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _280_ (.A(net29),
    .X(net149),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _281_ (.A(net30),
    .X(net150),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _282_ (.A(net31),
    .X(net151),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _283_ (.A(net32),
    .X(net152),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _284_ (.A(net33),
    .X(net153),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _285_ (.A(net34),
    .X(net154),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _286_ (.A(net4),
    .X(net124),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _287_ (.A(net5),
    .X(net125),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _288_ (.A(net6),
    .X(net126),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _289_ (.A(net7),
    .X(net127),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _290_ (.A(net8),
    .X(net128),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _291_ (.A(net9),
    .X(net129),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _292_ (.A(net10),
    .X(net130),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _293_ (.A(net11),
    .X(net131),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _294_ (.A(net12),
    .X(net132),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _295_ (.A(net13),
    .X(net133),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _296_ (.A(net15),
    .X(net135),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _297_ (.A(net16),
    .X(net136),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _298_ (.A(net17),
    .X(net137),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _299_ (.A(net18),
    .X(net138),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _300_ (.A(net19),
    .X(net139),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _301_ (.A(net20),
    .X(net140),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _302_ (.A(net21),
    .X(net141),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _303_ (.A(net22),
    .X(net142),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _304_ (.A(net23),
    .X(net143),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _305_ (.A(net24),
    .X(net144),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _306_ (.A(net26),
    .X(net146),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _307_ (.A(net27),
    .X(net147),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _308_ (.A(FrameStrobe[0]),
    .X(net155),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _309_ (.A(net82),
    .X(net166),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _310_ (.A(net79),
    .X(net167),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _311_ (.A(net75),
    .X(net168),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _312_ (.A(FrameStrobe[4]),
    .X(net169),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _313_ (.A(FrameStrobe[5]),
    .X(net170),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _314_ (.A(FrameStrobe[6]),
    .X(net171),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _315_ (.A(FrameStrobe[7]),
    .X(net172),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _316_ (.A(FrameStrobe[8]),
    .X(net173),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _317_ (.A(FrameStrobe[9]),
    .X(net174),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _318_ (.A(FrameStrobe[10]),
    .X(net156),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _319_ (.A(FrameStrobe[11]),
    .X(net157),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _320_ (.A(FrameStrobe[12]),
    .X(net158),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _321_ (.A(FrameStrobe[13]),
    .X(net159),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _322_ (.A(FrameStrobe[14]),
    .X(net160),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _323_ (.A(FrameStrobe[15]),
    .X(net161),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _324_ (.A(FrameStrobe[16]),
    .X(net162),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _325_ (.A(FrameStrobe[17]),
    .X(net163),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _326_ (.A(FrameStrobe[18]),
    .X(net164),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _327_ (.A(FrameStrobe[19]),
    .X(net165),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _328_ (.A(\Inst_N_IO_switch_matrix.S1BEG0 ),
    .X(net175),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _329_ (.A(\Inst_N_IO_switch_matrix.S1BEG1 ),
    .X(net176),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _330_ (.A(\Inst_N_IO_switch_matrix.S1BEG2 ),
    .X(net177),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _331_ (.A(\Inst_N_IO_switch_matrix.S1BEG3 ),
    .X(net178),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _332_ (.A(\Inst_N_IO_switch_matrix.S2BEG0 ),
    .X(net179),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _333_ (.A(\Inst_N_IO_switch_matrix.S2BEG1 ),
    .X(net180),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _334_ (.A(\Inst_N_IO_switch_matrix.S2BEG2 ),
    .X(net181),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _335_ (.A(\Inst_N_IO_switch_matrix.S2BEG3 ),
    .X(net182),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _336_ (.A(\Inst_N_IO_switch_matrix.S2BEG4 ),
    .X(net183),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _337_ (.A(\Inst_N_IO_switch_matrix.S2BEG5 ),
    .X(net184),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _338_ (.A(\Inst_N_IO_switch_matrix.S2BEG6 ),
    .X(net185),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _339_ (.A(\Inst_N_IO_switch_matrix.S2BEG7 ),
    .X(net186),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _340_ (.A(\Inst_N_IO_switch_matrix.S2BEGb0 ),
    .X(net187),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _341_ (.A(\Inst_N_IO_switch_matrix.S2BEGb1 ),
    .X(net188),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _342_ (.A(\Inst_N_IO_switch_matrix.S2BEGb2 ),
    .X(net189),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _343_ (.A(\Inst_N_IO_switch_matrix.S2BEGb3 ),
    .X(net190),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _344_ (.A(\Inst_N_IO_switch_matrix.S2BEGb4 ),
    .X(net191),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _345_ (.A(\Inst_N_IO_switch_matrix.S2BEGb5 ),
    .X(net192),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _346_ (.A(\Inst_N_IO_switch_matrix.S2BEGb6 ),
    .X(net193),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _347_ (.A(\Inst_N_IO_switch_matrix.S2BEGb7 ),
    .X(net194),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _348_ (.A(\Inst_N_IO_switch_matrix.S4BEG0 ),
    .X(net195),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _349_ (.A(\Inst_N_IO_switch_matrix.S4BEG1 ),
    .X(net202),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _350_ (.A(\Inst_N_IO_switch_matrix.S4BEG2 ),
    .X(net203),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _351_ (.A(\Inst_N_IO_switch_matrix.S4BEG3 ),
    .X(net204),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _352_ (.A(\Inst_N_IO_switch_matrix.S4BEG4 ),
    .X(net205),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _353_ (.A(\Inst_N_IO_switch_matrix.S4BEG5 ),
    .X(net206),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _354_ (.A(\Inst_N_IO_switch_matrix.S4BEG6 ),
    .X(net207),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _355_ (.A(\Inst_N_IO_switch_matrix.S4BEG7 ),
    .X(net208),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _356_ (.A(\Inst_N_IO_switch_matrix.S4BEG8 ),
    .X(net209),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _357_ (.A(\Inst_N_IO_switch_matrix.S4BEG9 ),
    .X(net210),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _358_ (.A(\Inst_N_IO_switch_matrix.S4BEG10 ),
    .X(net196),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _359_ (.A(\Inst_N_IO_switch_matrix.S4BEG11 ),
    .X(net197),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _360_ (.A(\Inst_N_IO_switch_matrix.S4BEG12 ),
    .X(net198),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _361_ (.A(\Inst_N_IO_switch_matrix.S4BEG13 ),
    .X(net199),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _362_ (.A(\Inst_N_IO_switch_matrix.S4BEG14 ),
    .X(net200),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _363_ (.A(\Inst_N_IO_switch_matrix.S4BEG15 ),
    .X(net201),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _364_ (.A(\Inst_N_IO_switch_matrix.SS4BEG0 ),
    .X(net211),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _365_ (.A(\Inst_N_IO_switch_matrix.SS4BEG1 ),
    .X(net218),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _366_ (.A(\Inst_N_IO_switch_matrix.SS4BEG2 ),
    .X(net219),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _367_ (.A(\Inst_N_IO_switch_matrix.SS4BEG3 ),
    .X(net220),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _368_ (.A(\Inst_N_IO_switch_matrix.SS4BEG4 ),
    .X(net221),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _369_ (.A(\Inst_N_IO_switch_matrix.SS4BEG5 ),
    .X(net222),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _370_ (.A(\Inst_N_IO_switch_matrix.SS4BEG6 ),
    .X(net223),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _371_ (.A(\Inst_N_IO_switch_matrix.SS4BEG7 ),
    .X(net224),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _372_ (.A(\Inst_N_IO_switch_matrix.SS4BEG8 ),
    .X(net225),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _373_ (.A(\Inst_N_IO_switch_matrix.SS4BEG9 ),
    .X(net226),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _374_ (.A(\Inst_N_IO_switch_matrix.SS4BEG10 ),
    .X(net212),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _375_ (.A(\Inst_N_IO_switch_matrix.SS4BEG11 ),
    .X(net213),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _376_ (.A(\Inst_N_IO_switch_matrix.SS4BEG12 ),
    .X(net214),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _377_ (.A(\Inst_N_IO_switch_matrix.SS4BEG13 ),
    .X(net215),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _378_ (.A(\Inst_N_IO_switch_matrix.SS4BEG14 ),
    .X(net216),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _379_ (.A(\Inst_N_IO_switch_matrix.SS4BEG15 ),
    .X(net217),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _380_ (.A(UserCLK),
    .X(net227),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout69 (.A(\Inst_N_IO_ConfigMem.Inst_frame0_bit25.Q ),
    .X(net69),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout70 (.A(\Inst_N_IO_ConfigMem.Inst_frame0_bit18.Q ),
    .X(net70),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout71 (.A(net74),
    .X(net71),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout72 (.A(net73),
    .X(net72),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout73 (.A(net74),
    .X(net73),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout74 (.A(net75),
    .X(net74),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout75 (.A(FrameStrobe[3]),
    .X(net75),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout76 (.A(net78),
    .X(net76),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout77 (.A(net78),
    .X(net77),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout78 (.A(FrameStrobe[2]),
    .X(net78),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout79 (.A(net81),
    .X(net79),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout80 (.A(net81),
    .X(net80),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout81 (.A(FrameStrobe[2]),
    .X(net81),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout82 (.A(net35),
    .X(net82),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout83 (.A(net86),
    .X(net83),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout84 (.A(net86),
    .X(net84),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout85 (.A(net86),
    .X(net85),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout86 (.A(net35),
    .X(net86),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout87 (.A(net89),
    .X(net87),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout88 (.A(net89),
    .X(net88),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout89 (.A(FrameStrobe[0]),
    .X(net89),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout90 (.A(net91),
    .X(net90),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout91 (.A(FrameStrobe[0]),
    .X(net91),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input1 (.A(A_O_top),
    .X(net1),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input2 (.A(B_O_top),
    .X(net2),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input3 (.A(FrameData[0]),
    .X(net3),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input4 (.A(FrameData[10]),
    .X(net4),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input5 (.A(FrameData[11]),
    .X(net5),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input6 (.A(FrameData[12]),
    .X(net6),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input7 (.A(FrameData[13]),
    .X(net7),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input8 (.A(FrameData[14]),
    .X(net8),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input9 (.A(FrameData[15]),
    .X(net9),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input10 (.A(FrameData[16]),
    .X(net10),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input11 (.A(FrameData[17]),
    .X(net11),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input12 (.A(FrameData[18]),
    .X(net12),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input13 (.A(FrameData[19]),
    .X(net13),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input14 (.A(FrameData[1]),
    .X(net14),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input15 (.A(FrameData[20]),
    .X(net15),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input16 (.A(FrameData[21]),
    .X(net16),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input17 (.A(FrameData[22]),
    .X(net17),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input18 (.A(FrameData[23]),
    .X(net18),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input19 (.A(FrameData[24]),
    .X(net19),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input20 (.A(FrameData[25]),
    .X(net20),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input21 (.A(FrameData[26]),
    .X(net21),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input22 (.A(FrameData[27]),
    .X(net22),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input23 (.A(FrameData[28]),
    .X(net23),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input24 (.A(FrameData[29]),
    .X(net24),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input25 (.A(FrameData[2]),
    .X(net25),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input26 (.A(FrameData[30]),
    .X(net26),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input27 (.A(FrameData[31]),
    .X(net27),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input28 (.A(FrameData[3]),
    .X(net28),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input29 (.A(FrameData[4]),
    .X(net29),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input30 (.A(FrameData[5]),
    .X(net30),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input31 (.A(FrameData[6]),
    .X(net31),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input32 (.A(FrameData[7]),
    .X(net32),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input33 (.A(FrameData[8]),
    .X(net33),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input34 (.A(FrameData[9]),
    .X(net34),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input35 (.A(FrameStrobe[1]),
    .X(net35),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input36 (.A(N1END[0]),
    .X(net36),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input37 (.A(N1END[1]),
    .X(net37),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input38 (.A(N1END[2]),
    .X(net38),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input39 (.A(N1END[3]),
    .X(net39),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input40 (.A(N2END[0]),
    .X(net40),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input41 (.A(N2END[1]),
    .X(net41),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input42 (.A(N2END[2]),
    .X(net42),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input43 (.A(N2END[3]),
    .X(net43),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input44 (.A(N2END[4]),
    .X(net44),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input45 (.A(N2END[5]),
    .X(net45),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input46 (.A(N2END[6]),
    .X(net46),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input47 (.A(N2END[7]),
    .X(net47),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input48 (.A(N2MID[0]),
    .X(net48),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input49 (.A(N2MID[1]),
    .X(net49),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input50 (.A(N2MID[2]),
    .X(net50),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input51 (.A(N2MID[3]),
    .X(net51),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input52 (.A(N2MID[4]),
    .X(net52),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input53 (.A(N2MID[5]),
    .X(net53),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input54 (.A(N2MID[6]),
    .X(net54),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input55 (.A(N2MID[7]),
    .X(net55),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input56 (.A(N4END[0]),
    .X(net56),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input57 (.A(N4END[10]),
    .X(net57),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input58 (.A(N4END[11]),
    .X(net58),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input59 (.A(N4END[12]),
    .X(net59),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input60 (.A(N4END[13]),
    .X(net60),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input61 (.A(N4END[14]),
    .X(net61),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input62 (.A(N4END[15]),
    .X(net62),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input63 (.A(N4END[1]),
    .X(net63),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input64 (.A(N4END[2]),
    .X(net64),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input65 (.A(N4END[3]),
    .X(net65),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input66 (.A(N4END[4]),
    .X(net66),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input67 (.A(N4END[5]),
    .X(net67),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input68 (.A(N4END[6]),
    .X(net68),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input69 (.A(N4END[7]),
    .X(net92),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input70 (.A(N4END[8]),
    .X(net93),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input71 (.A(N4END[9]),
    .X(net94),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input72 (.A(NN4END[0]),
    .X(net95),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input73 (.A(NN4END[10]),
    .X(net96),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input74 (.A(NN4END[11]),
    .X(net97),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input75 (.A(NN4END[12]),
    .X(net98),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input76 (.A(NN4END[13]),
    .X(net99),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input77 (.A(NN4END[14]),
    .X(net100),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input78 (.A(NN4END[15]),
    .X(net101),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input79 (.A(NN4END[1]),
    .X(net102),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input80 (.A(NN4END[2]),
    .X(net103),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input81 (.A(NN4END[3]),
    .X(net104),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input82 (.A(NN4END[4]),
    .X(net105),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input83 (.A(NN4END[5]),
    .X(net106),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input84 (.A(NN4END[6]),
    .X(net107),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input85 (.A(NN4END[7]),
    .X(net108),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input86 (.A(NN4END[8]),
    .X(net109),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input87 (.A(NN4END[9]),
    .X(net110),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output88 (.A(net111),
    .X(A_I_top),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output89 (.A(net112),
    .X(A_T_top),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output90 (.A(net113),
    .X(A_config_C_bit0),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output91 (.A(net114),
    .X(A_config_C_bit1),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output92 (.A(net115),
    .X(A_config_C_bit2),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output93 (.A(net116),
    .X(A_config_C_bit3),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output94 (.A(net117),
    .X(B_I_top),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output95 (.A(net118),
    .X(B_T_top),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output96 (.A(net119),
    .X(B_config_C_bit0),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output97 (.A(net120),
    .X(B_config_C_bit1),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output98 (.A(net121),
    .X(B_config_C_bit2),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output99 (.A(net122),
    .X(B_config_C_bit3),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output100 (.A(net123),
    .X(FrameData_O[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output101 (.A(net124),
    .X(FrameData_O[10]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output102 (.A(net125),
    .X(FrameData_O[11]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output103 (.A(net126),
    .X(FrameData_O[12]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output104 (.A(net127),
    .X(FrameData_O[13]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output105 (.A(net128),
    .X(FrameData_O[14]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output106 (.A(net129),
    .X(FrameData_O[15]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output107 (.A(net130),
    .X(FrameData_O[16]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output108 (.A(net131),
    .X(FrameData_O[17]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output109 (.A(net132),
    .X(FrameData_O[18]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output110 (.A(net133),
    .X(FrameData_O[19]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output111 (.A(net134),
    .X(FrameData_O[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output112 (.A(net135),
    .X(FrameData_O[20]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output113 (.A(net136),
    .X(FrameData_O[21]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output114 (.A(net137),
    .X(FrameData_O[22]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output115 (.A(net138),
    .X(FrameData_O[23]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output116 (.A(net139),
    .X(FrameData_O[24]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output117 (.A(net140),
    .X(FrameData_O[25]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output118 (.A(net141),
    .X(FrameData_O[26]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output119 (.A(net142),
    .X(FrameData_O[27]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output120 (.A(net143),
    .X(FrameData_O[28]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output121 (.A(net144),
    .X(FrameData_O[29]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output122 (.A(net145),
    .X(FrameData_O[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output123 (.A(net146),
    .X(FrameData_O[30]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output124 (.A(net147),
    .X(FrameData_O[31]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output125 (.A(net148),
    .X(FrameData_O[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output126 (.A(net149),
    .X(FrameData_O[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output127 (.A(net150),
    .X(FrameData_O[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output128 (.A(net151),
    .X(FrameData_O[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output129 (.A(net152),
    .X(FrameData_O[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output130 (.A(net153),
    .X(FrameData_O[8]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output131 (.A(net154),
    .X(FrameData_O[9]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output132 (.A(net155),
    .X(FrameStrobe_O[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output133 (.A(net156),
    .X(FrameStrobe_O[10]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output134 (.A(net157),
    .X(FrameStrobe_O[11]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output135 (.A(net158),
    .X(FrameStrobe_O[12]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output136 (.A(net159),
    .X(FrameStrobe_O[13]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output137 (.A(net160),
    .X(FrameStrobe_O[14]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output138 (.A(net161),
    .X(FrameStrobe_O[15]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output139 (.A(net162),
    .X(FrameStrobe_O[16]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output140 (.A(net163),
    .X(FrameStrobe_O[17]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output141 (.A(net164),
    .X(FrameStrobe_O[18]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output142 (.A(net165),
    .X(FrameStrobe_O[19]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output143 (.A(net166),
    .X(FrameStrobe_O[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output144 (.A(net167),
    .X(FrameStrobe_O[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output145 (.A(net168),
    .X(FrameStrobe_O[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output146 (.A(net169),
    .X(FrameStrobe_O[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output147 (.A(net170),
    .X(FrameStrobe_O[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output148 (.A(net171),
    .X(FrameStrobe_O[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output149 (.A(net172),
    .X(FrameStrobe_O[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output150 (.A(net173),
    .X(FrameStrobe_O[8]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output151 (.A(net174),
    .X(FrameStrobe_O[9]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output152 (.A(net175),
    .X(S1BEG[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output153 (.A(net176),
    .X(S1BEG[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output154 (.A(net177),
    .X(S1BEG[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output155 (.A(net178),
    .X(S1BEG[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output156 (.A(net179),
    .X(S2BEG[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output157 (.A(net180),
    .X(S2BEG[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output158 (.A(net181),
    .X(S2BEG[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output159 (.A(net182),
    .X(S2BEG[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output160 (.A(net183),
    .X(S2BEG[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output161 (.A(net184),
    .X(S2BEG[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output162 (.A(net185),
    .X(S2BEG[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output163 (.A(net186),
    .X(S2BEG[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output164 (.A(net187),
    .X(S2BEGb[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output165 (.A(net188),
    .X(S2BEGb[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output166 (.A(net189),
    .X(S2BEGb[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output167 (.A(net190),
    .X(S2BEGb[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output168 (.A(net191),
    .X(S2BEGb[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output169 (.A(net192),
    .X(S2BEGb[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output170 (.A(net193),
    .X(S2BEGb[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output171 (.A(net194),
    .X(S2BEGb[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output172 (.A(net195),
    .X(S4BEG[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output173 (.A(net196),
    .X(S4BEG[10]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output174 (.A(net197),
    .X(S4BEG[11]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output175 (.A(net198),
    .X(S4BEG[12]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output176 (.A(net199),
    .X(S4BEG[13]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output177 (.A(net200),
    .X(S4BEG[14]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output178 (.A(net201),
    .X(S4BEG[15]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output179 (.A(net202),
    .X(S4BEG[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output180 (.A(net203),
    .X(S4BEG[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output181 (.A(net204),
    .X(S4BEG[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output182 (.A(net205),
    .X(S4BEG[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output183 (.A(net206),
    .X(S4BEG[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output184 (.A(net207),
    .X(S4BEG[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output185 (.A(net208),
    .X(S4BEG[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output186 (.A(net209),
    .X(S4BEG[8]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output187 (.A(net210),
    .X(S4BEG[9]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output188 (.A(net211),
    .X(SS4BEG[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output189 (.A(net212),
    .X(SS4BEG[10]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output190 (.A(net213),
    .X(SS4BEG[11]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output191 (.A(net214),
    .X(SS4BEG[12]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output192 (.A(net215),
    .X(SS4BEG[13]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output193 (.A(net216),
    .X(SS4BEG[14]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output194 (.A(net217),
    .X(SS4BEG[15]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output195 (.A(net218),
    .X(SS4BEG[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output196 (.A(net219),
    .X(SS4BEG[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output197 (.A(net220),
    .X(SS4BEG[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output198 (.A(net221),
    .X(SS4BEG[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output199 (.A(net222),
    .X(SS4BEG[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output200 (.A(net223),
    .X(SS4BEG[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output201 (.A(net224),
    .X(SS4BEG[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output202 (.A(net225),
    .X(SS4BEG[8]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output203 (.A(net226),
    .X(SS4BEG[9]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output204 (.A(net227),
    .X(UserCLKo),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_tiehi _272__205 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net228));
 sg13g2_fill_1 FILLER_0_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_16 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_38 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_341 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_10 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_107 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_12 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_22 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_10 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_397 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_12 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_80 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_44 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_15 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_37 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_121 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_227 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_426 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_12 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_27 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_90 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_12 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_19 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_26 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_30 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_71 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_80 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_20 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_24 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_29 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_36 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_38 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_383 (.VDD(VPWR),
    .VSS(VGND));
endmodule
