magic
tech sky130A
magscale 1 2
timestamp 1740383483
<< viali >>
rect 1409 8585 1443 8619
rect 2973 8585 3007 8619
rect 4537 8585 4571 8619
rect 6469 8585 6503 8619
rect 7665 8585 7699 8619
rect 9229 8585 9263 8619
rect 10793 8585 10827 8619
rect 12357 8585 12391 8619
rect 14197 8585 14231 8619
rect 15485 8585 15519 8619
rect 17049 8585 17083 8619
rect 18613 8585 18647 8619
rect 20177 8585 20211 8619
rect 21925 8585 21959 8619
rect 23397 8585 23431 8619
rect 24961 8585 24995 8619
rect 26525 8585 26559 8619
rect 28089 8585 28123 8619
rect 29745 8585 29779 8619
rect 30113 8585 30147 8619
rect 30481 8585 30515 8619
rect 31217 8585 31251 8619
rect 1593 8449 1627 8483
rect 3157 8449 3191 8483
rect 4721 8449 4755 8483
rect 6653 8449 6687 8483
rect 7849 8449 7883 8483
rect 9413 8449 9447 8483
rect 10977 8449 11011 8483
rect 12541 8449 12575 8483
rect 14381 8449 14415 8483
rect 15662 8449 15696 8483
rect 17233 8449 17267 8483
rect 18797 8449 18831 8483
rect 20361 8449 20395 8483
rect 22109 8449 22143 8483
rect 23213 8449 23247 8483
rect 24777 8449 24811 8483
rect 26341 8449 26375 8483
rect 27905 8449 27939 8483
rect 29561 8449 29595 8483
rect 29929 8449 29963 8483
rect 30297 8449 30331 8483
rect 30665 8449 30699 8483
rect 31033 8449 31067 8483
rect 31677 8449 31711 8483
rect 30849 8313 30883 8347
rect 31861 8313 31895 8347
rect 30665 8041 30699 8075
rect 31033 8041 31067 8075
rect 31401 8041 31435 8075
rect 30481 7837 30515 7871
rect 30849 7837 30883 7871
rect 31217 7837 31251 7871
rect 31585 7837 31619 7871
rect 31953 7837 31987 7871
rect 31769 7701 31803 7735
rect 32137 7701 32171 7735
rect 4905 7497 4939 7531
rect 6745 7497 6779 7531
rect 7665 7497 7699 7531
rect 13369 7497 13403 7531
rect 15301 7497 15335 7531
rect 16037 7497 16071 7531
rect 16405 7497 16439 7531
rect 17785 7497 17819 7531
rect 18153 7497 18187 7531
rect 19717 7497 19751 7531
rect 20269 7497 20303 7531
rect 22937 7497 22971 7531
rect 24225 7497 24259 7531
rect 25145 7497 25179 7531
rect 25329 7497 25363 7531
rect 31493 7497 31527 7531
rect 13461 7429 13495 7463
rect 17141 7429 17175 7463
rect 4721 7361 4755 7395
rect 5733 7361 5767 7395
rect 6009 7361 6043 7395
rect 6561 7361 6595 7395
rect 6837 7361 6871 7395
rect 7205 7361 7239 7395
rect 7481 7361 7515 7395
rect 8769 7361 8803 7395
rect 9045 7361 9079 7395
rect 9321 7361 9355 7395
rect 11897 7361 11931 7395
rect 12173 7361 12207 7395
rect 12449 7361 12483 7395
rect 12817 7361 12851 7395
rect 12909 7361 12943 7395
rect 13645 7361 13679 7395
rect 13737 7361 13771 7395
rect 14013 7361 14047 7395
rect 14449 7361 14483 7395
rect 14565 7361 14599 7395
rect 14749 7361 14783 7395
rect 15025 7361 15059 7395
rect 15301 7361 15335 7395
rect 16129 7361 16163 7395
rect 16221 7361 16255 7395
rect 16681 7361 16715 7395
rect 16957 7361 16991 7395
rect 17233 7361 17267 7395
rect 17325 7361 17359 7395
rect 17877 7361 17911 7395
rect 17969 7361 18003 7395
rect 19901 7361 19935 7395
rect 20453 7361 20487 7395
rect 20913 7361 20947 7395
rect 23121 7361 23155 7395
rect 24409 7361 24443 7395
rect 24961 7361 24995 7395
rect 25513 7361 25547 7395
rect 31309 7361 31343 7395
rect 31677 7361 31711 7395
rect 13277 7293 13311 7327
rect 5917 7225 5951 7259
rect 8953 7225 8987 7259
rect 13553 7225 13587 7259
rect 13921 7225 13955 7259
rect 15209 7225 15243 7259
rect 6193 7157 6227 7191
rect 7021 7157 7055 7191
rect 7389 7157 7423 7191
rect 9229 7157 9263 7191
rect 9505 7157 9539 7191
rect 12081 7157 12115 7191
rect 12357 7157 12391 7191
rect 12633 7157 12667 7191
rect 12725 7157 12759 7191
rect 13093 7157 13127 7191
rect 14197 7157 14231 7191
rect 14289 7157 14323 7191
rect 14933 7157 14967 7191
rect 16865 7157 16899 7191
rect 17509 7157 17543 7191
rect 20729 7157 20763 7191
rect 31861 7157 31895 7191
rect 5733 6749 5767 6783
rect 8033 6749 8067 6783
rect 8401 6749 8435 6783
rect 8953 6749 8987 6783
rect 17233 6749 17267 6783
rect 19441 6749 19475 6783
rect 19533 6749 19567 6783
rect 25329 6749 25363 6783
rect 31217 6749 31251 6783
rect 31585 6749 31619 6783
rect 31953 6749 31987 6783
rect 5917 6613 5951 6647
rect 8217 6613 8251 6647
rect 8585 6613 8619 6647
rect 9137 6613 9171 6647
rect 17049 6613 17083 6647
rect 17417 6613 17451 6647
rect 19349 6613 19383 6647
rect 19717 6613 19751 6647
rect 25145 6613 25179 6647
rect 31401 6613 31435 6647
rect 31769 6613 31803 6647
rect 32137 6613 32171 6647
rect 31861 6409 31895 6443
rect 7205 6273 7239 6307
rect 9781 6273 9815 6307
rect 20637 6273 20671 6307
rect 21097 6273 21131 6307
rect 21189 6273 21223 6307
rect 31309 6273 31343 6307
rect 31677 6273 31711 6307
rect 20453 6137 20487 6171
rect 7389 6069 7423 6103
rect 9965 6069 9999 6103
rect 21005 6069 21039 6103
rect 21373 6069 21407 6103
rect 31493 6069 31527 6103
rect 29193 5797 29227 5831
rect 31401 5797 31435 5831
rect 32137 5797 32171 5831
rect 3801 5661 3835 5695
rect 10977 5661 11011 5695
rect 18153 5661 18187 5695
rect 18245 5661 18279 5695
rect 21189 5661 21223 5695
rect 22109 5661 22143 5695
rect 29009 5661 29043 5695
rect 30665 5661 30699 5695
rect 31217 5661 31251 5695
rect 31585 5661 31619 5695
rect 31953 5661 31987 5695
rect 3985 5525 4019 5559
rect 11161 5525 11195 5559
rect 18061 5525 18095 5559
rect 18429 5525 18463 5559
rect 21005 5525 21039 5559
rect 21925 5525 21959 5559
rect 30849 5525 30883 5559
rect 31769 5525 31803 5559
rect 23673 5321 23707 5355
rect 27169 5321 27203 5355
rect 5457 5185 5491 5219
rect 10609 5185 10643 5219
rect 23213 5185 23247 5219
rect 23305 5185 23339 5219
rect 23857 5185 23891 5219
rect 26985 5185 27019 5219
rect 31309 5185 31343 5219
rect 31677 5185 31711 5219
rect 5641 4981 5675 5015
rect 10793 4981 10827 5015
rect 23121 4981 23155 5015
rect 23489 4981 23523 5015
rect 31493 4981 31527 5015
rect 31861 4981 31895 5015
rect 12541 4777 12575 4811
rect 25053 4777 25087 4811
rect 11713 4709 11747 4743
rect 13001 4709 13035 4743
rect 2605 4573 2639 4607
rect 11529 4573 11563 4607
rect 12357 4573 12391 4607
rect 12817 4573 12851 4607
rect 14197 4573 14231 4607
rect 24869 4573 24903 4607
rect 25237 4573 25271 4607
rect 25329 4573 25363 4607
rect 31585 4573 31619 4607
rect 31953 4573 31987 4607
rect 2789 4437 2823 4471
rect 14381 4437 14415 4471
rect 25145 4437 25179 4471
rect 25513 4437 25547 4471
rect 31769 4437 31803 4471
rect 32137 4437 32171 4471
rect 13277 4233 13311 4267
rect 18245 4233 18279 4267
rect 12173 4097 12207 4131
rect 12449 4097 12483 4131
rect 12725 4097 12759 4131
rect 13093 4097 13127 4131
rect 13553 4097 13587 4131
rect 13829 4097 13863 4131
rect 14197 4097 14231 4131
rect 14473 4097 14507 4131
rect 15117 4097 15151 4131
rect 15761 4097 15795 4131
rect 16681 4097 16715 4131
rect 17141 4097 17175 4131
rect 17509 4097 17543 4131
rect 17601 4097 17635 4131
rect 18061 4097 18095 4131
rect 19073 4097 19107 4131
rect 19441 4097 19475 4131
rect 19717 4097 19751 4131
rect 22385 4097 22419 4131
rect 23305 4097 23339 4131
rect 23489 4097 23523 4131
rect 23857 4097 23891 4131
rect 31309 4097 31343 4131
rect 31677 4097 31711 4131
rect 18981 4029 19015 4063
rect 19349 3961 19383 3995
rect 22201 3961 22235 3995
rect 23121 3961 23155 3995
rect 23673 3961 23707 3995
rect 24041 3961 24075 3995
rect 12357 3893 12391 3927
rect 12633 3893 12667 3927
rect 12909 3893 12943 3927
rect 13737 3893 13771 3927
rect 14013 3893 14047 3927
rect 14381 3893 14415 3927
rect 14657 3893 14691 3927
rect 15301 3893 15335 3927
rect 15945 3893 15979 3927
rect 16865 3893 16899 3927
rect 17325 3893 17359 3927
rect 17417 3893 17451 3927
rect 17785 3893 17819 3927
rect 19625 3893 19659 3927
rect 19901 3893 19935 3927
rect 31493 3893 31527 3927
rect 31861 3893 31895 3927
rect 21925 3621 21959 3655
rect 25605 3621 25639 3655
rect 12449 3485 12483 3519
rect 19809 3485 19843 3519
rect 20085 3485 20119 3519
rect 20545 3485 20579 3519
rect 20637 3485 20671 3519
rect 21281 3485 21315 3519
rect 21465 3485 21499 3519
rect 21741 3485 21775 3519
rect 22017 3485 22051 3519
rect 25329 3485 25363 3519
rect 25421 3485 25455 3519
rect 25881 3485 25915 3519
rect 25973 3485 26007 3519
rect 26341 3485 26375 3519
rect 26433 3485 26467 3519
rect 31585 3485 31619 3519
rect 31953 3485 31987 3519
rect 25237 3417 25271 3451
rect 12633 3349 12667 3383
rect 19993 3349 20027 3383
rect 20269 3349 20303 3383
rect 20453 3349 20487 3383
rect 20821 3349 20855 3383
rect 21649 3349 21683 3383
rect 25789 3349 25823 3383
rect 26157 3349 26191 3383
rect 26249 3349 26283 3383
rect 26617 3349 26651 3383
rect 31769 3349 31803 3383
rect 32137 3349 32171 3383
rect 14473 3009 14507 3043
rect 15301 3009 15335 3043
rect 16129 3009 16163 3043
rect 19441 3009 19475 3043
rect 20545 3009 20579 3043
rect 20913 3009 20947 3043
rect 21833 3009 21867 3043
rect 22753 3009 22787 3043
rect 23305 3009 23339 3043
rect 23857 3009 23891 3043
rect 31309 3009 31343 3043
rect 31677 3009 31711 3043
rect 14657 2805 14691 2839
rect 15485 2805 15519 2839
rect 16313 2805 16347 2839
rect 19625 2805 19659 2839
rect 20729 2805 20763 2839
rect 21097 2805 21131 2839
rect 22017 2805 22051 2839
rect 22937 2805 22971 2839
rect 23489 2805 23523 2839
rect 24041 2805 24075 2839
rect 31493 2805 31527 2839
rect 31861 2805 31895 2839
rect 18613 2601 18647 2635
rect 20545 2601 20579 2635
rect 22385 2601 22419 2635
rect 23489 2601 23523 2635
rect 18981 2533 19015 2567
rect 20913 2533 20947 2567
rect 22753 2533 22787 2567
rect 23857 2533 23891 2567
rect 13645 2397 13679 2431
rect 14369 2397 14403 2431
rect 14749 2397 14783 2431
rect 15117 2397 15151 2431
rect 15485 2397 15519 2431
rect 15853 2397 15887 2431
rect 16221 2397 16255 2431
rect 16773 2397 16807 2431
rect 17141 2397 17175 2431
rect 17509 2397 17543 2431
rect 18061 2397 18095 2431
rect 18429 2397 18463 2431
rect 18785 2397 18819 2431
rect 19257 2397 19291 2431
rect 19625 2397 19659 2431
rect 19993 2397 20027 2431
rect 20361 2397 20395 2431
rect 20729 2397 20763 2431
rect 21097 2397 21131 2431
rect 21833 2397 21867 2431
rect 22201 2397 22235 2431
rect 22569 2397 22603 2431
rect 22937 2397 22971 2431
rect 23305 2397 23339 2431
rect 23673 2397 23707 2431
rect 24409 2397 24443 2431
rect 30573 2397 30607 2431
rect 30941 2397 30975 2431
rect 31309 2397 31343 2431
rect 31677 2397 31711 2431
rect 13829 2261 13863 2295
rect 14565 2261 14599 2295
rect 14933 2261 14967 2295
rect 15301 2261 15335 2295
rect 15669 2261 15703 2295
rect 16037 2261 16071 2295
rect 16405 2261 16439 2295
rect 16957 2261 16991 2295
rect 17325 2261 17359 2295
rect 17693 2261 17727 2295
rect 18245 2261 18279 2295
rect 19441 2261 19475 2295
rect 19809 2261 19843 2295
rect 20177 2261 20211 2295
rect 21281 2261 21315 2295
rect 22017 2261 22051 2295
rect 23121 2261 23155 2295
rect 24593 2261 24627 2295
rect 30757 2261 30791 2295
rect 31125 2261 31159 2295
rect 31493 2261 31527 2295
rect 31861 2261 31895 2295
<< metal1 >>
rect 16758 9392 16764 9444
rect 16816 9432 16822 9444
rect 24946 9432 24952 9444
rect 16816 9404 24952 9432
rect 16816 9392 16822 9404
rect 24946 9392 24952 9404
rect 25004 9392 25010 9444
rect 17310 9324 17316 9376
rect 17368 9364 17374 9376
rect 25314 9364 25320 9376
rect 17368 9336 25320 9364
rect 17368 9324 17374 9336
rect 25314 9324 25320 9336
rect 25372 9324 25378 9376
rect 14274 9256 14280 9308
rect 14332 9296 14338 9308
rect 30650 9296 30656 9308
rect 14332 9268 30656 9296
rect 14332 9256 14338 9268
rect 30650 9256 30656 9268
rect 30708 9256 30714 9308
rect 9398 9188 9404 9240
rect 9456 9228 9462 9240
rect 19518 9228 19524 9240
rect 9456 9200 19524 9228
rect 9456 9188 9462 9200
rect 19518 9188 19524 9200
rect 19576 9188 19582 9240
rect 12526 9120 12532 9172
rect 12584 9160 12590 9172
rect 17310 9160 17316 9172
rect 12584 9132 17316 9160
rect 12584 9120 12590 9132
rect 17310 9120 17316 9132
rect 17368 9120 17374 9172
rect 17402 9120 17408 9172
rect 17460 9160 17466 9172
rect 24210 9160 24216 9172
rect 17460 9132 24216 9160
rect 17460 9120 17466 9132
rect 24210 9120 24216 9132
rect 24268 9120 24274 9172
rect 12618 9052 12624 9104
rect 12676 9092 12682 9104
rect 30282 9092 30288 9104
rect 12676 9064 30288 9092
rect 12676 9052 12682 9064
rect 30282 9052 30288 9064
rect 30340 9052 30346 9104
rect 17862 9024 17868 9036
rect 4724 8996 17868 9024
rect 4724 8832 4752 8996
rect 17862 8984 17868 8996
rect 17920 8984 17926 9036
rect 4982 8916 4988 8968
rect 5040 8956 5046 8968
rect 17402 8956 17408 8968
rect 5040 8928 17408 8956
rect 5040 8916 5046 8928
rect 17402 8916 17408 8928
rect 17460 8916 17466 8968
rect 17494 8916 17500 8968
rect 17552 8956 17558 8968
rect 29914 8956 29920 8968
rect 17552 8928 29920 8956
rect 17552 8916 17558 8928
rect 29914 8916 29920 8928
rect 29972 8916 29978 8968
rect 10962 8848 10968 8900
rect 11020 8888 11026 8900
rect 11020 8860 16896 8888
rect 11020 8848 11026 8860
rect 4706 8780 4712 8832
rect 4764 8780 4770 8832
rect 14366 8780 14372 8832
rect 14424 8820 14430 8832
rect 16758 8820 16764 8832
rect 14424 8792 16764 8820
rect 14424 8780 14430 8792
rect 16758 8780 16764 8792
rect 16816 8780 16822 8832
rect 16868 8820 16896 8860
rect 17034 8848 17040 8900
rect 17092 8888 17098 8900
rect 23382 8888 23388 8900
rect 17092 8860 23388 8888
rect 17092 8848 17098 8860
rect 23382 8848 23388 8860
rect 23440 8848 23446 8900
rect 22922 8820 22928 8832
rect 16868 8792 22928 8820
rect 22922 8780 22928 8792
rect 22980 8780 22986 8832
rect 1104 8730 32568 8752
rect 1104 8678 3010 8730
rect 3062 8678 3074 8730
rect 3126 8678 3138 8730
rect 3190 8678 3202 8730
rect 3254 8678 3266 8730
rect 3318 8678 9010 8730
rect 9062 8678 9074 8730
rect 9126 8678 9138 8730
rect 9190 8678 9202 8730
rect 9254 8678 9266 8730
rect 9318 8678 15010 8730
rect 15062 8678 15074 8730
rect 15126 8678 15138 8730
rect 15190 8678 15202 8730
rect 15254 8678 15266 8730
rect 15318 8678 21010 8730
rect 21062 8678 21074 8730
rect 21126 8678 21138 8730
rect 21190 8678 21202 8730
rect 21254 8678 21266 8730
rect 21318 8678 27010 8730
rect 27062 8678 27074 8730
rect 27126 8678 27138 8730
rect 27190 8678 27202 8730
rect 27254 8678 27266 8730
rect 27318 8678 32568 8730
rect 1104 8656 32568 8678
rect 1210 8576 1216 8628
rect 1268 8616 1274 8628
rect 1397 8619 1455 8625
rect 1397 8616 1409 8619
rect 1268 8588 1409 8616
rect 1268 8576 1274 8588
rect 1397 8585 1409 8588
rect 1443 8585 1455 8619
rect 1397 8579 1455 8585
rect 2774 8576 2780 8628
rect 2832 8616 2838 8628
rect 2961 8619 3019 8625
rect 2961 8616 2973 8619
rect 2832 8588 2973 8616
rect 2832 8576 2838 8588
rect 2961 8585 2973 8588
rect 3007 8585 3019 8619
rect 2961 8579 3019 8585
rect 4338 8576 4344 8628
rect 4396 8616 4402 8628
rect 4525 8619 4583 8625
rect 4525 8616 4537 8619
rect 4396 8588 4537 8616
rect 4396 8576 4402 8588
rect 4525 8585 4537 8588
rect 4571 8585 4583 8619
rect 4525 8579 4583 8585
rect 4706 8576 4712 8628
rect 4764 8576 4770 8628
rect 5902 8576 5908 8628
rect 5960 8616 5966 8628
rect 6457 8619 6515 8625
rect 6457 8616 6469 8619
rect 5960 8588 6469 8616
rect 5960 8576 5966 8588
rect 6457 8585 6469 8588
rect 6503 8585 6515 8619
rect 6457 8579 6515 8585
rect 7466 8576 7472 8628
rect 7524 8616 7530 8628
rect 7653 8619 7711 8625
rect 7653 8616 7665 8619
rect 7524 8588 7665 8616
rect 7524 8576 7530 8588
rect 7653 8585 7665 8588
rect 7699 8585 7711 8619
rect 7653 8579 7711 8585
rect 8846 8576 8852 8628
rect 8904 8616 8910 8628
rect 9217 8619 9275 8625
rect 9217 8616 9229 8619
rect 8904 8588 9229 8616
rect 8904 8576 8910 8588
rect 9217 8585 9229 8588
rect 9263 8585 9275 8619
rect 9217 8579 9275 8585
rect 10594 8576 10600 8628
rect 10652 8616 10658 8628
rect 10781 8619 10839 8625
rect 10781 8616 10793 8619
rect 10652 8588 10793 8616
rect 10652 8576 10658 8588
rect 10781 8585 10793 8588
rect 10827 8585 10839 8619
rect 12066 8616 12072 8628
rect 10781 8579 10839 8585
rect 10888 8588 12072 8616
rect 1578 8440 1584 8492
rect 1636 8440 1642 8492
rect 4724 8489 4752 8576
rect 10888 8548 10916 8588
rect 12066 8576 12072 8588
rect 12124 8576 12130 8628
rect 12158 8576 12164 8628
rect 12216 8616 12222 8628
rect 12345 8619 12403 8625
rect 12345 8616 12357 8619
rect 12216 8588 12357 8616
rect 12216 8576 12222 8588
rect 12345 8585 12357 8588
rect 12391 8585 12403 8619
rect 12345 8579 12403 8585
rect 13722 8576 13728 8628
rect 13780 8616 13786 8628
rect 14185 8619 14243 8625
rect 14185 8616 14197 8619
rect 13780 8588 14197 8616
rect 13780 8576 13786 8588
rect 14185 8585 14197 8588
rect 14231 8585 14243 8619
rect 14185 8579 14243 8585
rect 15378 8576 15384 8628
rect 15436 8616 15442 8628
rect 15473 8619 15531 8625
rect 15473 8616 15485 8619
rect 15436 8588 15485 8616
rect 15436 8576 15442 8588
rect 15473 8585 15485 8588
rect 15519 8585 15531 8619
rect 15473 8579 15531 8585
rect 16850 8576 16856 8628
rect 16908 8616 16914 8628
rect 17037 8619 17095 8625
rect 17037 8616 17049 8619
rect 16908 8588 17049 8616
rect 16908 8576 16914 8588
rect 17037 8585 17049 8588
rect 17083 8585 17095 8619
rect 17037 8579 17095 8585
rect 18414 8576 18420 8628
rect 18472 8616 18478 8628
rect 18601 8619 18659 8625
rect 18601 8616 18613 8619
rect 18472 8588 18613 8616
rect 18472 8576 18478 8588
rect 18601 8585 18613 8588
rect 18647 8585 18659 8619
rect 18601 8579 18659 8585
rect 19978 8576 19984 8628
rect 20036 8616 20042 8628
rect 20165 8619 20223 8625
rect 20165 8616 20177 8619
rect 20036 8588 20177 8616
rect 20036 8576 20042 8588
rect 20165 8585 20177 8588
rect 20211 8585 20223 8619
rect 20165 8579 20223 8585
rect 21542 8576 21548 8628
rect 21600 8616 21606 8628
rect 21913 8619 21971 8625
rect 21913 8616 21925 8619
rect 21600 8588 21925 8616
rect 21600 8576 21606 8588
rect 21913 8585 21925 8588
rect 21959 8585 21971 8619
rect 21913 8579 21971 8585
rect 23106 8576 23112 8628
rect 23164 8616 23170 8628
rect 23385 8619 23443 8625
rect 23385 8616 23397 8619
rect 23164 8588 23397 8616
rect 23164 8576 23170 8588
rect 23385 8585 23397 8588
rect 23431 8585 23443 8619
rect 23385 8579 23443 8585
rect 24670 8576 24676 8628
rect 24728 8616 24734 8628
rect 24949 8619 25007 8625
rect 24949 8616 24961 8619
rect 24728 8588 24961 8616
rect 24728 8576 24734 8588
rect 24949 8585 24961 8588
rect 24995 8585 25007 8619
rect 24949 8579 25007 8585
rect 26234 8576 26240 8628
rect 26292 8616 26298 8628
rect 26513 8619 26571 8625
rect 26513 8616 26525 8619
rect 26292 8588 26525 8616
rect 26292 8576 26298 8588
rect 26513 8585 26525 8588
rect 26559 8585 26571 8619
rect 26513 8579 26571 8585
rect 27798 8576 27804 8628
rect 27856 8616 27862 8628
rect 28077 8619 28135 8625
rect 28077 8616 28089 8619
rect 27856 8588 28089 8616
rect 27856 8576 27862 8588
rect 28077 8585 28089 8588
rect 28123 8585 28135 8619
rect 28077 8579 28135 8585
rect 29362 8576 29368 8628
rect 29420 8616 29426 8628
rect 29733 8619 29791 8625
rect 29733 8616 29745 8619
rect 29420 8588 29745 8616
rect 29420 8576 29426 8588
rect 29733 8585 29745 8588
rect 29779 8585 29791 8619
rect 29733 8579 29791 8585
rect 30098 8576 30104 8628
rect 30156 8576 30162 8628
rect 30466 8576 30472 8628
rect 30524 8576 30530 8628
rect 30926 8576 30932 8628
rect 30984 8616 30990 8628
rect 31205 8619 31263 8625
rect 31205 8616 31217 8619
rect 30984 8588 31217 8616
rect 30984 8576 30990 8588
rect 31205 8585 31217 8588
rect 31251 8585 31263 8619
rect 31205 8579 31263 8585
rect 19150 8548 19156 8560
rect 7852 8520 10916 8548
rect 17052 8520 19156 8548
rect 7852 8489 7880 8520
rect 3145 8483 3203 8489
rect 3145 8449 3157 8483
rect 3191 8449 3203 8483
rect 3145 8443 3203 8449
rect 4709 8483 4767 8489
rect 4709 8449 4721 8483
rect 4755 8449 4767 8483
rect 4709 8443 4767 8449
rect 6641 8483 6699 8489
rect 6641 8449 6653 8483
rect 6687 8480 6699 8483
rect 7837 8483 7895 8489
rect 6687 8452 6914 8480
rect 6687 8449 6699 8452
rect 6641 8443 6699 8449
rect 3160 8412 3188 8443
rect 4982 8412 4988 8424
rect 3160 8384 4988 8412
rect 4982 8372 4988 8384
rect 5040 8372 5046 8424
rect 6886 8412 6914 8452
rect 7837 8449 7849 8483
rect 7883 8449 7895 8483
rect 7837 8443 7895 8449
rect 9398 8440 9404 8492
rect 9456 8440 9462 8492
rect 10962 8440 10968 8492
rect 11020 8440 11026 8492
rect 12526 8440 12532 8492
rect 12584 8440 12590 8492
rect 14366 8440 14372 8492
rect 14424 8440 14430 8492
rect 15654 8489 15660 8492
rect 15650 8443 15660 8489
rect 15654 8440 15660 8443
rect 15712 8440 15718 8492
rect 17052 8480 17080 8520
rect 19150 8508 19156 8520
rect 19208 8508 19214 8560
rect 21376 8520 31708 8548
rect 15764 8452 17080 8480
rect 17221 8483 17279 8489
rect 15764 8412 15792 8452
rect 17221 8449 17233 8483
rect 17267 8449 17279 8483
rect 17221 8443 17279 8449
rect 6886 8384 15792 8412
rect 15838 8372 15844 8424
rect 15896 8412 15902 8424
rect 17034 8412 17040 8424
rect 15896 8384 17040 8412
rect 15896 8372 15902 8384
rect 17034 8372 17040 8384
rect 17092 8372 17098 8424
rect 17236 8412 17264 8443
rect 18782 8440 18788 8492
rect 18840 8440 18846 8492
rect 20346 8440 20352 8492
rect 20404 8440 20410 8492
rect 20530 8412 20536 8424
rect 17236 8384 20536 8412
rect 20530 8372 20536 8384
rect 20588 8372 20594 8424
rect 14918 8304 14924 8356
rect 14976 8344 14982 8356
rect 21376 8344 21404 8520
rect 22097 8483 22155 8489
rect 22097 8449 22109 8483
rect 22143 8480 22155 8483
rect 22186 8480 22192 8492
rect 22143 8452 22192 8480
rect 22143 8449 22155 8452
rect 22097 8443 22155 8449
rect 22186 8440 22192 8452
rect 22244 8440 22250 8492
rect 23106 8440 23112 8492
rect 23164 8480 23170 8492
rect 23201 8483 23259 8489
rect 23201 8480 23213 8483
rect 23164 8452 23213 8480
rect 23164 8440 23170 8452
rect 23201 8449 23213 8452
rect 23247 8449 23259 8483
rect 23201 8443 23259 8449
rect 23658 8440 23664 8492
rect 23716 8480 23722 8492
rect 24765 8483 24823 8489
rect 24765 8480 24777 8483
rect 23716 8452 24777 8480
rect 23716 8440 23722 8452
rect 24765 8449 24777 8452
rect 24811 8449 24823 8483
rect 24765 8443 24823 8449
rect 26329 8483 26387 8489
rect 26329 8449 26341 8483
rect 26375 8480 26387 8483
rect 26418 8480 26424 8492
rect 26375 8452 26424 8480
rect 26375 8449 26387 8452
rect 26329 8443 26387 8449
rect 26418 8440 26424 8452
rect 26476 8440 26482 8492
rect 27893 8483 27951 8489
rect 27893 8449 27905 8483
rect 27939 8449 27951 8483
rect 27893 8443 27951 8449
rect 25038 8372 25044 8424
rect 25096 8412 25102 8424
rect 27908 8412 27936 8443
rect 28994 8440 29000 8492
rect 29052 8480 29058 8492
rect 29549 8483 29607 8489
rect 29549 8480 29561 8483
rect 29052 8452 29561 8480
rect 29052 8440 29058 8452
rect 29549 8449 29561 8452
rect 29595 8449 29607 8483
rect 29549 8443 29607 8449
rect 29914 8440 29920 8492
rect 29972 8440 29978 8492
rect 30282 8440 30288 8492
rect 30340 8440 30346 8492
rect 30650 8440 30656 8492
rect 30708 8440 30714 8492
rect 31680 8489 31708 8520
rect 31021 8483 31079 8489
rect 31021 8449 31033 8483
rect 31067 8449 31079 8483
rect 31021 8443 31079 8449
rect 31665 8483 31723 8489
rect 31665 8449 31677 8483
rect 31711 8449 31723 8483
rect 31665 8443 31723 8449
rect 25096 8384 27936 8412
rect 25096 8372 25102 8384
rect 30466 8372 30472 8424
rect 30524 8412 30530 8424
rect 31036 8412 31064 8443
rect 32398 8412 32404 8424
rect 30524 8384 31064 8412
rect 31726 8384 32404 8412
rect 30524 8372 30530 8384
rect 14976 8316 21404 8344
rect 30837 8347 30895 8353
rect 14976 8304 14982 8316
rect 30837 8313 30849 8347
rect 30883 8344 30895 8347
rect 31726 8344 31754 8384
rect 32398 8372 32404 8384
rect 32456 8372 32462 8424
rect 30883 8316 31754 8344
rect 30883 8313 30895 8316
rect 30837 8307 30895 8313
rect 31846 8304 31852 8356
rect 31904 8304 31910 8356
rect 1104 8186 32568 8208
rect 1104 8134 1950 8186
rect 2002 8134 2014 8186
rect 2066 8134 2078 8186
rect 2130 8134 2142 8186
rect 2194 8134 2206 8186
rect 2258 8134 7950 8186
rect 8002 8134 8014 8186
rect 8066 8134 8078 8186
rect 8130 8134 8142 8186
rect 8194 8134 8206 8186
rect 8258 8134 13950 8186
rect 14002 8134 14014 8186
rect 14066 8134 14078 8186
rect 14130 8134 14142 8186
rect 14194 8134 14206 8186
rect 14258 8134 19950 8186
rect 20002 8134 20014 8186
rect 20066 8134 20078 8186
rect 20130 8134 20142 8186
rect 20194 8134 20206 8186
rect 20258 8134 25950 8186
rect 26002 8134 26014 8186
rect 26066 8134 26078 8186
rect 26130 8134 26142 8186
rect 26194 8134 26206 8186
rect 26258 8134 31950 8186
rect 32002 8134 32014 8186
rect 32066 8134 32078 8186
rect 32130 8134 32142 8186
rect 32194 8134 32206 8186
rect 32258 8134 32568 8186
rect 1104 8112 32568 8134
rect 15562 8072 15568 8084
rect 6886 8044 15568 8072
rect 4890 7964 4896 8016
rect 4948 8004 4954 8016
rect 6886 8004 6914 8044
rect 15562 8032 15568 8044
rect 15620 8032 15626 8084
rect 21634 8032 21640 8084
rect 21692 8072 21698 8084
rect 30374 8072 30380 8084
rect 21692 8044 30380 8072
rect 21692 8032 21698 8044
rect 30374 8032 30380 8044
rect 30432 8032 30438 8084
rect 30653 8075 30711 8081
rect 30653 8041 30665 8075
rect 30699 8072 30711 8075
rect 30834 8072 30840 8084
rect 30699 8044 30840 8072
rect 30699 8041 30711 8044
rect 30653 8035 30711 8041
rect 30834 8032 30840 8044
rect 30892 8032 30898 8084
rect 31018 8032 31024 8084
rect 31076 8032 31082 8084
rect 31386 8032 31392 8084
rect 31444 8032 31450 8084
rect 4948 7976 6914 8004
rect 4948 7964 4954 7976
rect 7006 7964 7012 8016
rect 7064 8004 7070 8016
rect 7064 7976 15608 8004
rect 7064 7964 7070 7976
rect 7650 7896 7656 7948
rect 7708 7936 7714 7948
rect 13354 7936 13360 7948
rect 7708 7908 13360 7936
rect 7708 7896 7714 7908
rect 13354 7896 13360 7908
rect 13412 7896 13418 7948
rect 7558 7828 7564 7880
rect 7616 7868 7622 7880
rect 15470 7868 15476 7880
rect 7616 7840 15476 7868
rect 7616 7828 7622 7840
rect 15470 7828 15476 7840
rect 15528 7828 15534 7880
rect 7374 7760 7380 7812
rect 7432 7800 7438 7812
rect 12158 7800 12164 7812
rect 7432 7772 12164 7800
rect 7432 7760 7438 7772
rect 12158 7760 12164 7772
rect 12216 7760 12222 7812
rect 15580 7800 15608 7976
rect 19150 7964 19156 8016
rect 19208 8004 19214 8016
rect 20254 8004 20260 8016
rect 19208 7976 20260 8004
rect 19208 7964 19214 7976
rect 20254 7964 20260 7976
rect 20312 7964 20318 8016
rect 26786 7964 26792 8016
rect 26844 8004 26850 8016
rect 26844 7976 31616 8004
rect 26844 7964 26850 7976
rect 16390 7896 16396 7948
rect 16448 7936 16454 7948
rect 16448 7908 31248 7936
rect 16448 7896 16454 7908
rect 18138 7828 18144 7880
rect 18196 7868 18202 7880
rect 21634 7868 21640 7880
rect 18196 7840 21640 7868
rect 18196 7828 18202 7840
rect 21634 7828 21640 7840
rect 21692 7828 21698 7880
rect 23934 7828 23940 7880
rect 23992 7868 23998 7880
rect 30469 7871 30527 7877
rect 30469 7868 30481 7871
rect 23992 7840 30481 7868
rect 23992 7828 23998 7840
rect 30469 7837 30481 7840
rect 30515 7837 30527 7871
rect 30469 7831 30527 7837
rect 30834 7828 30840 7880
rect 30892 7828 30898 7880
rect 31220 7877 31248 7908
rect 31588 7877 31616 7976
rect 31205 7871 31263 7877
rect 31205 7837 31217 7871
rect 31251 7837 31263 7871
rect 31205 7831 31263 7837
rect 31573 7871 31631 7877
rect 31573 7837 31585 7871
rect 31619 7837 31631 7871
rect 31573 7831 31631 7837
rect 31941 7871 31999 7877
rect 31941 7837 31953 7871
rect 31987 7837 31999 7871
rect 31941 7831 31999 7837
rect 31956 7800 31984 7831
rect 15580 7772 31984 7800
rect 5626 7692 5632 7744
rect 5684 7732 5690 7744
rect 8110 7732 8116 7744
rect 5684 7704 8116 7732
rect 5684 7692 5690 7704
rect 8110 7692 8116 7704
rect 8168 7692 8174 7744
rect 12066 7692 12072 7744
rect 12124 7732 12130 7744
rect 14274 7732 14280 7744
rect 12124 7704 14280 7732
rect 12124 7692 12130 7704
rect 14274 7692 14280 7704
rect 14332 7692 14338 7744
rect 16850 7692 16856 7744
rect 16908 7732 16914 7744
rect 26786 7732 26792 7744
rect 16908 7704 26792 7732
rect 16908 7692 16914 7704
rect 26786 7692 26792 7704
rect 26844 7692 26850 7744
rect 31754 7692 31760 7744
rect 31812 7692 31818 7744
rect 32122 7692 32128 7744
rect 32180 7692 32186 7744
rect 1104 7642 32568 7664
rect 1104 7590 3010 7642
rect 3062 7590 3074 7642
rect 3126 7590 3138 7642
rect 3190 7590 3202 7642
rect 3254 7590 3266 7642
rect 3318 7590 9010 7642
rect 9062 7590 9074 7642
rect 9126 7590 9138 7642
rect 9190 7590 9202 7642
rect 9254 7590 9266 7642
rect 9318 7590 15010 7642
rect 15062 7590 15074 7642
rect 15126 7590 15138 7642
rect 15190 7590 15202 7642
rect 15254 7590 15266 7642
rect 15318 7590 21010 7642
rect 21062 7590 21074 7642
rect 21126 7590 21138 7642
rect 21190 7590 21202 7642
rect 21254 7590 21266 7642
rect 21318 7590 27010 7642
rect 27062 7590 27074 7642
rect 27126 7590 27138 7642
rect 27190 7590 27202 7642
rect 27254 7590 27266 7642
rect 27318 7590 32568 7642
rect 1104 7568 32568 7590
rect 4890 7488 4896 7540
rect 4948 7488 4954 7540
rect 6086 7488 6092 7540
rect 6144 7528 6150 7540
rect 6733 7531 6791 7537
rect 6144 7500 6684 7528
rect 6144 7488 6150 7500
rect 5534 7420 5540 7472
rect 5592 7460 5598 7472
rect 6656 7460 6684 7500
rect 6733 7497 6745 7531
rect 6779 7528 6791 7531
rect 7558 7528 7564 7540
rect 6779 7500 7564 7528
rect 6779 7497 6791 7500
rect 6733 7491 6791 7497
rect 7558 7488 7564 7500
rect 7616 7488 7622 7540
rect 7653 7531 7711 7537
rect 7653 7497 7665 7531
rect 7699 7528 7711 7531
rect 12618 7528 12624 7540
rect 7699 7500 12624 7528
rect 7699 7497 7711 7500
rect 7653 7491 7711 7497
rect 12618 7488 12624 7500
rect 12676 7488 12682 7540
rect 13354 7488 13360 7540
rect 13412 7488 13418 7540
rect 13722 7488 13728 7540
rect 13780 7528 13786 7540
rect 15289 7531 15347 7537
rect 15289 7528 15301 7531
rect 13780 7500 15301 7528
rect 13780 7488 13786 7500
rect 15289 7497 15301 7500
rect 15335 7497 15347 7531
rect 15289 7491 15347 7497
rect 15378 7488 15384 7540
rect 15436 7528 15442 7540
rect 16025 7531 16083 7537
rect 16025 7528 16037 7531
rect 15436 7500 16037 7528
rect 15436 7488 15442 7500
rect 16025 7497 16037 7500
rect 16071 7497 16083 7531
rect 16025 7491 16083 7497
rect 16390 7488 16396 7540
rect 16448 7488 16454 7540
rect 16574 7488 16580 7540
rect 16632 7528 16638 7540
rect 17773 7531 17831 7537
rect 17773 7528 17785 7531
rect 16632 7500 17785 7528
rect 16632 7488 16638 7500
rect 17773 7497 17785 7500
rect 17819 7497 17831 7531
rect 17773 7491 17831 7497
rect 18138 7488 18144 7540
rect 18196 7488 18202 7540
rect 19705 7531 19763 7537
rect 19705 7497 19717 7531
rect 19751 7497 19763 7531
rect 19705 7491 19763 7497
rect 5592 7432 6592 7460
rect 6656 7432 7512 7460
rect 5592 7420 5598 7432
rect 4706 7352 4712 7404
rect 4764 7352 4770 7404
rect 4798 7352 4804 7404
rect 4856 7392 4862 7404
rect 6564 7401 6592 7432
rect 5721 7395 5779 7401
rect 5721 7392 5733 7395
rect 4856 7364 5733 7392
rect 4856 7352 4862 7364
rect 5721 7361 5733 7364
rect 5767 7361 5779 7395
rect 5721 7355 5779 7361
rect 5997 7395 6055 7401
rect 5997 7361 6009 7395
rect 6043 7361 6055 7395
rect 5997 7355 6055 7361
rect 6549 7395 6607 7401
rect 6549 7361 6561 7395
rect 6595 7361 6607 7395
rect 6549 7355 6607 7361
rect 6012 7324 6040 7355
rect 6822 7352 6828 7404
rect 6880 7352 6886 7404
rect 7484 7401 7512 7432
rect 8110 7420 8116 7472
rect 8168 7460 8174 7472
rect 13449 7463 13507 7469
rect 8168 7432 9352 7460
rect 8168 7420 8174 7432
rect 9324 7401 9352 7432
rect 13449 7429 13461 7463
rect 13495 7460 13507 7463
rect 13495 7432 13860 7460
rect 13495 7429 13507 7432
rect 13449 7423 13507 7429
rect 7193 7395 7251 7401
rect 7193 7361 7205 7395
rect 7239 7361 7251 7395
rect 7193 7355 7251 7361
rect 7469 7395 7527 7401
rect 7469 7361 7481 7395
rect 7515 7361 7527 7395
rect 7469 7355 7527 7361
rect 8757 7395 8815 7401
rect 8757 7361 8769 7395
rect 8803 7361 8815 7395
rect 9033 7395 9091 7401
rect 9033 7392 9045 7395
rect 8757 7355 8815 7361
rect 8864 7364 9045 7392
rect 7098 7324 7104 7336
rect 6012 7296 7104 7324
rect 7098 7284 7104 7296
rect 7156 7284 7162 7336
rect 7208 7324 7236 7355
rect 7834 7324 7840 7336
rect 7208 7296 7840 7324
rect 7834 7284 7840 7296
rect 7892 7284 7898 7336
rect 5902 7216 5908 7268
rect 5960 7216 5966 7268
rect 6270 7216 6276 7268
rect 6328 7256 6334 7268
rect 8772 7256 8800 7355
rect 6328 7228 8800 7256
rect 6328 7216 6334 7228
rect 6178 7148 6184 7200
rect 6236 7148 6242 7200
rect 7006 7148 7012 7200
rect 7064 7148 7070 7200
rect 7374 7148 7380 7200
rect 7432 7148 7438 7200
rect 7742 7148 7748 7200
rect 7800 7188 7806 7200
rect 8864 7188 8892 7364
rect 9033 7361 9045 7364
rect 9079 7361 9091 7395
rect 9033 7355 9091 7361
rect 9309 7395 9367 7401
rect 9309 7361 9321 7395
rect 9355 7361 9367 7395
rect 9309 7355 9367 7361
rect 11882 7352 11888 7404
rect 11940 7352 11946 7404
rect 12158 7352 12164 7404
rect 12216 7352 12222 7404
rect 12434 7352 12440 7404
rect 12492 7352 12498 7404
rect 12805 7395 12863 7401
rect 12805 7361 12817 7395
rect 12851 7392 12863 7395
rect 12897 7395 12955 7401
rect 12897 7392 12909 7395
rect 12851 7364 12909 7392
rect 12851 7361 12863 7364
rect 12805 7355 12863 7361
rect 12897 7361 12909 7364
rect 12943 7361 12955 7395
rect 12897 7355 12955 7361
rect 13633 7395 13691 7401
rect 13633 7361 13645 7395
rect 13679 7392 13691 7395
rect 13725 7395 13783 7401
rect 13725 7392 13737 7395
rect 13679 7364 13737 7392
rect 13679 7361 13691 7364
rect 13633 7355 13691 7361
rect 13725 7361 13737 7364
rect 13771 7361 13783 7395
rect 13832 7392 13860 7432
rect 13906 7420 13912 7472
rect 13964 7460 13970 7472
rect 13964 7432 16712 7460
rect 13964 7420 13970 7432
rect 14458 7401 14464 7404
rect 14001 7395 14059 7401
rect 14001 7392 14013 7395
rect 13832 7364 14013 7392
rect 13725 7355 13783 7361
rect 14001 7361 14013 7364
rect 14047 7361 14059 7395
rect 14437 7395 14464 7401
rect 14437 7392 14449 7395
rect 14001 7355 14059 7361
rect 14108 7364 14449 7392
rect 13265 7327 13323 7333
rect 13265 7293 13277 7327
rect 13311 7324 13323 7327
rect 14108 7324 14136 7364
rect 14437 7361 14449 7364
rect 14437 7355 14464 7361
rect 14458 7352 14464 7355
rect 14516 7352 14522 7404
rect 14550 7352 14556 7404
rect 14608 7392 14614 7404
rect 14737 7395 14795 7401
rect 14737 7392 14749 7395
rect 14608 7364 14749 7392
rect 14608 7352 14614 7364
rect 14737 7361 14749 7364
rect 14783 7361 14795 7395
rect 14737 7355 14795 7361
rect 15013 7395 15071 7401
rect 15013 7361 15025 7395
rect 15059 7392 15071 7395
rect 15289 7395 15347 7401
rect 15289 7392 15301 7395
rect 15059 7364 15301 7392
rect 15059 7361 15071 7364
rect 15013 7355 15071 7361
rect 15289 7361 15301 7364
rect 15335 7361 15347 7395
rect 15289 7355 15347 7361
rect 16117 7395 16175 7401
rect 16117 7361 16129 7395
rect 16163 7392 16175 7395
rect 16209 7395 16267 7401
rect 16209 7392 16221 7395
rect 16163 7364 16221 7392
rect 16163 7361 16175 7364
rect 16117 7355 16175 7361
rect 16209 7361 16221 7364
rect 16255 7361 16267 7395
rect 16209 7355 16267 7361
rect 16298 7352 16304 7404
rect 16356 7392 16362 7404
rect 16684 7401 16712 7432
rect 17126 7420 17132 7472
rect 17184 7420 17190 7472
rect 19518 7420 19524 7472
rect 19576 7460 19582 7472
rect 19720 7460 19748 7491
rect 20254 7488 20260 7540
rect 20312 7488 20318 7540
rect 21634 7528 21640 7540
rect 20456 7500 21640 7528
rect 19576 7432 19748 7460
rect 19576 7420 19582 7432
rect 16669 7395 16727 7401
rect 16356 7364 16574 7392
rect 16356 7352 16362 7364
rect 16390 7324 16396 7336
rect 13311 7296 14136 7324
rect 15120 7296 16396 7324
rect 13311 7293 13323 7296
rect 13265 7287 13323 7293
rect 8941 7259 8999 7265
rect 8941 7225 8953 7259
rect 8987 7256 8999 7259
rect 9306 7256 9312 7268
rect 8987 7228 9312 7256
rect 8987 7225 8999 7228
rect 8941 7219 8999 7225
rect 9306 7216 9312 7228
rect 9364 7216 9370 7268
rect 10962 7216 10968 7268
rect 11020 7256 11026 7268
rect 13541 7259 13599 7265
rect 13541 7256 13553 7259
rect 11020 7228 13553 7256
rect 11020 7216 11026 7228
rect 13541 7225 13553 7228
rect 13587 7225 13599 7259
rect 13541 7219 13599 7225
rect 13909 7259 13967 7265
rect 13909 7225 13921 7259
rect 13955 7256 13967 7259
rect 15120 7256 15148 7296
rect 16390 7284 16396 7296
rect 16448 7284 16454 7336
rect 16546 7324 16574 7364
rect 16669 7361 16681 7395
rect 16715 7392 16727 7395
rect 16945 7395 17003 7401
rect 16945 7392 16957 7395
rect 16715 7364 16957 7392
rect 16715 7361 16727 7364
rect 16669 7355 16727 7361
rect 16945 7361 16957 7364
rect 16991 7361 17003 7395
rect 16945 7355 17003 7361
rect 17221 7395 17279 7401
rect 17221 7361 17233 7395
rect 17267 7392 17279 7395
rect 17313 7395 17371 7401
rect 17313 7392 17325 7395
rect 17267 7364 17325 7392
rect 17267 7361 17279 7364
rect 17221 7355 17279 7361
rect 17313 7361 17325 7364
rect 17359 7361 17371 7395
rect 17313 7355 17371 7361
rect 17865 7395 17923 7401
rect 17865 7361 17877 7395
rect 17911 7392 17923 7395
rect 17957 7395 18015 7401
rect 17957 7392 17969 7395
rect 17911 7364 17969 7392
rect 17911 7361 17923 7364
rect 17865 7355 17923 7361
rect 17957 7361 17969 7364
rect 18003 7361 18015 7395
rect 17957 7355 18015 7361
rect 19610 7352 19616 7404
rect 19668 7392 19674 7404
rect 20456 7401 20484 7500
rect 21634 7488 21640 7500
rect 21692 7488 21698 7540
rect 22922 7488 22928 7540
rect 22980 7488 22986 7540
rect 24210 7488 24216 7540
rect 24268 7488 24274 7540
rect 25130 7488 25136 7540
rect 25188 7488 25194 7540
rect 25314 7488 25320 7540
rect 25372 7488 25378 7540
rect 31478 7488 31484 7540
rect 31536 7488 31542 7540
rect 25682 7460 25688 7472
rect 23124 7432 25688 7460
rect 19889 7395 19947 7401
rect 19889 7392 19901 7395
rect 19668 7364 19901 7392
rect 19668 7352 19674 7364
rect 19889 7361 19901 7364
rect 19935 7361 19947 7395
rect 19889 7355 19947 7361
rect 20441 7395 20499 7401
rect 20441 7361 20453 7395
rect 20487 7361 20499 7395
rect 20441 7355 20499 7361
rect 20898 7352 20904 7404
rect 20956 7352 20962 7404
rect 23124 7401 23152 7432
rect 25682 7420 25688 7432
rect 25740 7420 25746 7472
rect 23109 7395 23167 7401
rect 23109 7361 23121 7395
rect 23155 7361 23167 7395
rect 23109 7355 23167 7361
rect 24302 7352 24308 7404
rect 24360 7392 24366 7404
rect 24397 7395 24455 7401
rect 24397 7392 24409 7395
rect 24360 7364 24409 7392
rect 24360 7352 24366 7364
rect 24397 7361 24409 7364
rect 24443 7361 24455 7395
rect 24397 7355 24455 7361
rect 24949 7395 25007 7401
rect 24949 7361 24961 7395
rect 24995 7361 25007 7395
rect 24949 7355 25007 7361
rect 25501 7395 25559 7401
rect 25501 7361 25513 7395
rect 25547 7392 25559 7395
rect 25866 7392 25872 7404
rect 25547 7364 25872 7392
rect 25547 7361 25559 7364
rect 25501 7355 25559 7361
rect 23934 7324 23940 7336
rect 16546 7296 23940 7324
rect 23934 7284 23940 7296
rect 23992 7284 23998 7336
rect 24026 7284 24032 7336
rect 24084 7324 24090 7336
rect 24964 7324 24992 7355
rect 25866 7352 25872 7364
rect 25924 7352 25930 7404
rect 31294 7352 31300 7404
rect 31352 7352 31358 7404
rect 31665 7395 31723 7401
rect 31665 7361 31677 7395
rect 31711 7361 31723 7395
rect 31665 7355 31723 7361
rect 24084 7296 24992 7324
rect 24084 7284 24090 7296
rect 13955 7228 15148 7256
rect 15197 7259 15255 7265
rect 13955 7225 13967 7228
rect 13909 7219 13967 7225
rect 15197 7225 15209 7259
rect 15243 7256 15255 7259
rect 15378 7256 15384 7268
rect 15243 7228 15384 7256
rect 15243 7225 15255 7228
rect 15197 7219 15255 7225
rect 15378 7216 15384 7228
rect 15436 7216 15442 7268
rect 15470 7216 15476 7268
rect 15528 7256 15534 7268
rect 31680 7256 31708 7355
rect 15528 7228 31708 7256
rect 15528 7216 15534 7228
rect 7800 7160 8892 7188
rect 7800 7148 7806 7160
rect 9214 7148 9220 7200
rect 9272 7148 9278 7200
rect 9490 7148 9496 7200
rect 9548 7148 9554 7200
rect 12066 7148 12072 7200
rect 12124 7148 12130 7200
rect 12342 7148 12348 7200
rect 12400 7148 12406 7200
rect 12526 7148 12532 7200
rect 12584 7188 12590 7200
rect 12621 7191 12679 7197
rect 12621 7188 12633 7191
rect 12584 7160 12633 7188
rect 12584 7148 12590 7160
rect 12621 7157 12633 7160
rect 12667 7157 12679 7191
rect 12621 7151 12679 7157
rect 12710 7148 12716 7200
rect 12768 7148 12774 7200
rect 13078 7148 13084 7200
rect 13136 7148 13142 7200
rect 14182 7148 14188 7200
rect 14240 7148 14246 7200
rect 14274 7148 14280 7200
rect 14332 7148 14338 7200
rect 14918 7148 14924 7200
rect 14976 7148 14982 7200
rect 16850 7148 16856 7200
rect 16908 7148 16914 7200
rect 17494 7148 17500 7200
rect 17552 7148 17558 7200
rect 17862 7148 17868 7200
rect 17920 7188 17926 7200
rect 20717 7191 20775 7197
rect 20717 7188 20729 7191
rect 17920 7160 20729 7188
rect 17920 7148 17926 7160
rect 20717 7157 20729 7160
rect 20763 7157 20775 7191
rect 20717 7151 20775 7157
rect 31849 7191 31907 7197
rect 31849 7157 31861 7191
rect 31895 7188 31907 7191
rect 32766 7188 32772 7200
rect 31895 7160 32772 7188
rect 31895 7157 31907 7160
rect 31849 7151 31907 7157
rect 32766 7148 32772 7160
rect 32824 7148 32830 7200
rect 1104 7098 32568 7120
rect 1104 7046 1950 7098
rect 2002 7046 2014 7098
rect 2066 7046 2078 7098
rect 2130 7046 2142 7098
rect 2194 7046 2206 7098
rect 2258 7046 7950 7098
rect 8002 7046 8014 7098
rect 8066 7046 8078 7098
rect 8130 7046 8142 7098
rect 8194 7046 8206 7098
rect 8258 7046 13950 7098
rect 14002 7046 14014 7098
rect 14066 7046 14078 7098
rect 14130 7046 14142 7098
rect 14194 7046 14206 7098
rect 14258 7046 19950 7098
rect 20002 7046 20014 7098
rect 20066 7046 20078 7098
rect 20130 7046 20142 7098
rect 20194 7046 20206 7098
rect 20258 7046 25950 7098
rect 26002 7046 26014 7098
rect 26066 7046 26078 7098
rect 26130 7046 26142 7098
rect 26194 7046 26206 7098
rect 26258 7046 31950 7098
rect 32002 7046 32014 7098
rect 32066 7046 32078 7098
rect 32130 7046 32142 7098
rect 32194 7046 32206 7098
rect 32258 7046 32568 7098
rect 1104 7024 32568 7046
rect 4706 6944 4712 6996
rect 4764 6984 4770 6996
rect 7466 6984 7472 6996
rect 4764 6956 7472 6984
rect 4764 6944 4770 6956
rect 7466 6944 7472 6956
rect 7524 6944 7530 6996
rect 12342 6944 12348 6996
rect 12400 6984 12406 6996
rect 30834 6984 30840 6996
rect 12400 6956 30840 6984
rect 12400 6944 12406 6956
rect 30834 6944 30840 6956
rect 30892 6944 30898 6996
rect 7098 6876 7104 6928
rect 7156 6916 7162 6928
rect 7742 6916 7748 6928
rect 7156 6888 7748 6916
rect 7156 6876 7162 6888
rect 7742 6876 7748 6888
rect 7800 6876 7806 6928
rect 9214 6876 9220 6928
rect 9272 6916 9278 6928
rect 16298 6916 16304 6928
rect 9272 6888 16304 6916
rect 9272 6876 9278 6888
rect 16298 6876 16304 6888
rect 16356 6876 16362 6928
rect 20898 6876 20904 6928
rect 20956 6916 20962 6928
rect 24578 6916 24584 6928
rect 20956 6888 24584 6916
rect 20956 6876 20962 6888
rect 24578 6876 24584 6888
rect 24636 6876 24642 6928
rect 9306 6808 9312 6860
rect 9364 6848 9370 6860
rect 17034 6848 17040 6860
rect 9364 6820 17040 6848
rect 9364 6808 9370 6820
rect 17034 6808 17040 6820
rect 17092 6808 17098 6860
rect 17144 6820 31248 6848
rect 5721 6783 5779 6789
rect 5721 6749 5733 6783
rect 5767 6780 5779 6783
rect 5810 6780 5816 6792
rect 5767 6752 5816 6780
rect 5767 6749 5779 6752
rect 5721 6743 5779 6749
rect 5810 6740 5816 6752
rect 5868 6740 5874 6792
rect 8021 6783 8079 6789
rect 8021 6780 8033 6783
rect 5920 6752 8033 6780
rect 4706 6672 4712 6724
rect 4764 6712 4770 6724
rect 5920 6712 5948 6752
rect 8021 6749 8033 6752
rect 8067 6749 8079 6783
rect 8021 6743 8079 6749
rect 8294 6740 8300 6792
rect 8352 6780 8358 6792
rect 8389 6783 8447 6789
rect 8389 6780 8401 6783
rect 8352 6752 8401 6780
rect 8352 6740 8358 6752
rect 8389 6749 8401 6752
rect 8435 6749 8447 6783
rect 8389 6743 8447 6749
rect 8941 6783 8999 6789
rect 8941 6749 8953 6783
rect 8987 6749 8999 6783
rect 15562 6780 15568 6792
rect 8941 6743 8999 6749
rect 9048 6752 15568 6780
rect 4764 6684 5948 6712
rect 4764 6672 4770 6684
rect 6362 6672 6368 6724
rect 6420 6712 6426 6724
rect 8956 6712 8984 6743
rect 6420 6684 8984 6712
rect 6420 6672 6426 6684
rect 5902 6604 5908 6656
rect 5960 6604 5966 6656
rect 8202 6604 8208 6656
rect 8260 6604 8266 6656
rect 8573 6647 8631 6653
rect 8573 6613 8585 6647
rect 8619 6644 8631 6647
rect 9048 6644 9076 6752
rect 15562 6740 15568 6752
rect 15620 6740 15626 6792
rect 16482 6740 16488 6792
rect 16540 6780 16546 6792
rect 17144 6780 17172 6820
rect 16540 6752 17172 6780
rect 16540 6740 16546 6752
rect 17218 6740 17224 6792
rect 17276 6740 17282 6792
rect 19429 6783 19487 6789
rect 19429 6749 19441 6783
rect 19475 6780 19487 6783
rect 19521 6783 19579 6789
rect 19521 6780 19533 6783
rect 19475 6752 19533 6780
rect 19475 6749 19487 6752
rect 19429 6743 19487 6749
rect 19521 6749 19533 6752
rect 19567 6749 19579 6783
rect 19521 6743 19579 6749
rect 25317 6783 25375 6789
rect 25317 6749 25329 6783
rect 25363 6780 25375 6783
rect 26326 6780 26332 6792
rect 25363 6752 26332 6780
rect 25363 6749 25375 6752
rect 25317 6743 25375 6749
rect 26326 6740 26332 6752
rect 26384 6740 26390 6792
rect 31220 6789 31248 6820
rect 31205 6783 31263 6789
rect 31205 6749 31217 6783
rect 31251 6749 31263 6783
rect 31205 6743 31263 6749
rect 31570 6740 31576 6792
rect 31628 6740 31634 6792
rect 31662 6740 31668 6792
rect 31720 6780 31726 6792
rect 31941 6783 31999 6789
rect 31941 6780 31953 6783
rect 31720 6752 31953 6780
rect 31720 6740 31726 6752
rect 31941 6749 31953 6752
rect 31987 6749 31999 6783
rect 31941 6743 31999 6749
rect 9490 6672 9496 6724
rect 9548 6712 9554 6724
rect 31478 6712 31484 6724
rect 9548 6684 31484 6712
rect 9548 6672 9554 6684
rect 31478 6672 31484 6684
rect 31536 6672 31542 6724
rect 8619 6616 9076 6644
rect 9125 6647 9183 6653
rect 8619 6613 8631 6616
rect 8573 6607 8631 6613
rect 9125 6613 9137 6647
rect 9171 6644 9183 6647
rect 16114 6644 16120 6656
rect 9171 6616 16120 6644
rect 9171 6613 9183 6616
rect 9125 6607 9183 6613
rect 16114 6604 16120 6616
rect 16172 6604 16178 6656
rect 16942 6604 16948 6656
rect 17000 6644 17006 6656
rect 17037 6647 17095 6653
rect 17037 6644 17049 6647
rect 17000 6616 17049 6644
rect 17000 6604 17006 6616
rect 17037 6613 17049 6616
rect 17083 6644 17095 6647
rect 17218 6644 17224 6656
rect 17083 6616 17224 6644
rect 17083 6613 17095 6616
rect 17037 6607 17095 6613
rect 17218 6604 17224 6616
rect 17276 6604 17282 6656
rect 17405 6647 17463 6653
rect 17405 6613 17417 6647
rect 17451 6644 17463 6647
rect 19242 6644 19248 6656
rect 17451 6616 19248 6644
rect 17451 6613 17463 6616
rect 17405 6607 17463 6613
rect 19242 6604 19248 6616
rect 19300 6604 19306 6656
rect 19334 6604 19340 6656
rect 19392 6604 19398 6656
rect 19702 6604 19708 6656
rect 19760 6604 19766 6656
rect 24946 6604 24952 6656
rect 25004 6644 25010 6656
rect 25133 6647 25191 6653
rect 25133 6644 25145 6647
rect 25004 6616 25145 6644
rect 25004 6604 25010 6616
rect 25133 6613 25145 6616
rect 25179 6613 25191 6647
rect 25133 6607 25191 6613
rect 31386 6604 31392 6656
rect 31444 6604 31450 6656
rect 31754 6604 31760 6656
rect 31812 6604 31818 6656
rect 32125 6647 32183 6653
rect 32125 6613 32137 6647
rect 32171 6644 32183 6647
rect 32306 6644 32312 6656
rect 32171 6616 32312 6644
rect 32171 6613 32183 6616
rect 32125 6607 32183 6613
rect 32306 6604 32312 6616
rect 32364 6604 32370 6656
rect 1104 6554 32568 6576
rect 1104 6502 3010 6554
rect 3062 6502 3074 6554
rect 3126 6502 3138 6554
rect 3190 6502 3202 6554
rect 3254 6502 3266 6554
rect 3318 6502 9010 6554
rect 9062 6502 9074 6554
rect 9126 6502 9138 6554
rect 9190 6502 9202 6554
rect 9254 6502 9266 6554
rect 9318 6502 15010 6554
rect 15062 6502 15074 6554
rect 15126 6502 15138 6554
rect 15190 6502 15202 6554
rect 15254 6502 15266 6554
rect 15318 6502 21010 6554
rect 21062 6502 21074 6554
rect 21126 6502 21138 6554
rect 21190 6502 21202 6554
rect 21254 6502 21266 6554
rect 21318 6502 27010 6554
rect 27062 6502 27074 6554
rect 27126 6502 27138 6554
rect 27190 6502 27202 6554
rect 27254 6502 27266 6554
rect 27318 6502 32568 6554
rect 1104 6480 32568 6502
rect 8202 6400 8208 6452
rect 8260 6440 8266 6452
rect 14734 6440 14740 6452
rect 8260 6412 14740 6440
rect 8260 6400 8266 6412
rect 14734 6400 14740 6412
rect 14792 6400 14798 6452
rect 19702 6400 19708 6452
rect 19760 6440 19766 6452
rect 27614 6440 27620 6452
rect 19760 6412 27620 6440
rect 19760 6400 19766 6412
rect 27614 6400 27620 6412
rect 27672 6400 27678 6452
rect 31846 6400 31852 6452
rect 31904 6400 31910 6452
rect 17034 6332 17040 6384
rect 17092 6372 17098 6384
rect 31570 6372 31576 6384
rect 17092 6344 31576 6372
rect 17092 6332 17098 6344
rect 31570 6332 31576 6344
rect 31628 6332 31634 6384
rect 4430 6264 4436 6316
rect 4488 6304 4494 6316
rect 7193 6307 7251 6313
rect 7193 6304 7205 6307
rect 4488 6276 7205 6304
rect 4488 6264 4494 6276
rect 7193 6273 7205 6276
rect 7239 6273 7251 6307
rect 7193 6267 7251 6273
rect 8570 6264 8576 6316
rect 8628 6304 8634 6316
rect 9769 6307 9827 6313
rect 9769 6304 9781 6307
rect 8628 6276 9781 6304
rect 8628 6264 8634 6276
rect 9769 6273 9781 6276
rect 9815 6273 9827 6307
rect 9769 6267 9827 6273
rect 20625 6307 20683 6313
rect 20625 6273 20637 6307
rect 20671 6273 20683 6307
rect 20625 6267 20683 6273
rect 21085 6307 21143 6313
rect 21085 6273 21097 6307
rect 21131 6304 21143 6307
rect 21177 6307 21235 6313
rect 21177 6304 21189 6307
rect 21131 6276 21189 6304
rect 21131 6273 21143 6276
rect 21085 6267 21143 6273
rect 21177 6273 21189 6276
rect 21223 6273 21235 6307
rect 21177 6267 21235 6273
rect 5902 6196 5908 6248
rect 5960 6236 5966 6248
rect 13354 6236 13360 6248
rect 5960 6208 13360 6236
rect 5960 6196 5966 6208
rect 13354 6196 13360 6208
rect 13412 6196 13418 6248
rect 14458 6196 14464 6248
rect 14516 6236 14522 6248
rect 20640 6236 20668 6267
rect 30374 6264 30380 6316
rect 30432 6304 30438 6316
rect 31297 6307 31355 6313
rect 31297 6304 31309 6307
rect 30432 6276 31309 6304
rect 30432 6264 30438 6276
rect 31297 6273 31309 6276
rect 31343 6273 31355 6307
rect 31297 6267 31355 6273
rect 31478 6264 31484 6316
rect 31536 6304 31542 6316
rect 31665 6307 31723 6313
rect 31665 6304 31677 6307
rect 31536 6276 31677 6304
rect 31536 6264 31542 6276
rect 31665 6273 31677 6276
rect 31711 6273 31723 6307
rect 31665 6267 31723 6273
rect 22830 6236 22836 6248
rect 14516 6208 20576 6236
rect 20640 6208 22836 6236
rect 14516 6196 14522 6208
rect 18782 6128 18788 6180
rect 18840 6168 18846 6180
rect 20441 6171 20499 6177
rect 20441 6168 20453 6171
rect 18840 6140 20453 6168
rect 18840 6128 18846 6140
rect 20441 6137 20453 6140
rect 20487 6137 20499 6171
rect 20548 6168 20576 6208
rect 22830 6196 22836 6208
rect 22888 6196 22894 6248
rect 25130 6168 25136 6180
rect 20548 6140 25136 6168
rect 20441 6131 20499 6137
rect 25130 6128 25136 6140
rect 25188 6128 25194 6180
rect 26896 6140 31754 6168
rect 7377 6103 7435 6109
rect 7377 6069 7389 6103
rect 7423 6100 7435 6103
rect 9582 6100 9588 6112
rect 7423 6072 9588 6100
rect 7423 6069 7435 6072
rect 7377 6063 7435 6069
rect 9582 6060 9588 6072
rect 9640 6060 9646 6112
rect 9953 6103 10011 6109
rect 9953 6069 9965 6103
rect 9999 6100 10011 6103
rect 17770 6100 17776 6112
rect 9999 6072 17776 6100
rect 9999 6069 10011 6072
rect 9953 6063 10011 6069
rect 17770 6060 17776 6072
rect 17828 6060 17834 6112
rect 20898 6060 20904 6112
rect 20956 6100 20962 6112
rect 20993 6103 21051 6109
rect 20993 6100 21005 6103
rect 20956 6072 21005 6100
rect 20956 6060 20962 6072
rect 20993 6069 21005 6072
rect 21039 6069 21051 6103
rect 20993 6063 21051 6069
rect 21361 6103 21419 6109
rect 21361 6069 21373 6103
rect 21407 6100 21419 6103
rect 26896 6100 26924 6140
rect 21407 6072 26924 6100
rect 21407 6069 21419 6072
rect 21361 6063 21419 6069
rect 31478 6060 31484 6112
rect 31536 6060 31542 6112
rect 31726 6100 31754 6140
rect 31846 6100 31852 6112
rect 31726 6072 31852 6100
rect 31846 6060 31852 6072
rect 31904 6060 31910 6112
rect 1104 6010 32568 6032
rect 1104 5958 1950 6010
rect 2002 5958 2014 6010
rect 2066 5958 2078 6010
rect 2130 5958 2142 6010
rect 2194 5958 2206 6010
rect 2258 5958 7950 6010
rect 8002 5958 8014 6010
rect 8066 5958 8078 6010
rect 8130 5958 8142 6010
rect 8194 5958 8206 6010
rect 8258 5958 13950 6010
rect 14002 5958 14014 6010
rect 14066 5958 14078 6010
rect 14130 5958 14142 6010
rect 14194 5958 14206 6010
rect 14258 5958 19950 6010
rect 20002 5958 20014 6010
rect 20066 5958 20078 6010
rect 20130 5958 20142 6010
rect 20194 5958 20206 6010
rect 20258 5958 25950 6010
rect 26002 5958 26014 6010
rect 26066 5958 26078 6010
rect 26130 5958 26142 6010
rect 26194 5958 26206 6010
rect 26258 5958 31950 6010
rect 32002 5958 32014 6010
rect 32066 5958 32078 6010
rect 32130 5958 32142 6010
rect 32194 5958 32206 6010
rect 32258 5958 32568 6010
rect 1104 5936 32568 5958
rect 12066 5856 12072 5908
rect 12124 5896 12130 5908
rect 31202 5896 31208 5908
rect 12124 5868 31208 5896
rect 12124 5856 12130 5868
rect 31202 5856 31208 5868
rect 31260 5856 31266 5908
rect 15378 5788 15384 5840
rect 15436 5828 15442 5840
rect 29181 5831 29239 5837
rect 15436 5800 28396 5828
rect 15436 5788 15442 5800
rect 13078 5720 13084 5772
rect 13136 5760 13142 5772
rect 28368 5760 28396 5800
rect 29181 5797 29193 5831
rect 29227 5828 29239 5831
rect 30466 5828 30472 5840
rect 29227 5800 30472 5828
rect 29227 5797 29239 5800
rect 29181 5791 29239 5797
rect 30466 5788 30472 5800
rect 30524 5788 30530 5840
rect 31389 5831 31447 5837
rect 31389 5797 31401 5831
rect 31435 5828 31447 5831
rect 32030 5828 32036 5840
rect 31435 5800 32036 5828
rect 31435 5797 31447 5800
rect 31389 5791 31447 5797
rect 32030 5788 32036 5800
rect 32088 5788 32094 5840
rect 32122 5788 32128 5840
rect 32180 5788 32186 5840
rect 13136 5732 26464 5760
rect 28368 5732 31984 5760
rect 13136 5720 13142 5732
rect 3789 5695 3847 5701
rect 3789 5661 3801 5695
rect 3835 5692 3847 5695
rect 5534 5692 5540 5704
rect 3835 5664 5540 5692
rect 3835 5661 3847 5664
rect 3789 5655 3847 5661
rect 5534 5652 5540 5664
rect 5592 5652 5598 5704
rect 8846 5652 8852 5704
rect 8904 5692 8910 5704
rect 10965 5695 11023 5701
rect 10965 5692 10977 5695
rect 8904 5664 10977 5692
rect 8904 5652 8910 5664
rect 10965 5661 10977 5664
rect 11011 5661 11023 5695
rect 10965 5655 11023 5661
rect 18141 5695 18199 5701
rect 18141 5661 18153 5695
rect 18187 5692 18199 5695
rect 18233 5695 18291 5701
rect 18233 5692 18245 5695
rect 18187 5664 18245 5692
rect 18187 5661 18199 5664
rect 18141 5655 18199 5661
rect 18233 5661 18245 5664
rect 18279 5661 18291 5695
rect 18233 5655 18291 5661
rect 21177 5695 21235 5701
rect 21177 5661 21189 5695
rect 21223 5661 21235 5695
rect 21177 5655 21235 5661
rect 22097 5695 22155 5701
rect 22097 5661 22109 5695
rect 22143 5692 22155 5695
rect 22143 5664 26188 5692
rect 22143 5661 22155 5664
rect 22097 5655 22155 5661
rect 16758 5624 16764 5636
rect 6886 5596 16764 5624
rect 3973 5559 4031 5565
rect 3973 5525 3985 5559
rect 4019 5556 4031 5559
rect 6886 5556 6914 5596
rect 16758 5584 16764 5596
rect 16816 5584 16822 5636
rect 20530 5584 20536 5636
rect 20588 5624 20594 5636
rect 21192 5624 21220 5655
rect 20588 5596 21128 5624
rect 21192 5596 22094 5624
rect 20588 5584 20594 5596
rect 4019 5528 6914 5556
rect 4019 5525 4031 5528
rect 3973 5519 4031 5525
rect 7374 5516 7380 5568
rect 7432 5556 7438 5568
rect 8386 5556 8392 5568
rect 7432 5528 8392 5556
rect 7432 5516 7438 5528
rect 8386 5516 8392 5528
rect 8444 5516 8450 5568
rect 11149 5559 11207 5565
rect 11149 5525 11161 5559
rect 11195 5556 11207 5559
rect 17954 5556 17960 5568
rect 11195 5528 17960 5556
rect 11195 5525 11207 5528
rect 11149 5519 11207 5525
rect 17954 5516 17960 5528
rect 18012 5516 18018 5568
rect 18046 5516 18052 5568
rect 18104 5516 18110 5568
rect 18417 5559 18475 5565
rect 18417 5525 18429 5559
rect 18463 5556 18475 5559
rect 19794 5556 19800 5568
rect 18463 5528 19800 5556
rect 18463 5525 18475 5528
rect 18417 5519 18475 5525
rect 19794 5516 19800 5528
rect 19852 5516 19858 5568
rect 20346 5516 20352 5568
rect 20404 5556 20410 5568
rect 20993 5559 21051 5565
rect 20993 5556 21005 5559
rect 20404 5528 21005 5556
rect 20404 5516 20410 5528
rect 20993 5525 21005 5528
rect 21039 5525 21051 5559
rect 21100 5556 21128 5596
rect 21913 5559 21971 5565
rect 21913 5556 21925 5559
rect 21100 5528 21925 5556
rect 20993 5519 21051 5525
rect 21913 5525 21925 5528
rect 21959 5525 21971 5559
rect 22066 5556 22094 5596
rect 26050 5556 26056 5568
rect 22066 5528 26056 5556
rect 21913 5519 21971 5525
rect 26050 5516 26056 5528
rect 26108 5516 26114 5568
rect 26160 5556 26188 5664
rect 26436 5624 26464 5732
rect 28997 5695 29055 5701
rect 28997 5661 29009 5695
rect 29043 5692 29055 5695
rect 29270 5692 29276 5704
rect 29043 5664 29276 5692
rect 29043 5661 29055 5664
rect 28997 5655 29055 5661
rect 29270 5652 29276 5664
rect 29328 5652 29334 5704
rect 29546 5652 29552 5704
rect 29604 5692 29610 5704
rect 30653 5695 30711 5701
rect 30653 5692 30665 5695
rect 29604 5664 30665 5692
rect 29604 5652 29610 5664
rect 30653 5661 30665 5664
rect 30699 5661 30711 5695
rect 30653 5655 30711 5661
rect 31202 5652 31208 5704
rect 31260 5652 31266 5704
rect 31956 5701 31984 5732
rect 31573 5695 31631 5701
rect 31573 5661 31585 5695
rect 31619 5661 31631 5695
rect 31573 5655 31631 5661
rect 31941 5695 31999 5701
rect 31941 5661 31953 5695
rect 31987 5661 31999 5695
rect 31941 5655 31999 5661
rect 31588 5624 31616 5655
rect 26436 5596 31616 5624
rect 26786 5556 26792 5568
rect 26160 5528 26792 5556
rect 26786 5516 26792 5528
rect 26844 5516 26850 5568
rect 30837 5559 30895 5565
rect 30837 5525 30849 5559
rect 30883 5556 30895 5559
rect 31662 5556 31668 5568
rect 30883 5528 31668 5556
rect 30883 5525 30895 5528
rect 30837 5519 30895 5525
rect 31662 5516 31668 5528
rect 31720 5516 31726 5568
rect 31754 5516 31760 5568
rect 31812 5516 31818 5568
rect 1104 5466 32568 5488
rect 1104 5414 3010 5466
rect 3062 5414 3074 5466
rect 3126 5414 3138 5466
rect 3190 5414 3202 5466
rect 3254 5414 3266 5466
rect 3318 5414 9010 5466
rect 9062 5414 9074 5466
rect 9126 5414 9138 5466
rect 9190 5414 9202 5466
rect 9254 5414 9266 5466
rect 9318 5414 15010 5466
rect 15062 5414 15074 5466
rect 15126 5414 15138 5466
rect 15190 5414 15202 5466
rect 15254 5414 15266 5466
rect 15318 5414 21010 5466
rect 21062 5414 21074 5466
rect 21126 5414 21138 5466
rect 21190 5414 21202 5466
rect 21254 5414 21266 5466
rect 21318 5414 27010 5466
rect 27062 5414 27074 5466
rect 27126 5414 27138 5466
rect 27190 5414 27202 5466
rect 27254 5414 27266 5466
rect 27318 5414 32568 5466
rect 1104 5392 32568 5414
rect 12526 5312 12532 5364
rect 12584 5352 12590 5364
rect 18046 5352 18052 5364
rect 12584 5324 18052 5352
rect 12584 5312 12590 5324
rect 18046 5312 18052 5324
rect 18104 5312 18110 5364
rect 23382 5312 23388 5364
rect 23440 5352 23446 5364
rect 23661 5355 23719 5361
rect 23661 5352 23673 5355
rect 23440 5324 23673 5352
rect 23440 5312 23446 5324
rect 23661 5321 23673 5324
rect 23707 5321 23719 5355
rect 23661 5315 23719 5321
rect 27157 5355 27215 5361
rect 27157 5321 27169 5355
rect 27203 5352 27215 5355
rect 28994 5352 29000 5364
rect 27203 5324 29000 5352
rect 27203 5321 27215 5324
rect 27157 5315 27215 5321
rect 28994 5312 29000 5324
rect 29052 5312 29058 5364
rect 19426 5244 19432 5296
rect 19484 5284 19490 5296
rect 19484 5256 31708 5284
rect 19484 5244 19490 5256
rect 4154 5176 4160 5228
rect 4212 5216 4218 5228
rect 5445 5219 5503 5225
rect 5445 5216 5457 5219
rect 4212 5188 5457 5216
rect 4212 5176 4218 5188
rect 5445 5185 5457 5188
rect 5491 5185 5503 5219
rect 10597 5219 10655 5225
rect 10597 5216 10609 5219
rect 5445 5179 5503 5185
rect 6886 5188 10609 5216
rect 4982 5108 4988 5160
rect 5040 5148 5046 5160
rect 6886 5148 6914 5188
rect 10597 5185 10609 5188
rect 10643 5185 10655 5219
rect 10597 5179 10655 5185
rect 23201 5219 23259 5225
rect 23201 5185 23213 5219
rect 23247 5216 23259 5219
rect 23293 5219 23351 5225
rect 23293 5216 23305 5219
rect 23247 5188 23305 5216
rect 23247 5185 23259 5188
rect 23201 5179 23259 5185
rect 23293 5185 23305 5188
rect 23339 5185 23351 5219
rect 23293 5179 23351 5185
rect 23845 5219 23903 5225
rect 23845 5185 23857 5219
rect 23891 5216 23903 5219
rect 26510 5216 26516 5228
rect 23891 5188 26516 5216
rect 23891 5185 23903 5188
rect 23845 5179 23903 5185
rect 26510 5176 26516 5188
rect 26568 5176 26574 5228
rect 26973 5219 27031 5225
rect 26973 5185 26985 5219
rect 27019 5216 27031 5219
rect 29086 5216 29092 5228
rect 27019 5188 29092 5216
rect 27019 5185 27031 5188
rect 26973 5179 27031 5185
rect 29086 5176 29092 5188
rect 29144 5176 29150 5228
rect 31680 5225 31708 5256
rect 31297 5219 31355 5225
rect 31297 5185 31309 5219
rect 31343 5185 31355 5219
rect 31297 5179 31355 5185
rect 31665 5219 31723 5225
rect 31665 5185 31677 5219
rect 31711 5185 31723 5219
rect 31665 5179 31723 5185
rect 5040 5120 6914 5148
rect 5040 5108 5046 5120
rect 26234 5108 26240 5160
rect 26292 5148 26298 5160
rect 27338 5148 27344 5160
rect 26292 5120 27344 5148
rect 26292 5108 26298 5120
rect 27338 5108 27344 5120
rect 27396 5108 27402 5160
rect 27614 5108 27620 5160
rect 27672 5148 27678 5160
rect 31312 5148 31340 5179
rect 27672 5120 31340 5148
rect 27672 5108 27678 5120
rect 5629 5015 5687 5021
rect 5629 4981 5641 5015
rect 5675 5012 5687 5015
rect 9490 5012 9496 5024
rect 5675 4984 9496 5012
rect 5675 4981 5687 4984
rect 5629 4975 5687 4981
rect 9490 4972 9496 4984
rect 9548 4972 9554 5024
rect 10781 5015 10839 5021
rect 10781 4981 10793 5015
rect 10827 5012 10839 5015
rect 13630 5012 13636 5024
rect 10827 4984 13636 5012
rect 10827 4981 10839 4984
rect 10781 4975 10839 4981
rect 13630 4972 13636 4984
rect 13688 4972 13694 5024
rect 15470 4972 15476 5024
rect 15528 5012 15534 5024
rect 19426 5012 19432 5024
rect 15528 4984 19432 5012
rect 15528 4972 15534 4984
rect 19426 4972 19432 4984
rect 19484 4972 19490 5024
rect 23014 4972 23020 5024
rect 23072 5012 23078 5024
rect 23109 5015 23167 5021
rect 23109 5012 23121 5015
rect 23072 4984 23121 5012
rect 23072 4972 23078 4984
rect 23109 4981 23121 4984
rect 23155 4981 23167 5015
rect 23109 4975 23167 4981
rect 23474 4972 23480 5024
rect 23532 4972 23538 5024
rect 31478 4972 31484 5024
rect 31536 4972 31542 5024
rect 31849 5015 31907 5021
rect 31849 4981 31861 5015
rect 31895 5012 31907 5015
rect 32858 5012 32864 5024
rect 31895 4984 32864 5012
rect 31895 4981 31907 4984
rect 31849 4975 31907 4981
rect 32858 4972 32864 4984
rect 32916 4972 32922 5024
rect 1104 4922 32568 4944
rect 1104 4870 1950 4922
rect 2002 4870 2014 4922
rect 2066 4870 2078 4922
rect 2130 4870 2142 4922
rect 2194 4870 2206 4922
rect 2258 4870 7950 4922
rect 8002 4870 8014 4922
rect 8066 4870 8078 4922
rect 8130 4870 8142 4922
rect 8194 4870 8206 4922
rect 8258 4870 13950 4922
rect 14002 4870 14014 4922
rect 14066 4870 14078 4922
rect 14130 4870 14142 4922
rect 14194 4870 14206 4922
rect 14258 4870 19950 4922
rect 20002 4870 20014 4922
rect 20066 4870 20078 4922
rect 20130 4870 20142 4922
rect 20194 4870 20206 4922
rect 20258 4870 25950 4922
rect 26002 4870 26014 4922
rect 26066 4870 26078 4922
rect 26130 4870 26142 4922
rect 26194 4870 26206 4922
rect 26258 4870 31950 4922
rect 32002 4870 32014 4922
rect 32066 4870 32078 4922
rect 32130 4870 32142 4922
rect 32194 4870 32206 4922
rect 32258 4870 32568 4922
rect 1104 4848 32568 4870
rect 12529 4811 12587 4817
rect 12529 4777 12541 4811
rect 12575 4808 12587 4811
rect 14918 4808 14924 4820
rect 12575 4780 14924 4808
rect 12575 4777 12587 4780
rect 12529 4771 12587 4777
rect 14918 4768 14924 4780
rect 14976 4768 14982 4820
rect 25038 4768 25044 4820
rect 25096 4768 25102 4820
rect 11701 4743 11759 4749
rect 11701 4709 11713 4743
rect 11747 4740 11759 4743
rect 12802 4740 12808 4752
rect 11747 4712 12808 4740
rect 11747 4709 11759 4712
rect 11701 4703 11759 4709
rect 12802 4700 12808 4712
rect 12860 4700 12866 4752
rect 12989 4743 13047 4749
rect 12989 4709 13001 4743
rect 13035 4740 13047 4743
rect 15378 4740 15384 4752
rect 13035 4712 15384 4740
rect 13035 4709 13047 4712
rect 12989 4703 13047 4709
rect 15378 4700 15384 4712
rect 15436 4700 15442 4752
rect 11882 4632 11888 4684
rect 11940 4672 11946 4684
rect 11940 4644 14228 4672
rect 11940 4632 11946 4644
rect 2593 4607 2651 4613
rect 2593 4573 2605 4607
rect 2639 4604 2651 4607
rect 5258 4604 5264 4616
rect 2639 4576 5264 4604
rect 2639 4573 2651 4576
rect 2593 4567 2651 4573
rect 5258 4564 5264 4576
rect 5316 4564 5322 4616
rect 6638 4564 6644 4616
rect 6696 4604 6702 4616
rect 14200 4613 14228 4644
rect 23474 4632 23480 4684
rect 23532 4672 23538 4684
rect 23532 4644 31616 4672
rect 23532 4632 23538 4644
rect 31588 4613 31616 4644
rect 11517 4607 11575 4613
rect 11517 4604 11529 4607
rect 6696 4576 11529 4604
rect 6696 4564 6702 4576
rect 11517 4573 11529 4576
rect 11563 4573 11575 4607
rect 11517 4567 11575 4573
rect 12345 4607 12403 4613
rect 12345 4573 12357 4607
rect 12391 4573 12403 4607
rect 12805 4607 12863 4613
rect 12805 4604 12817 4607
rect 12345 4567 12403 4573
rect 12452 4576 12817 4604
rect 6914 4496 6920 4548
rect 6972 4536 6978 4548
rect 12360 4536 12388 4567
rect 6972 4508 12388 4536
rect 6972 4496 6978 4508
rect 2777 4471 2835 4477
rect 2777 4437 2789 4471
rect 2823 4468 2835 4471
rect 7098 4468 7104 4480
rect 2823 4440 7104 4468
rect 2823 4437 2835 4440
rect 2777 4431 2835 4437
rect 7098 4428 7104 4440
rect 7156 4428 7162 4480
rect 7190 4428 7196 4480
rect 7248 4468 7254 4480
rect 12452 4468 12480 4576
rect 12805 4573 12817 4576
rect 12851 4573 12863 4607
rect 12805 4567 12863 4573
rect 14185 4607 14243 4613
rect 14185 4573 14197 4607
rect 14231 4573 14243 4607
rect 24857 4607 24915 4613
rect 14185 4567 14243 4573
rect 14292 4576 16574 4604
rect 7248 4440 12480 4468
rect 7248 4428 7254 4440
rect 13078 4428 13084 4480
rect 13136 4468 13142 4480
rect 14292 4468 14320 4576
rect 16546 4536 16574 4576
rect 24857 4573 24869 4607
rect 24903 4604 24915 4607
rect 25225 4607 25283 4613
rect 24903 4576 25176 4604
rect 24903 4573 24915 4576
rect 24857 4567 24915 4573
rect 25148 4536 25176 4576
rect 25225 4573 25237 4607
rect 25271 4604 25283 4607
rect 25317 4607 25375 4613
rect 25317 4604 25329 4607
rect 25271 4576 25329 4604
rect 25271 4573 25283 4576
rect 25225 4567 25283 4573
rect 25317 4573 25329 4576
rect 25363 4573 25375 4607
rect 25317 4567 25375 4573
rect 31573 4607 31631 4613
rect 31573 4573 31585 4607
rect 31619 4573 31631 4607
rect 31573 4567 31631 4573
rect 31846 4564 31852 4616
rect 31904 4604 31910 4616
rect 31941 4607 31999 4613
rect 31941 4604 31953 4607
rect 31904 4576 31953 4604
rect 31904 4564 31910 4576
rect 31941 4573 31953 4576
rect 31987 4573 31999 4607
rect 31941 4567 31999 4573
rect 28718 4536 28724 4548
rect 16546 4508 22094 4536
rect 25148 4508 28724 4536
rect 13136 4440 14320 4468
rect 14369 4471 14427 4477
rect 13136 4428 13142 4440
rect 14369 4437 14381 4471
rect 14415 4468 14427 4471
rect 20346 4468 20352 4480
rect 14415 4440 20352 4468
rect 14415 4437 14427 4440
rect 14369 4431 14427 4437
rect 20346 4428 20352 4440
rect 20404 4428 20410 4480
rect 22066 4468 22094 4508
rect 28718 4496 28724 4508
rect 28776 4496 28782 4548
rect 25133 4471 25191 4477
rect 25133 4468 25145 4471
rect 22066 4440 25145 4468
rect 25133 4437 25145 4440
rect 25179 4437 25191 4471
rect 25133 4431 25191 4437
rect 25501 4471 25559 4477
rect 25501 4437 25513 4471
rect 25547 4468 25559 4471
rect 31294 4468 31300 4480
rect 25547 4440 31300 4468
rect 25547 4437 25559 4440
rect 25501 4431 25559 4437
rect 31294 4428 31300 4440
rect 31352 4428 31358 4480
rect 31754 4428 31760 4480
rect 31812 4428 31818 4480
rect 32122 4428 32128 4480
rect 32180 4428 32186 4480
rect 1104 4378 32568 4400
rect 1104 4326 3010 4378
rect 3062 4326 3074 4378
rect 3126 4326 3138 4378
rect 3190 4326 3202 4378
rect 3254 4326 3266 4378
rect 3318 4326 9010 4378
rect 9062 4326 9074 4378
rect 9126 4326 9138 4378
rect 9190 4326 9202 4378
rect 9254 4326 9266 4378
rect 9318 4326 15010 4378
rect 15062 4326 15074 4378
rect 15126 4326 15138 4378
rect 15190 4326 15202 4378
rect 15254 4326 15266 4378
rect 15318 4326 21010 4378
rect 21062 4326 21074 4378
rect 21126 4326 21138 4378
rect 21190 4326 21202 4378
rect 21254 4326 21266 4378
rect 21318 4326 27010 4378
rect 27062 4326 27074 4378
rect 27126 4326 27138 4378
rect 27190 4326 27202 4378
rect 27254 4326 27266 4378
rect 27318 4326 32568 4378
rect 1104 4304 32568 4326
rect 7098 4224 7104 4276
rect 7156 4264 7162 4276
rect 10134 4264 10140 4276
rect 7156 4236 10140 4264
rect 7156 4224 7162 4236
rect 10134 4224 10140 4236
rect 10192 4224 10198 4276
rect 13265 4267 13323 4273
rect 13265 4233 13277 4267
rect 13311 4233 13323 4267
rect 13265 4227 13323 4233
rect 18233 4267 18291 4273
rect 18233 4233 18245 4267
rect 18279 4264 18291 4267
rect 18279 4236 19840 4264
rect 18279 4233 18291 4236
rect 18233 4227 18291 4233
rect 12161 4131 12219 4137
rect 12161 4097 12173 4131
rect 12207 4097 12219 4131
rect 12161 4091 12219 4097
rect 12176 4060 12204 4091
rect 12434 4088 12440 4140
rect 12492 4088 12498 4140
rect 12713 4131 12771 4137
rect 12713 4097 12725 4131
rect 12759 4128 12771 4131
rect 12986 4128 12992 4140
rect 12759 4100 12992 4128
rect 12759 4097 12771 4100
rect 12713 4091 12771 4097
rect 12986 4088 12992 4100
rect 13044 4088 13050 4140
rect 13081 4131 13139 4137
rect 13081 4097 13093 4131
rect 13127 4097 13139 4131
rect 13081 4091 13139 4097
rect 12894 4060 12900 4072
rect 12176 4032 12900 4060
rect 12894 4020 12900 4032
rect 12952 4020 12958 4072
rect 12710 3952 12716 4004
rect 12768 3992 12774 4004
rect 13096 3992 13124 4091
rect 13280 4060 13308 4227
rect 13832 4168 14596 4196
rect 13538 4088 13544 4140
rect 13596 4088 13602 4140
rect 13832 4137 13860 4168
rect 14568 4140 14596 4168
rect 19352 4168 19656 4196
rect 13817 4131 13875 4137
rect 13817 4097 13829 4131
rect 13863 4097 13875 4131
rect 13817 4091 13875 4097
rect 13906 4088 13912 4140
rect 13964 4128 13970 4140
rect 14185 4131 14243 4137
rect 14185 4128 14197 4131
rect 13964 4100 14197 4128
rect 13964 4088 13970 4100
rect 14185 4097 14197 4100
rect 14231 4097 14243 4131
rect 14185 4091 14243 4097
rect 14458 4088 14464 4140
rect 14516 4088 14522 4140
rect 14550 4088 14556 4140
rect 14608 4088 14614 4140
rect 14826 4088 14832 4140
rect 14884 4128 14890 4140
rect 15105 4131 15163 4137
rect 15105 4128 15117 4131
rect 14884 4100 15117 4128
rect 14884 4088 14890 4100
rect 15105 4097 15117 4100
rect 15151 4097 15163 4131
rect 15105 4091 15163 4097
rect 15194 4088 15200 4140
rect 15252 4128 15258 4140
rect 15749 4131 15807 4137
rect 15749 4128 15761 4131
rect 15252 4100 15761 4128
rect 15252 4088 15258 4100
rect 15749 4097 15761 4100
rect 15795 4097 15807 4131
rect 15749 4091 15807 4097
rect 16666 4088 16672 4140
rect 16724 4088 16730 4140
rect 17126 4088 17132 4140
rect 17184 4088 17190 4140
rect 17497 4131 17555 4137
rect 17497 4097 17509 4131
rect 17543 4128 17555 4131
rect 17589 4131 17647 4137
rect 17589 4128 17601 4131
rect 17543 4100 17601 4128
rect 17543 4097 17555 4100
rect 17497 4091 17555 4097
rect 17589 4097 17601 4100
rect 17635 4097 17647 4131
rect 17589 4091 17647 4097
rect 18046 4088 18052 4140
rect 18104 4088 18110 4140
rect 19061 4131 19119 4137
rect 19061 4097 19073 4131
rect 19107 4128 19119 4131
rect 19352 4128 19380 4168
rect 19107 4100 19380 4128
rect 19429 4131 19487 4137
rect 19107 4097 19119 4100
rect 19061 4091 19119 4097
rect 19429 4097 19441 4131
rect 19475 4097 19487 4131
rect 19628 4128 19656 4168
rect 19705 4131 19763 4137
rect 19705 4128 19717 4131
rect 19628 4100 19717 4128
rect 19429 4091 19487 4097
rect 19705 4097 19717 4100
rect 19751 4097 19763 4131
rect 19812 4128 19840 4236
rect 22002 4128 22008 4140
rect 19812 4100 22008 4128
rect 19705 4091 19763 4097
rect 13280 4032 18828 4060
rect 18506 3992 18512 4004
rect 12768 3964 13124 3992
rect 13188 3964 18512 3992
rect 12768 3952 12774 3964
rect 12342 3884 12348 3936
rect 12400 3884 12406 3936
rect 12618 3884 12624 3936
rect 12676 3884 12682 3936
rect 12897 3927 12955 3933
rect 12897 3893 12909 3927
rect 12943 3924 12955 3927
rect 13188 3924 13216 3964
rect 18506 3952 18512 3964
rect 18564 3952 18570 4004
rect 12943 3896 13216 3924
rect 12943 3893 12955 3896
rect 12897 3887 12955 3893
rect 13722 3884 13728 3936
rect 13780 3884 13786 3936
rect 14001 3927 14059 3933
rect 14001 3893 14013 3927
rect 14047 3924 14059 3927
rect 14274 3924 14280 3936
rect 14047 3896 14280 3924
rect 14047 3893 14059 3896
rect 14001 3887 14059 3893
rect 14274 3884 14280 3896
rect 14332 3884 14338 3936
rect 14366 3884 14372 3936
rect 14424 3884 14430 3936
rect 14642 3884 14648 3936
rect 14700 3884 14706 3936
rect 15286 3884 15292 3936
rect 15344 3884 15350 3936
rect 15930 3884 15936 3936
rect 15988 3884 15994 3936
rect 16850 3884 16856 3936
rect 16908 3884 16914 3936
rect 17310 3884 17316 3936
rect 17368 3884 17374 3936
rect 17402 3884 17408 3936
rect 17460 3884 17466 3936
rect 17773 3927 17831 3933
rect 17773 3893 17785 3927
rect 17819 3924 17831 3927
rect 18690 3924 18696 3936
rect 17819 3896 18696 3924
rect 17819 3893 17831 3896
rect 17773 3887 17831 3893
rect 18690 3884 18696 3896
rect 18748 3884 18754 3936
rect 18800 3924 18828 4032
rect 18966 4020 18972 4072
rect 19024 4020 19030 4072
rect 19444 4060 19472 4091
rect 22002 4088 22008 4100
rect 22060 4088 22066 4140
rect 22370 4088 22376 4140
rect 22428 4088 22434 4140
rect 23290 4088 23296 4140
rect 23348 4088 23354 4140
rect 23477 4131 23535 4137
rect 23477 4097 23489 4131
rect 23523 4097 23535 4131
rect 23477 4091 23535 4097
rect 23845 4131 23903 4137
rect 23845 4097 23857 4131
rect 23891 4128 23903 4131
rect 28442 4128 28448 4140
rect 23891 4100 28448 4128
rect 23891 4097 23903 4100
rect 23845 4091 23903 4097
rect 19352 4032 19472 4060
rect 23492 4060 23520 4091
rect 28442 4088 28448 4100
rect 28500 4088 28506 4140
rect 31294 4088 31300 4140
rect 31352 4088 31358 4140
rect 31665 4131 31723 4137
rect 31665 4097 31677 4131
rect 31711 4097 31723 4131
rect 31665 4091 31723 4097
rect 28166 4060 28172 4072
rect 23492 4032 28172 4060
rect 18874 3952 18880 4004
rect 18932 3992 18938 4004
rect 19352 4001 19380 4032
rect 28166 4020 28172 4032
rect 28224 4020 28230 4072
rect 28994 4020 29000 4072
rect 29052 4060 29058 4072
rect 31680 4060 31708 4091
rect 29052 4032 31708 4060
rect 29052 4020 29058 4032
rect 19337 3995 19395 4001
rect 19337 3992 19349 3995
rect 18932 3964 19349 3992
rect 18932 3952 18938 3964
rect 19337 3961 19349 3964
rect 19383 3961 19395 3995
rect 20898 3992 20904 4004
rect 19337 3955 19395 3961
rect 19536 3964 20904 3992
rect 19536 3924 19564 3964
rect 20898 3952 20904 3964
rect 20956 3952 20962 4004
rect 22186 3952 22192 4004
rect 22244 3952 22250 4004
rect 23106 3952 23112 4004
rect 23164 3952 23170 4004
rect 23658 3952 23664 4004
rect 23716 3952 23722 4004
rect 24029 3995 24087 4001
rect 24029 3961 24041 3995
rect 24075 3992 24087 3995
rect 26418 3992 26424 4004
rect 24075 3964 26424 3992
rect 24075 3961 24087 3964
rect 24029 3955 24087 3961
rect 26418 3952 26424 3964
rect 26476 3952 26482 4004
rect 18800 3896 19564 3924
rect 19613 3927 19671 3933
rect 19613 3893 19625 3927
rect 19659 3924 19671 3927
rect 19794 3924 19800 3936
rect 19659 3896 19800 3924
rect 19659 3893 19671 3896
rect 19613 3887 19671 3893
rect 19794 3884 19800 3896
rect 19852 3884 19858 3936
rect 19889 3927 19947 3933
rect 19889 3893 19901 3927
rect 19935 3924 19947 3927
rect 31294 3924 31300 3936
rect 19935 3896 31300 3924
rect 19935 3893 19947 3896
rect 19889 3887 19947 3893
rect 31294 3884 31300 3896
rect 31352 3884 31358 3936
rect 31478 3884 31484 3936
rect 31536 3884 31542 3936
rect 31849 3927 31907 3933
rect 31849 3893 31861 3927
rect 31895 3924 31907 3927
rect 32858 3924 32864 3936
rect 31895 3896 32864 3924
rect 31895 3893 31907 3896
rect 31849 3887 31907 3893
rect 32858 3884 32864 3896
rect 32916 3884 32922 3936
rect 1104 3834 32568 3856
rect 1104 3782 1950 3834
rect 2002 3782 2014 3834
rect 2066 3782 2078 3834
rect 2130 3782 2142 3834
rect 2194 3782 2206 3834
rect 2258 3782 7950 3834
rect 8002 3782 8014 3834
rect 8066 3782 8078 3834
rect 8130 3782 8142 3834
rect 8194 3782 8206 3834
rect 8258 3782 13950 3834
rect 14002 3782 14014 3834
rect 14066 3782 14078 3834
rect 14130 3782 14142 3834
rect 14194 3782 14206 3834
rect 14258 3782 19950 3834
rect 20002 3782 20014 3834
rect 20066 3782 20078 3834
rect 20130 3782 20142 3834
rect 20194 3782 20206 3834
rect 20258 3782 25950 3834
rect 26002 3782 26014 3834
rect 26066 3782 26078 3834
rect 26130 3782 26142 3834
rect 26194 3782 26206 3834
rect 26258 3782 31950 3834
rect 32002 3782 32014 3834
rect 32066 3782 32078 3834
rect 32130 3782 32142 3834
rect 32194 3782 32206 3834
rect 32258 3782 32568 3834
rect 1104 3760 32568 3782
rect 9398 3680 9404 3732
rect 9456 3720 9462 3732
rect 13538 3720 13544 3732
rect 9456 3692 13544 3720
rect 9456 3680 9462 3692
rect 13538 3680 13544 3692
rect 13596 3680 13602 3732
rect 13722 3680 13728 3732
rect 13780 3720 13786 3732
rect 15470 3720 15476 3732
rect 13780 3692 15476 3720
rect 13780 3680 13786 3692
rect 15470 3680 15476 3692
rect 15528 3680 15534 3732
rect 15930 3680 15936 3732
rect 15988 3720 15994 3732
rect 17218 3720 17224 3732
rect 15988 3692 17224 3720
rect 15988 3680 15994 3692
rect 17218 3680 17224 3692
rect 17276 3680 17282 3732
rect 17310 3680 17316 3732
rect 17368 3720 17374 3732
rect 22738 3720 22744 3732
rect 17368 3692 22744 3720
rect 17368 3680 17374 3692
rect 22738 3680 22744 3692
rect 22796 3680 22802 3732
rect 23290 3680 23296 3732
rect 23348 3720 23354 3732
rect 27890 3720 27896 3732
rect 23348 3692 27896 3720
rect 23348 3680 23354 3692
rect 27890 3680 27896 3692
rect 27948 3680 27954 3732
rect 12618 3612 12624 3664
rect 12676 3652 12682 3664
rect 19886 3652 19892 3664
rect 12676 3624 19892 3652
rect 12676 3612 12682 3624
rect 19886 3612 19892 3624
rect 19944 3612 19950 3664
rect 21450 3652 21456 3664
rect 20088 3624 21456 3652
rect 12158 3544 12164 3596
rect 12216 3584 12222 3596
rect 13722 3584 13728 3596
rect 12216 3556 13728 3584
rect 12216 3544 12222 3556
rect 13722 3544 13728 3556
rect 13780 3544 13786 3596
rect 14274 3544 14280 3596
rect 14332 3584 14338 3596
rect 17494 3584 17500 3596
rect 14332 3556 17500 3584
rect 14332 3544 14338 3556
rect 17494 3544 17500 3556
rect 17552 3544 17558 3596
rect 20088 3584 20116 3624
rect 21450 3612 21456 3624
rect 21508 3612 21514 3664
rect 21913 3655 21971 3661
rect 21913 3621 21925 3655
rect 21959 3652 21971 3655
rect 24118 3652 24124 3664
rect 21959 3624 24124 3652
rect 21959 3621 21971 3624
rect 21913 3615 21971 3621
rect 24118 3612 24124 3624
rect 24176 3612 24182 3664
rect 25593 3655 25651 3661
rect 25593 3621 25605 3655
rect 25639 3652 25651 3655
rect 25639 3624 31984 3652
rect 25639 3621 25651 3624
rect 25593 3615 25651 3621
rect 22278 3584 22284 3596
rect 19260 3556 20116 3584
rect 20180 3556 22284 3584
rect 12437 3519 12495 3525
rect 12437 3485 12449 3519
rect 12483 3516 12495 3519
rect 13814 3516 13820 3528
rect 12483 3488 13820 3516
rect 12483 3485 12495 3488
rect 12437 3479 12495 3485
rect 13814 3476 13820 3488
rect 13872 3476 13878 3528
rect 14182 3476 14188 3528
rect 14240 3516 14246 3528
rect 15102 3516 15108 3528
rect 14240 3488 15108 3516
rect 14240 3476 14246 3488
rect 15102 3476 15108 3488
rect 15160 3476 15166 3528
rect 15286 3476 15292 3528
rect 15344 3516 15350 3528
rect 19260 3516 19288 3556
rect 15344 3488 19288 3516
rect 15344 3476 15350 3488
rect 19334 3476 19340 3528
rect 19392 3516 19398 3528
rect 19797 3519 19855 3525
rect 19797 3516 19809 3519
rect 19392 3488 19809 3516
rect 19392 3476 19398 3488
rect 19797 3485 19809 3488
rect 19843 3485 19855 3519
rect 19797 3479 19855 3485
rect 20073 3519 20131 3525
rect 20073 3485 20085 3519
rect 20119 3485 20131 3519
rect 20073 3479 20131 3485
rect 12526 3408 12532 3460
rect 12584 3448 12590 3460
rect 14458 3448 14464 3460
rect 12584 3420 14464 3448
rect 12584 3408 12590 3420
rect 14458 3408 14464 3420
rect 14516 3408 14522 3460
rect 14642 3408 14648 3460
rect 14700 3448 14706 3460
rect 17862 3448 17868 3460
rect 14700 3420 17868 3448
rect 14700 3408 14706 3420
rect 17862 3408 17868 3420
rect 17920 3408 17926 3460
rect 19518 3408 19524 3460
rect 19576 3448 19582 3460
rect 20088 3448 20116 3479
rect 19576 3420 20116 3448
rect 19576 3408 19582 3420
rect 12621 3383 12679 3389
rect 12621 3349 12633 3383
rect 12667 3380 12679 3383
rect 15930 3380 15936 3392
rect 12667 3352 15936 3380
rect 12667 3349 12679 3352
rect 12621 3343 12679 3349
rect 15930 3340 15936 3352
rect 15988 3340 15994 3392
rect 17218 3340 17224 3392
rect 17276 3380 17282 3392
rect 19150 3380 19156 3392
rect 17276 3352 19156 3380
rect 17276 3340 17282 3352
rect 19150 3340 19156 3352
rect 19208 3340 19214 3392
rect 19981 3383 20039 3389
rect 19981 3349 19993 3383
rect 20027 3380 20039 3383
rect 20180 3380 20208 3556
rect 22278 3544 22284 3556
rect 22336 3544 22342 3596
rect 22370 3544 22376 3596
rect 22428 3584 22434 3596
rect 27614 3584 27620 3596
rect 22428 3556 27620 3584
rect 22428 3544 22434 3556
rect 27614 3544 27620 3556
rect 27672 3544 27678 3596
rect 20533 3519 20591 3525
rect 20533 3485 20545 3519
rect 20579 3516 20591 3519
rect 20625 3519 20683 3525
rect 20625 3516 20637 3519
rect 20579 3488 20637 3516
rect 20579 3485 20591 3488
rect 20533 3479 20591 3485
rect 20625 3485 20637 3488
rect 20671 3485 20683 3519
rect 20625 3479 20683 3485
rect 20714 3476 20720 3528
rect 20772 3516 20778 3528
rect 21269 3519 21327 3525
rect 21269 3516 21281 3519
rect 20772 3488 21281 3516
rect 20772 3476 20778 3488
rect 21269 3485 21281 3488
rect 21315 3516 21327 3519
rect 21453 3519 21511 3525
rect 21453 3516 21465 3519
rect 21315 3488 21465 3516
rect 21315 3485 21327 3488
rect 21269 3479 21327 3485
rect 21453 3485 21465 3488
rect 21499 3485 21511 3519
rect 21453 3479 21511 3485
rect 21726 3476 21732 3528
rect 21784 3516 21790 3528
rect 31956 3525 31984 3624
rect 22005 3519 22063 3525
rect 22005 3516 22017 3519
rect 21784 3488 22017 3516
rect 21784 3476 21790 3488
rect 22005 3485 22017 3488
rect 22051 3485 22063 3519
rect 22005 3479 22063 3485
rect 25317 3519 25375 3525
rect 25317 3485 25329 3519
rect 25363 3516 25375 3519
rect 25409 3519 25467 3525
rect 25409 3516 25421 3519
rect 25363 3488 25421 3516
rect 25363 3485 25375 3488
rect 25317 3479 25375 3485
rect 25409 3485 25421 3488
rect 25455 3485 25467 3519
rect 25409 3479 25467 3485
rect 25869 3519 25927 3525
rect 25869 3485 25881 3519
rect 25915 3516 25927 3519
rect 25961 3519 26019 3525
rect 25961 3516 25973 3519
rect 25915 3488 25973 3516
rect 25915 3485 25927 3488
rect 25869 3479 25927 3485
rect 25961 3485 25973 3488
rect 26007 3485 26019 3519
rect 25961 3479 26019 3485
rect 26329 3519 26387 3525
rect 26329 3485 26341 3519
rect 26375 3516 26387 3519
rect 26421 3519 26479 3525
rect 26421 3516 26433 3519
rect 26375 3488 26433 3516
rect 26375 3485 26387 3488
rect 26329 3479 26387 3485
rect 26421 3485 26433 3488
rect 26467 3485 26479 3519
rect 26421 3479 26479 3485
rect 31573 3519 31631 3525
rect 31573 3485 31585 3519
rect 31619 3485 31631 3519
rect 31573 3479 31631 3485
rect 31941 3519 31999 3525
rect 31941 3485 31953 3519
rect 31987 3485 31999 3519
rect 31941 3479 31999 3485
rect 20346 3408 20352 3460
rect 20404 3448 20410 3460
rect 21358 3448 21364 3460
rect 20404 3420 21364 3448
rect 20404 3408 20410 3420
rect 21358 3408 21364 3420
rect 21416 3408 21422 3460
rect 23934 3448 23940 3460
rect 21652 3420 23940 3448
rect 20027 3352 20208 3380
rect 20027 3349 20039 3352
rect 19981 3343 20039 3349
rect 20254 3340 20260 3392
rect 20312 3340 20318 3392
rect 20438 3340 20444 3392
rect 20496 3340 20502 3392
rect 20806 3340 20812 3392
rect 20864 3340 20870 3392
rect 21652 3389 21680 3420
rect 23934 3408 23940 3420
rect 23992 3408 23998 3460
rect 25222 3408 25228 3460
rect 25280 3408 25286 3460
rect 31588 3448 31616 3479
rect 26160 3420 31616 3448
rect 21637 3383 21695 3389
rect 21637 3349 21649 3383
rect 21683 3349 21695 3383
rect 21637 3343 21695 3349
rect 25774 3340 25780 3392
rect 25832 3340 25838 3392
rect 26160 3389 26188 3420
rect 26145 3383 26203 3389
rect 26145 3349 26157 3383
rect 26191 3349 26203 3383
rect 26145 3343 26203 3349
rect 26234 3340 26240 3392
rect 26292 3340 26298 3392
rect 26605 3383 26663 3389
rect 26605 3349 26617 3383
rect 26651 3380 26663 3383
rect 31662 3380 31668 3392
rect 26651 3352 31668 3380
rect 26651 3349 26663 3352
rect 26605 3343 26663 3349
rect 31662 3340 31668 3352
rect 31720 3340 31726 3392
rect 31754 3340 31760 3392
rect 31812 3340 31818 3392
rect 32122 3340 32128 3392
rect 32180 3340 32186 3392
rect 1104 3290 32568 3312
rect 1104 3238 3010 3290
rect 3062 3238 3074 3290
rect 3126 3238 3138 3290
rect 3190 3238 3202 3290
rect 3254 3238 3266 3290
rect 3318 3238 9010 3290
rect 9062 3238 9074 3290
rect 9126 3238 9138 3290
rect 9190 3238 9202 3290
rect 9254 3238 9266 3290
rect 9318 3238 15010 3290
rect 15062 3238 15074 3290
rect 15126 3238 15138 3290
rect 15190 3238 15202 3290
rect 15254 3238 15266 3290
rect 15318 3238 21010 3290
rect 21062 3238 21074 3290
rect 21126 3238 21138 3290
rect 21190 3238 21202 3290
rect 21254 3238 21266 3290
rect 21318 3238 27010 3290
rect 27062 3238 27074 3290
rect 27126 3238 27138 3290
rect 27190 3238 27202 3290
rect 27254 3238 27266 3290
rect 27318 3238 32568 3290
rect 1104 3216 32568 3238
rect 14366 3136 14372 3188
rect 14424 3176 14430 3188
rect 20622 3176 20628 3188
rect 14424 3148 20628 3176
rect 14424 3136 14430 3148
rect 20622 3136 20628 3148
rect 20680 3136 20686 3188
rect 20806 3136 20812 3188
rect 20864 3176 20870 3188
rect 30926 3176 30932 3188
rect 20864 3148 30932 3176
rect 20864 3136 20870 3148
rect 30926 3136 30932 3148
rect 30984 3136 30990 3188
rect 11606 3068 11612 3120
rect 11664 3108 11670 3120
rect 14826 3108 14832 3120
rect 11664 3080 14832 3108
rect 11664 3068 11670 3080
rect 14826 3068 14832 3080
rect 14884 3068 14890 3120
rect 18506 3068 18512 3120
rect 18564 3108 18570 3120
rect 18564 3080 19564 3108
rect 18564 3068 18570 3080
rect 14461 3043 14519 3049
rect 14461 3009 14473 3043
rect 14507 3040 14519 3043
rect 14734 3040 14740 3052
rect 14507 3012 14740 3040
rect 14507 3009 14519 3012
rect 14461 3003 14519 3009
rect 14734 3000 14740 3012
rect 14792 3000 14798 3052
rect 15289 3043 15347 3049
rect 15289 3009 15301 3043
rect 15335 3040 15347 3043
rect 15378 3040 15384 3052
rect 15335 3012 15384 3040
rect 15335 3009 15347 3012
rect 15289 3003 15347 3009
rect 15378 3000 15384 3012
rect 15436 3000 15442 3052
rect 16114 3000 16120 3052
rect 16172 3000 16178 3052
rect 19426 3000 19432 3052
rect 19484 3000 19490 3052
rect 19536 3040 19564 3080
rect 20254 3068 20260 3120
rect 20312 3108 20318 3120
rect 20312 3080 23888 3108
rect 20312 3068 20318 3080
rect 20533 3043 20591 3049
rect 20533 3040 20545 3043
rect 19536 3012 20545 3040
rect 20533 3009 20545 3012
rect 20579 3009 20591 3043
rect 20533 3003 20591 3009
rect 20898 3000 20904 3052
rect 20956 3000 20962 3052
rect 21358 3000 21364 3052
rect 21416 3040 21422 3052
rect 21821 3043 21879 3049
rect 21821 3040 21833 3043
rect 21416 3012 21833 3040
rect 21416 3000 21422 3012
rect 21821 3009 21833 3012
rect 21867 3009 21879 3043
rect 21821 3003 21879 3009
rect 22738 3000 22744 3052
rect 22796 3000 22802 3052
rect 23860 3049 23888 3080
rect 23293 3043 23351 3049
rect 23293 3009 23305 3043
rect 23339 3009 23351 3043
rect 23293 3003 23351 3009
rect 23845 3043 23903 3049
rect 23845 3009 23857 3043
rect 23891 3009 23903 3043
rect 23845 3003 23903 3009
rect 12342 2932 12348 2984
rect 12400 2972 12406 2984
rect 19702 2972 19708 2984
rect 12400 2944 19708 2972
rect 12400 2932 12406 2944
rect 19702 2932 19708 2944
rect 19760 2932 19766 2984
rect 19794 2932 19800 2984
rect 19852 2972 19858 2984
rect 23308 2972 23336 3003
rect 31294 3000 31300 3052
rect 31352 3000 31358 3052
rect 31662 3000 31668 3052
rect 31720 3000 31726 3052
rect 19852 2944 23336 2972
rect 19852 2932 19858 2944
rect 12894 2864 12900 2916
rect 12952 2904 12958 2916
rect 13538 2904 13544 2916
rect 12952 2876 13544 2904
rect 12952 2864 12958 2876
rect 13538 2864 13544 2876
rect 13596 2864 13602 2916
rect 16850 2864 16856 2916
rect 16908 2904 16914 2916
rect 16908 2876 19840 2904
rect 16908 2864 16914 2876
rect 19812 2848 19840 2876
rect 19886 2864 19892 2916
rect 19944 2904 19950 2916
rect 20530 2904 20536 2916
rect 19944 2876 20536 2904
rect 19944 2864 19950 2876
rect 20530 2864 20536 2876
rect 20588 2864 20594 2916
rect 21450 2864 21456 2916
rect 21508 2904 21514 2916
rect 22370 2904 22376 2916
rect 21508 2876 22376 2904
rect 21508 2864 21514 2876
rect 22370 2864 22376 2876
rect 22428 2864 22434 2916
rect 12434 2796 12440 2848
rect 12492 2836 12498 2848
rect 13262 2836 13268 2848
rect 12492 2808 13268 2836
rect 12492 2796 12498 2808
rect 13262 2796 13268 2808
rect 13320 2796 13326 2848
rect 14366 2796 14372 2848
rect 14424 2836 14430 2848
rect 14645 2839 14703 2845
rect 14645 2836 14657 2839
rect 14424 2808 14657 2836
rect 14424 2796 14430 2808
rect 14645 2805 14657 2808
rect 14691 2805 14703 2839
rect 14645 2799 14703 2805
rect 15378 2796 15384 2848
rect 15436 2836 15442 2848
rect 15473 2839 15531 2845
rect 15473 2836 15485 2839
rect 15436 2808 15485 2836
rect 15436 2796 15442 2808
rect 15473 2805 15485 2808
rect 15519 2805 15531 2839
rect 15473 2799 15531 2805
rect 16022 2796 16028 2848
rect 16080 2836 16086 2848
rect 16301 2839 16359 2845
rect 16301 2836 16313 2839
rect 16080 2808 16313 2836
rect 16080 2796 16086 2808
rect 16301 2805 16313 2808
rect 16347 2805 16359 2839
rect 16301 2799 16359 2805
rect 17770 2796 17776 2848
rect 17828 2836 17834 2848
rect 18506 2836 18512 2848
rect 17828 2808 18512 2836
rect 17828 2796 17834 2808
rect 18506 2796 18512 2808
rect 18564 2796 18570 2848
rect 19334 2796 19340 2848
rect 19392 2836 19398 2848
rect 19613 2839 19671 2845
rect 19613 2836 19625 2839
rect 19392 2808 19625 2836
rect 19392 2796 19398 2808
rect 19613 2805 19625 2808
rect 19659 2805 19671 2839
rect 19613 2799 19671 2805
rect 19794 2796 19800 2848
rect 19852 2796 19858 2848
rect 20438 2796 20444 2848
rect 20496 2836 20502 2848
rect 20717 2839 20775 2845
rect 20717 2836 20729 2839
rect 20496 2808 20729 2836
rect 20496 2796 20502 2808
rect 20717 2805 20729 2808
rect 20763 2805 20775 2839
rect 20717 2799 20775 2805
rect 20806 2796 20812 2848
rect 20864 2836 20870 2848
rect 21085 2839 21143 2845
rect 21085 2836 21097 2839
rect 20864 2808 21097 2836
rect 20864 2796 20870 2808
rect 21085 2805 21097 2808
rect 21131 2805 21143 2839
rect 21085 2799 21143 2805
rect 21542 2796 21548 2848
rect 21600 2836 21606 2848
rect 22005 2839 22063 2845
rect 22005 2836 22017 2839
rect 21600 2808 22017 2836
rect 21600 2796 21606 2808
rect 22005 2805 22017 2808
rect 22051 2805 22063 2839
rect 22005 2799 22063 2805
rect 22646 2796 22652 2848
rect 22704 2836 22710 2848
rect 22925 2839 22983 2845
rect 22925 2836 22937 2839
rect 22704 2808 22937 2836
rect 22704 2796 22710 2808
rect 22925 2805 22937 2808
rect 22971 2805 22983 2839
rect 22925 2799 22983 2805
rect 23198 2796 23204 2848
rect 23256 2836 23262 2848
rect 23477 2839 23535 2845
rect 23477 2836 23489 2839
rect 23256 2808 23489 2836
rect 23256 2796 23262 2808
rect 23477 2805 23489 2808
rect 23523 2805 23535 2839
rect 23477 2799 23535 2805
rect 23750 2796 23756 2848
rect 23808 2836 23814 2848
rect 24029 2839 24087 2845
rect 24029 2836 24041 2839
rect 23808 2808 24041 2836
rect 23808 2796 23814 2808
rect 24029 2805 24041 2808
rect 24075 2805 24087 2839
rect 24029 2799 24087 2805
rect 31481 2839 31539 2845
rect 31481 2805 31493 2839
rect 31527 2836 31539 2839
rect 31754 2836 31760 2848
rect 31527 2808 31760 2836
rect 31527 2805 31539 2808
rect 31481 2799 31539 2805
rect 31754 2796 31760 2808
rect 31812 2796 31818 2848
rect 31849 2839 31907 2845
rect 31849 2805 31861 2839
rect 31895 2836 31907 2839
rect 32858 2836 32864 2848
rect 31895 2808 32864 2836
rect 31895 2805 31907 2808
rect 31849 2799 31907 2805
rect 32858 2796 32864 2808
rect 32916 2796 32922 2848
rect 1104 2746 32568 2768
rect 1104 2694 1950 2746
rect 2002 2694 2014 2746
rect 2066 2694 2078 2746
rect 2130 2694 2142 2746
rect 2194 2694 2206 2746
rect 2258 2694 7950 2746
rect 8002 2694 8014 2746
rect 8066 2694 8078 2746
rect 8130 2694 8142 2746
rect 8194 2694 8206 2746
rect 8258 2694 13950 2746
rect 14002 2694 14014 2746
rect 14066 2694 14078 2746
rect 14130 2694 14142 2746
rect 14194 2694 14206 2746
rect 14258 2694 19950 2746
rect 20002 2694 20014 2746
rect 20066 2694 20078 2746
rect 20130 2694 20142 2746
rect 20194 2694 20206 2746
rect 20258 2694 25950 2746
rect 26002 2694 26014 2746
rect 26066 2694 26078 2746
rect 26130 2694 26142 2746
rect 26194 2694 26206 2746
rect 26258 2694 31950 2746
rect 32002 2694 32014 2746
rect 32066 2694 32078 2746
rect 32130 2694 32142 2746
rect 32194 2694 32206 2746
rect 32258 2694 32568 2746
rect 1104 2672 32568 2694
rect 9490 2592 9496 2644
rect 9548 2632 9554 2644
rect 14182 2632 14188 2644
rect 9548 2604 14188 2632
rect 9548 2592 9554 2604
rect 14182 2592 14188 2604
rect 14240 2592 14246 2644
rect 17678 2592 17684 2644
rect 17736 2632 17742 2644
rect 18601 2635 18659 2641
rect 18601 2632 18613 2635
rect 17736 2604 18613 2632
rect 17736 2592 17742 2604
rect 18601 2601 18613 2604
rect 18647 2601 18659 2635
rect 18601 2595 18659 2601
rect 18874 2592 18880 2644
rect 18932 2632 18938 2644
rect 19518 2632 19524 2644
rect 18932 2604 19524 2632
rect 18932 2592 18938 2604
rect 19518 2592 19524 2604
rect 19576 2592 19582 2644
rect 20533 2635 20591 2641
rect 20533 2632 20545 2635
rect 19720 2604 20545 2632
rect 13170 2524 13176 2576
rect 13228 2564 13234 2576
rect 13228 2536 14596 2564
rect 13228 2524 13234 2536
rect 9582 2456 9588 2508
rect 9640 2496 9646 2508
rect 14568 2496 14596 2536
rect 15470 2524 15476 2576
rect 15528 2564 15534 2576
rect 15528 2536 15976 2564
rect 15528 2524 15534 2536
rect 15948 2496 15976 2536
rect 18230 2524 18236 2576
rect 18288 2564 18294 2576
rect 18969 2567 19027 2573
rect 18969 2564 18981 2567
rect 18288 2536 18981 2564
rect 18288 2524 18294 2536
rect 18969 2533 18981 2536
rect 19015 2533 19027 2567
rect 18969 2527 19027 2533
rect 19058 2524 19064 2576
rect 19116 2564 19122 2576
rect 19426 2564 19432 2576
rect 19116 2536 19432 2564
rect 19116 2524 19122 2536
rect 19426 2524 19432 2536
rect 19484 2524 19490 2576
rect 9640 2468 14320 2496
rect 14568 2468 15884 2496
rect 15948 2468 18460 2496
rect 9640 2456 9646 2468
rect 13630 2388 13636 2440
rect 13688 2388 13694 2440
rect 14292 2428 14320 2468
rect 14357 2431 14415 2437
rect 14357 2428 14369 2431
rect 14292 2400 14369 2428
rect 14357 2397 14369 2400
rect 14403 2397 14415 2431
rect 14357 2391 14415 2397
rect 14458 2388 14464 2440
rect 14516 2428 14522 2440
rect 14737 2431 14795 2437
rect 14737 2428 14749 2431
rect 14516 2400 14749 2428
rect 14516 2388 14522 2400
rect 14737 2397 14749 2400
rect 14783 2397 14795 2431
rect 14737 2391 14795 2397
rect 14918 2388 14924 2440
rect 14976 2428 14982 2440
rect 15856 2437 15884 2468
rect 15105 2431 15163 2437
rect 15105 2428 15117 2431
rect 14976 2400 15117 2428
rect 14976 2388 14982 2400
rect 15105 2397 15117 2400
rect 15151 2397 15163 2431
rect 15105 2391 15163 2397
rect 15473 2431 15531 2437
rect 15473 2397 15485 2431
rect 15519 2397 15531 2431
rect 15473 2391 15531 2397
rect 15841 2431 15899 2437
rect 15841 2397 15853 2431
rect 15887 2397 15899 2431
rect 15841 2391 15899 2397
rect 12802 2320 12808 2372
rect 12860 2360 12866 2372
rect 15488 2360 15516 2391
rect 16206 2388 16212 2440
rect 16264 2388 16270 2440
rect 16758 2388 16764 2440
rect 16816 2388 16822 2440
rect 16942 2388 16948 2440
rect 17000 2428 17006 2440
rect 17129 2431 17187 2437
rect 17129 2428 17141 2431
rect 17000 2400 17141 2428
rect 17000 2388 17006 2400
rect 17129 2397 17141 2400
rect 17175 2397 17187 2431
rect 17129 2391 17187 2397
rect 17494 2388 17500 2440
rect 17552 2388 17558 2440
rect 17954 2388 17960 2440
rect 18012 2428 18018 2440
rect 18432 2437 18460 2468
rect 18049 2431 18107 2437
rect 18049 2428 18061 2431
rect 18012 2400 18061 2428
rect 18012 2388 18018 2400
rect 18049 2397 18061 2400
rect 18095 2397 18107 2431
rect 18049 2391 18107 2397
rect 18417 2431 18475 2437
rect 18417 2397 18429 2431
rect 18463 2397 18475 2431
rect 18417 2391 18475 2397
rect 18506 2388 18512 2440
rect 18564 2428 18570 2440
rect 18773 2431 18831 2437
rect 18773 2428 18785 2431
rect 18564 2400 18785 2428
rect 18564 2388 18570 2400
rect 18773 2397 18785 2400
rect 18819 2397 18831 2431
rect 19245 2431 19303 2437
rect 19245 2428 19257 2431
rect 18773 2391 18831 2397
rect 18892 2400 19257 2428
rect 12860 2332 15516 2360
rect 12860 2320 12866 2332
rect 15562 2320 15568 2372
rect 15620 2360 15626 2372
rect 18892 2360 18920 2400
rect 19245 2397 19257 2400
rect 19291 2397 19303 2431
rect 19245 2391 19303 2397
rect 19426 2388 19432 2440
rect 19484 2428 19490 2440
rect 19613 2431 19671 2437
rect 19613 2428 19625 2431
rect 19484 2400 19625 2428
rect 19484 2388 19490 2400
rect 19613 2397 19625 2400
rect 19659 2397 19671 2431
rect 19613 2391 19671 2397
rect 19720 2360 19748 2604
rect 20533 2601 20545 2604
rect 20579 2601 20591 2635
rect 20533 2595 20591 2601
rect 21450 2592 21456 2644
rect 21508 2632 21514 2644
rect 22373 2635 22431 2641
rect 22373 2632 22385 2635
rect 21508 2604 22385 2632
rect 21508 2592 21514 2604
rect 22373 2601 22385 2604
rect 22419 2601 22431 2635
rect 22373 2595 22431 2601
rect 22462 2592 22468 2644
rect 22520 2632 22526 2644
rect 23477 2635 23535 2641
rect 23477 2632 23489 2635
rect 22520 2604 23489 2632
rect 22520 2592 22526 2604
rect 23477 2601 23489 2604
rect 23523 2601 23535 2635
rect 23477 2595 23535 2601
rect 19886 2524 19892 2576
rect 19944 2564 19950 2576
rect 20901 2567 20959 2573
rect 20901 2564 20913 2567
rect 19944 2536 20913 2564
rect 19944 2524 19950 2536
rect 20901 2533 20913 2536
rect 20947 2533 20959 2567
rect 20901 2527 20959 2533
rect 21818 2524 21824 2576
rect 21876 2564 21882 2576
rect 22741 2567 22799 2573
rect 22741 2564 22753 2567
rect 21876 2536 22753 2564
rect 21876 2524 21882 2536
rect 22741 2533 22753 2536
rect 22787 2533 22799 2567
rect 22741 2527 22799 2533
rect 22922 2524 22928 2576
rect 22980 2564 22986 2576
rect 23845 2567 23903 2573
rect 23845 2564 23857 2567
rect 22980 2536 23857 2564
rect 22980 2524 22986 2536
rect 23845 2533 23857 2536
rect 23891 2533 23903 2567
rect 23845 2527 23903 2533
rect 24118 2524 24124 2576
rect 24176 2564 24182 2576
rect 24176 2536 30604 2564
rect 24176 2524 24182 2536
rect 20530 2456 20536 2508
rect 20588 2496 20594 2508
rect 20588 2468 21128 2496
rect 20588 2456 20594 2468
rect 19978 2388 19984 2440
rect 20036 2388 20042 2440
rect 20346 2388 20352 2440
rect 20404 2388 20410 2440
rect 21100 2437 21128 2468
rect 22278 2456 22284 2508
rect 22336 2496 22342 2508
rect 22336 2468 23796 2496
rect 22336 2456 22342 2468
rect 20717 2431 20775 2437
rect 20717 2428 20729 2431
rect 20548 2400 20729 2428
rect 20548 2372 20576 2400
rect 20717 2397 20729 2400
rect 20763 2397 20775 2431
rect 20717 2391 20775 2397
rect 21085 2431 21143 2437
rect 21085 2397 21097 2431
rect 21131 2397 21143 2431
rect 21085 2391 21143 2397
rect 21634 2388 21640 2440
rect 21692 2428 21698 2440
rect 21821 2431 21879 2437
rect 21821 2428 21833 2431
rect 21692 2400 21833 2428
rect 21692 2388 21698 2400
rect 21821 2397 21833 2400
rect 21867 2397 21879 2431
rect 22189 2431 22247 2437
rect 22189 2428 22201 2431
rect 21821 2391 21879 2397
rect 22066 2400 22201 2428
rect 15620 2332 18920 2360
rect 19628 2332 19748 2360
rect 15620 2320 15626 2332
rect 19628 2304 19656 2332
rect 20530 2320 20536 2372
rect 20588 2320 20594 2372
rect 20622 2320 20628 2372
rect 20680 2360 20686 2372
rect 22066 2360 22094 2400
rect 22189 2397 22201 2400
rect 22235 2397 22247 2431
rect 22189 2391 22247 2397
rect 22370 2388 22376 2440
rect 22428 2428 22434 2440
rect 22557 2431 22615 2437
rect 22557 2428 22569 2431
rect 22428 2400 22569 2428
rect 22428 2388 22434 2400
rect 22557 2397 22569 2400
rect 22603 2397 22615 2431
rect 22557 2391 22615 2397
rect 22738 2388 22744 2440
rect 22796 2428 22802 2440
rect 22925 2431 22983 2437
rect 22925 2428 22937 2431
rect 22796 2400 22937 2428
rect 22796 2388 22802 2400
rect 22925 2397 22937 2400
rect 22971 2397 22983 2431
rect 22925 2391 22983 2397
rect 23290 2388 23296 2440
rect 23348 2388 23354 2440
rect 23658 2388 23664 2440
rect 23716 2388 23722 2440
rect 23768 2428 23796 2468
rect 23934 2456 23940 2508
rect 23992 2496 23998 2508
rect 23992 2468 26234 2496
rect 23992 2456 23998 2468
rect 24397 2431 24455 2437
rect 24397 2428 24409 2431
rect 23768 2400 24409 2428
rect 24397 2397 24409 2400
rect 24443 2397 24455 2431
rect 24397 2391 24455 2397
rect 20680 2332 22094 2360
rect 26206 2360 26234 2468
rect 30576 2437 30604 2536
rect 30561 2431 30619 2437
rect 30561 2397 30573 2431
rect 30607 2397 30619 2431
rect 30561 2391 30619 2397
rect 30926 2388 30932 2440
rect 30984 2388 30990 2440
rect 31294 2388 31300 2440
rect 31352 2388 31358 2440
rect 31665 2431 31723 2437
rect 31665 2397 31677 2431
rect 31711 2397 31723 2431
rect 31665 2391 31723 2397
rect 31680 2360 31708 2391
rect 26206 2332 31708 2360
rect 20680 2320 20686 2332
rect 13817 2295 13875 2301
rect 13817 2261 13829 2295
rect 13863 2292 13875 2295
rect 14090 2292 14096 2304
rect 13863 2264 14096 2292
rect 13863 2261 13875 2264
rect 13817 2255 13875 2261
rect 14090 2252 14096 2264
rect 14148 2252 14154 2304
rect 14182 2252 14188 2304
rect 14240 2292 14246 2304
rect 14458 2292 14464 2304
rect 14240 2264 14464 2292
rect 14240 2252 14246 2264
rect 14458 2252 14464 2264
rect 14516 2252 14522 2304
rect 14553 2295 14611 2301
rect 14553 2261 14565 2295
rect 14599 2292 14611 2295
rect 14642 2292 14648 2304
rect 14599 2264 14648 2292
rect 14599 2261 14611 2264
rect 14553 2255 14611 2261
rect 14642 2252 14648 2264
rect 14700 2252 14706 2304
rect 14918 2252 14924 2304
rect 14976 2252 14982 2304
rect 15289 2295 15347 2301
rect 15289 2261 15301 2295
rect 15335 2292 15347 2295
rect 15470 2292 15476 2304
rect 15335 2264 15476 2292
rect 15335 2261 15347 2264
rect 15289 2255 15347 2261
rect 15470 2252 15476 2264
rect 15528 2252 15534 2304
rect 15657 2295 15715 2301
rect 15657 2261 15669 2295
rect 15703 2292 15715 2295
rect 15746 2292 15752 2304
rect 15703 2264 15752 2292
rect 15703 2261 15715 2264
rect 15657 2255 15715 2261
rect 15746 2252 15752 2264
rect 15804 2252 15810 2304
rect 16025 2295 16083 2301
rect 16025 2261 16037 2295
rect 16071 2292 16083 2295
rect 16298 2292 16304 2304
rect 16071 2264 16304 2292
rect 16071 2261 16083 2264
rect 16025 2255 16083 2261
rect 16298 2252 16304 2264
rect 16356 2252 16362 2304
rect 16393 2295 16451 2301
rect 16393 2261 16405 2295
rect 16439 2292 16451 2295
rect 16574 2292 16580 2304
rect 16439 2264 16580 2292
rect 16439 2261 16451 2264
rect 16393 2255 16451 2261
rect 16574 2252 16580 2264
rect 16632 2252 16638 2304
rect 16850 2252 16856 2304
rect 16908 2292 16914 2304
rect 16945 2295 17003 2301
rect 16945 2292 16957 2295
rect 16908 2264 16957 2292
rect 16908 2252 16914 2264
rect 16945 2261 16957 2264
rect 16991 2261 17003 2295
rect 16945 2255 17003 2261
rect 17126 2252 17132 2304
rect 17184 2292 17190 2304
rect 17313 2295 17371 2301
rect 17313 2292 17325 2295
rect 17184 2264 17325 2292
rect 17184 2252 17190 2264
rect 17313 2261 17325 2264
rect 17359 2261 17371 2295
rect 17313 2255 17371 2261
rect 17402 2252 17408 2304
rect 17460 2292 17466 2304
rect 17681 2295 17739 2301
rect 17681 2292 17693 2295
rect 17460 2264 17693 2292
rect 17460 2252 17466 2264
rect 17681 2261 17693 2264
rect 17727 2261 17739 2295
rect 17681 2255 17739 2261
rect 17954 2252 17960 2304
rect 18012 2292 18018 2304
rect 18233 2295 18291 2301
rect 18233 2292 18245 2295
rect 18012 2264 18245 2292
rect 18012 2252 18018 2264
rect 18233 2261 18245 2264
rect 18279 2261 18291 2295
rect 18233 2255 18291 2261
rect 18506 2252 18512 2304
rect 18564 2292 18570 2304
rect 19429 2295 19487 2301
rect 19429 2292 19441 2295
rect 18564 2264 19441 2292
rect 18564 2252 18570 2264
rect 19429 2261 19441 2264
rect 19475 2261 19487 2295
rect 19429 2255 19487 2261
rect 19610 2252 19616 2304
rect 19668 2252 19674 2304
rect 19702 2252 19708 2304
rect 19760 2292 19766 2304
rect 19797 2295 19855 2301
rect 19797 2292 19809 2295
rect 19760 2264 19809 2292
rect 19760 2252 19766 2264
rect 19797 2261 19809 2264
rect 19843 2261 19855 2295
rect 19797 2255 19855 2261
rect 20162 2252 20168 2304
rect 20220 2252 20226 2304
rect 20254 2252 20260 2304
rect 20312 2292 20318 2304
rect 21269 2295 21327 2301
rect 21269 2292 21281 2295
rect 20312 2264 21281 2292
rect 20312 2252 20318 2264
rect 21269 2261 21281 2264
rect 21315 2261 21327 2295
rect 21269 2255 21327 2261
rect 21358 2252 21364 2304
rect 21416 2292 21422 2304
rect 22005 2295 22063 2301
rect 22005 2292 22017 2295
rect 21416 2264 22017 2292
rect 21416 2252 21422 2264
rect 22005 2261 22017 2264
rect 22051 2261 22063 2295
rect 22005 2255 22063 2261
rect 22094 2252 22100 2304
rect 22152 2292 22158 2304
rect 23109 2295 23167 2301
rect 23109 2292 23121 2295
rect 22152 2264 23121 2292
rect 22152 2252 22158 2264
rect 23109 2261 23121 2264
rect 23155 2261 23167 2295
rect 23109 2255 23167 2261
rect 23566 2252 23572 2304
rect 23624 2292 23630 2304
rect 24581 2295 24639 2301
rect 24581 2292 24593 2295
rect 23624 2264 24593 2292
rect 23624 2252 23630 2264
rect 24581 2261 24593 2264
rect 24627 2261 24639 2295
rect 24581 2255 24639 2261
rect 30742 2252 30748 2304
rect 30800 2252 30806 2304
rect 31110 2252 31116 2304
rect 31168 2252 31174 2304
rect 31478 2252 31484 2304
rect 31536 2252 31542 2304
rect 31846 2252 31852 2304
rect 31904 2252 31910 2304
rect 1104 2202 32568 2224
rect 1104 2150 3010 2202
rect 3062 2150 3074 2202
rect 3126 2150 3138 2202
rect 3190 2150 3202 2202
rect 3254 2150 3266 2202
rect 3318 2150 9010 2202
rect 9062 2150 9074 2202
rect 9126 2150 9138 2202
rect 9190 2150 9202 2202
rect 9254 2150 9266 2202
rect 9318 2150 15010 2202
rect 15062 2150 15074 2202
rect 15126 2150 15138 2202
rect 15190 2150 15202 2202
rect 15254 2150 15266 2202
rect 15318 2150 21010 2202
rect 21062 2150 21074 2202
rect 21126 2150 21138 2202
rect 21190 2150 21202 2202
rect 21254 2150 21266 2202
rect 21318 2150 27010 2202
rect 27062 2150 27074 2202
rect 27126 2150 27138 2202
rect 27190 2150 27202 2202
rect 27254 2150 27266 2202
rect 27318 2150 32568 2202
rect 1104 2128 32568 2150
rect 11330 2048 11336 2100
rect 11388 2088 11394 2100
rect 14274 2088 14280 2100
rect 11388 2060 14280 2088
rect 11388 2048 11394 2060
rect 14274 2048 14280 2060
rect 14332 2048 14338 2100
rect 17862 2048 17868 2100
rect 17920 2088 17926 2100
rect 21634 2088 21640 2100
rect 17920 2060 21640 2088
rect 17920 2048 17926 2060
rect 21634 2048 21640 2060
rect 21692 2048 21698 2100
rect 22002 2048 22008 2100
rect 22060 2088 22066 2100
rect 23658 2088 23664 2100
rect 22060 2060 23664 2088
rect 22060 2048 22066 2060
rect 23658 2048 23664 2060
rect 23716 2048 23722 2100
rect 9674 1980 9680 2032
rect 9732 2020 9738 2032
rect 18874 2020 18880 2032
rect 9732 1992 14320 2020
rect 9732 1980 9738 1992
rect 6178 1912 6184 1964
rect 6236 1952 6242 1964
rect 14292 1952 14320 1992
rect 14568 1992 18880 2020
rect 14568 1952 14596 1992
rect 18874 1980 18880 1992
rect 18932 1980 18938 2032
rect 18966 1980 18972 2032
rect 19024 2020 19030 2032
rect 19702 2020 19708 2032
rect 19024 1992 19708 2020
rect 19024 1980 19030 1992
rect 19702 1980 19708 1992
rect 19760 1980 19766 2032
rect 19794 1980 19800 2032
rect 19852 2020 19858 2032
rect 23290 2020 23296 2032
rect 19852 1992 23296 2020
rect 19852 1980 19858 1992
rect 23290 1980 23296 1992
rect 23348 1980 23354 2032
rect 6236 1924 12434 1952
rect 14292 1924 14596 1952
rect 6236 1912 6242 1924
rect 12406 1884 12434 1924
rect 15930 1912 15936 1964
rect 15988 1952 15994 1964
rect 20346 1952 20352 1964
rect 15988 1924 20352 1952
rect 15988 1912 15994 1924
rect 20346 1912 20352 1924
rect 20404 1912 20410 1964
rect 19978 1884 19984 1896
rect 12406 1856 19984 1884
rect 19978 1844 19984 1856
rect 20036 1844 20042 1896
rect 22738 1884 22744 1896
rect 22066 1856 22744 1884
rect 8386 1776 8392 1828
rect 8444 1816 8450 1828
rect 19426 1816 19432 1828
rect 8444 1788 19432 1816
rect 8444 1776 8450 1788
rect 19426 1776 19432 1788
rect 19484 1776 19490 1828
rect 9950 1708 9956 1760
rect 10008 1748 10014 1760
rect 19058 1748 19064 1760
rect 10008 1720 19064 1748
rect 10008 1708 10014 1720
rect 19058 1708 19064 1720
rect 19116 1708 19122 1760
rect 19150 1708 19156 1760
rect 19208 1748 19214 1760
rect 22066 1748 22094 1856
rect 22738 1844 22744 1856
rect 22796 1844 22802 1896
rect 19208 1720 22094 1748
rect 19208 1708 19214 1720
rect 10134 1640 10140 1692
rect 10192 1680 10198 1692
rect 16942 1680 16948 1692
rect 10192 1652 16948 1680
rect 10192 1640 10198 1652
rect 16942 1640 16948 1652
rect 17000 1640 17006 1692
rect 18690 1640 18696 1692
rect 18748 1680 18754 1692
rect 31294 1680 31300 1692
rect 18748 1652 31300 1680
rect 18748 1640 18754 1652
rect 31294 1640 31300 1652
rect 31352 1640 31358 1692
rect 13354 1572 13360 1624
rect 13412 1612 13418 1624
rect 16206 1612 16212 1624
rect 13412 1584 16212 1612
rect 13412 1572 13418 1584
rect 16206 1572 16212 1584
rect 16264 1572 16270 1624
rect 19058 1368 19064 1420
rect 19116 1408 19122 1420
rect 20162 1408 20168 1420
rect 19116 1380 20168 1408
rect 19116 1368 19122 1380
rect 20162 1368 20168 1380
rect 20220 1368 20226 1420
rect 9490 1300 9496 1352
rect 9548 1340 9554 1352
rect 14550 1340 14556 1352
rect 9548 1312 14556 1340
rect 9548 1300 9554 1312
rect 14550 1300 14556 1312
rect 14608 1300 14614 1352
rect 19518 1300 19524 1352
rect 19576 1340 19582 1352
rect 25406 1340 25412 1352
rect 19576 1312 25412 1340
rect 19576 1300 19582 1312
rect 25406 1300 25412 1312
rect 25464 1300 25470 1352
rect 11054 1232 11060 1284
rect 11112 1272 11118 1284
rect 16666 1272 16672 1284
rect 11112 1244 16672 1272
rect 11112 1232 11118 1244
rect 16666 1232 16672 1244
rect 16724 1232 16730 1284
rect 22830 1096 22836 1148
rect 22888 1136 22894 1148
rect 27062 1136 27068 1148
rect 22888 1108 27068 1136
rect 22888 1096 22894 1108
rect 27062 1096 27068 1108
rect 27120 1096 27126 1148
<< via1 >>
rect 16764 9392 16816 9444
rect 24952 9392 25004 9444
rect 17316 9324 17368 9376
rect 25320 9324 25372 9376
rect 14280 9256 14332 9308
rect 30656 9256 30708 9308
rect 9404 9188 9456 9240
rect 19524 9188 19576 9240
rect 12532 9120 12584 9172
rect 17316 9120 17368 9172
rect 17408 9120 17460 9172
rect 24216 9120 24268 9172
rect 12624 9052 12676 9104
rect 30288 9052 30340 9104
rect 17868 8984 17920 9036
rect 4988 8916 5040 8968
rect 17408 8916 17460 8968
rect 17500 8916 17552 8968
rect 29920 8916 29972 8968
rect 10968 8848 11020 8900
rect 4712 8780 4764 8832
rect 14372 8780 14424 8832
rect 16764 8780 16816 8832
rect 17040 8848 17092 8900
rect 23388 8848 23440 8900
rect 22928 8780 22980 8832
rect 3010 8678 3062 8730
rect 3074 8678 3126 8730
rect 3138 8678 3190 8730
rect 3202 8678 3254 8730
rect 3266 8678 3318 8730
rect 9010 8678 9062 8730
rect 9074 8678 9126 8730
rect 9138 8678 9190 8730
rect 9202 8678 9254 8730
rect 9266 8678 9318 8730
rect 15010 8678 15062 8730
rect 15074 8678 15126 8730
rect 15138 8678 15190 8730
rect 15202 8678 15254 8730
rect 15266 8678 15318 8730
rect 21010 8678 21062 8730
rect 21074 8678 21126 8730
rect 21138 8678 21190 8730
rect 21202 8678 21254 8730
rect 21266 8678 21318 8730
rect 27010 8678 27062 8730
rect 27074 8678 27126 8730
rect 27138 8678 27190 8730
rect 27202 8678 27254 8730
rect 27266 8678 27318 8730
rect 1216 8576 1268 8628
rect 2780 8576 2832 8628
rect 4344 8576 4396 8628
rect 4712 8576 4764 8628
rect 5908 8576 5960 8628
rect 7472 8576 7524 8628
rect 8852 8576 8904 8628
rect 10600 8576 10652 8628
rect 1584 8483 1636 8492
rect 1584 8449 1593 8483
rect 1593 8449 1627 8483
rect 1627 8449 1636 8483
rect 1584 8440 1636 8449
rect 12072 8576 12124 8628
rect 12164 8576 12216 8628
rect 13728 8576 13780 8628
rect 15384 8576 15436 8628
rect 16856 8576 16908 8628
rect 18420 8576 18472 8628
rect 19984 8576 20036 8628
rect 21548 8576 21600 8628
rect 23112 8576 23164 8628
rect 24676 8576 24728 8628
rect 26240 8576 26292 8628
rect 27804 8576 27856 8628
rect 29368 8576 29420 8628
rect 30104 8619 30156 8628
rect 30104 8585 30113 8619
rect 30113 8585 30147 8619
rect 30147 8585 30156 8619
rect 30104 8576 30156 8585
rect 30472 8619 30524 8628
rect 30472 8585 30481 8619
rect 30481 8585 30515 8619
rect 30515 8585 30524 8619
rect 30472 8576 30524 8585
rect 30932 8576 30984 8628
rect 4988 8372 5040 8424
rect 9404 8483 9456 8492
rect 9404 8449 9413 8483
rect 9413 8449 9447 8483
rect 9447 8449 9456 8483
rect 9404 8440 9456 8449
rect 10968 8483 11020 8492
rect 10968 8449 10977 8483
rect 10977 8449 11011 8483
rect 11011 8449 11020 8483
rect 10968 8440 11020 8449
rect 12532 8483 12584 8492
rect 12532 8449 12541 8483
rect 12541 8449 12575 8483
rect 12575 8449 12584 8483
rect 12532 8440 12584 8449
rect 14372 8483 14424 8492
rect 14372 8449 14381 8483
rect 14381 8449 14415 8483
rect 14415 8449 14424 8483
rect 14372 8440 14424 8449
rect 15660 8483 15712 8492
rect 15660 8449 15662 8483
rect 15662 8449 15696 8483
rect 15696 8449 15712 8483
rect 15660 8440 15712 8449
rect 19156 8508 19208 8560
rect 15844 8372 15896 8424
rect 17040 8372 17092 8424
rect 18788 8483 18840 8492
rect 18788 8449 18797 8483
rect 18797 8449 18831 8483
rect 18831 8449 18840 8483
rect 18788 8440 18840 8449
rect 20352 8483 20404 8492
rect 20352 8449 20361 8483
rect 20361 8449 20395 8483
rect 20395 8449 20404 8483
rect 20352 8440 20404 8449
rect 20536 8372 20588 8424
rect 14924 8304 14976 8356
rect 22192 8440 22244 8492
rect 23112 8440 23164 8492
rect 23664 8440 23716 8492
rect 26424 8440 26476 8492
rect 25044 8372 25096 8424
rect 29000 8440 29052 8492
rect 29920 8483 29972 8492
rect 29920 8449 29929 8483
rect 29929 8449 29963 8483
rect 29963 8449 29972 8483
rect 29920 8440 29972 8449
rect 30288 8483 30340 8492
rect 30288 8449 30297 8483
rect 30297 8449 30331 8483
rect 30331 8449 30340 8483
rect 30288 8440 30340 8449
rect 30656 8483 30708 8492
rect 30656 8449 30665 8483
rect 30665 8449 30699 8483
rect 30699 8449 30708 8483
rect 30656 8440 30708 8449
rect 30472 8372 30524 8424
rect 32404 8372 32456 8424
rect 31852 8347 31904 8356
rect 31852 8313 31861 8347
rect 31861 8313 31895 8347
rect 31895 8313 31904 8347
rect 31852 8304 31904 8313
rect 1950 8134 2002 8186
rect 2014 8134 2066 8186
rect 2078 8134 2130 8186
rect 2142 8134 2194 8186
rect 2206 8134 2258 8186
rect 7950 8134 8002 8186
rect 8014 8134 8066 8186
rect 8078 8134 8130 8186
rect 8142 8134 8194 8186
rect 8206 8134 8258 8186
rect 13950 8134 14002 8186
rect 14014 8134 14066 8186
rect 14078 8134 14130 8186
rect 14142 8134 14194 8186
rect 14206 8134 14258 8186
rect 19950 8134 20002 8186
rect 20014 8134 20066 8186
rect 20078 8134 20130 8186
rect 20142 8134 20194 8186
rect 20206 8134 20258 8186
rect 25950 8134 26002 8186
rect 26014 8134 26066 8186
rect 26078 8134 26130 8186
rect 26142 8134 26194 8186
rect 26206 8134 26258 8186
rect 31950 8134 32002 8186
rect 32014 8134 32066 8186
rect 32078 8134 32130 8186
rect 32142 8134 32194 8186
rect 32206 8134 32258 8186
rect 4896 7964 4948 8016
rect 15568 8032 15620 8084
rect 21640 8032 21692 8084
rect 30380 8032 30432 8084
rect 30840 8032 30892 8084
rect 31024 8075 31076 8084
rect 31024 8041 31033 8075
rect 31033 8041 31067 8075
rect 31067 8041 31076 8075
rect 31024 8032 31076 8041
rect 31392 8075 31444 8084
rect 31392 8041 31401 8075
rect 31401 8041 31435 8075
rect 31435 8041 31444 8075
rect 31392 8032 31444 8041
rect 7012 7964 7064 8016
rect 7656 7896 7708 7948
rect 13360 7896 13412 7948
rect 7564 7828 7616 7880
rect 15476 7828 15528 7880
rect 7380 7760 7432 7812
rect 12164 7760 12216 7812
rect 19156 7964 19208 8016
rect 20260 7964 20312 8016
rect 26792 7964 26844 8016
rect 16396 7896 16448 7948
rect 18144 7828 18196 7880
rect 21640 7828 21692 7880
rect 23940 7828 23992 7880
rect 30840 7871 30892 7880
rect 30840 7837 30849 7871
rect 30849 7837 30883 7871
rect 30883 7837 30892 7871
rect 30840 7828 30892 7837
rect 5632 7692 5684 7744
rect 8116 7692 8168 7744
rect 12072 7692 12124 7744
rect 14280 7692 14332 7744
rect 16856 7692 16908 7744
rect 26792 7692 26844 7744
rect 31760 7735 31812 7744
rect 31760 7701 31769 7735
rect 31769 7701 31803 7735
rect 31803 7701 31812 7735
rect 31760 7692 31812 7701
rect 32128 7735 32180 7744
rect 32128 7701 32137 7735
rect 32137 7701 32171 7735
rect 32171 7701 32180 7735
rect 32128 7692 32180 7701
rect 3010 7590 3062 7642
rect 3074 7590 3126 7642
rect 3138 7590 3190 7642
rect 3202 7590 3254 7642
rect 3266 7590 3318 7642
rect 9010 7590 9062 7642
rect 9074 7590 9126 7642
rect 9138 7590 9190 7642
rect 9202 7590 9254 7642
rect 9266 7590 9318 7642
rect 15010 7590 15062 7642
rect 15074 7590 15126 7642
rect 15138 7590 15190 7642
rect 15202 7590 15254 7642
rect 15266 7590 15318 7642
rect 21010 7590 21062 7642
rect 21074 7590 21126 7642
rect 21138 7590 21190 7642
rect 21202 7590 21254 7642
rect 21266 7590 21318 7642
rect 27010 7590 27062 7642
rect 27074 7590 27126 7642
rect 27138 7590 27190 7642
rect 27202 7590 27254 7642
rect 27266 7590 27318 7642
rect 4896 7531 4948 7540
rect 4896 7497 4905 7531
rect 4905 7497 4939 7531
rect 4939 7497 4948 7531
rect 4896 7488 4948 7497
rect 6092 7488 6144 7540
rect 5540 7420 5592 7472
rect 7564 7488 7616 7540
rect 12624 7488 12676 7540
rect 13360 7531 13412 7540
rect 13360 7497 13369 7531
rect 13369 7497 13403 7531
rect 13403 7497 13412 7531
rect 13360 7488 13412 7497
rect 13728 7488 13780 7540
rect 15384 7488 15436 7540
rect 16396 7531 16448 7540
rect 16396 7497 16405 7531
rect 16405 7497 16439 7531
rect 16439 7497 16448 7531
rect 16396 7488 16448 7497
rect 16580 7488 16632 7540
rect 18144 7531 18196 7540
rect 18144 7497 18153 7531
rect 18153 7497 18187 7531
rect 18187 7497 18196 7531
rect 18144 7488 18196 7497
rect 4712 7395 4764 7404
rect 4712 7361 4721 7395
rect 4721 7361 4755 7395
rect 4755 7361 4764 7395
rect 4712 7352 4764 7361
rect 4804 7352 4856 7404
rect 6828 7395 6880 7404
rect 6828 7361 6837 7395
rect 6837 7361 6871 7395
rect 6871 7361 6880 7395
rect 6828 7352 6880 7361
rect 8116 7420 8168 7472
rect 7104 7284 7156 7336
rect 7840 7284 7892 7336
rect 5908 7259 5960 7268
rect 5908 7225 5917 7259
rect 5917 7225 5951 7259
rect 5951 7225 5960 7259
rect 5908 7216 5960 7225
rect 6276 7216 6328 7268
rect 6184 7191 6236 7200
rect 6184 7157 6193 7191
rect 6193 7157 6227 7191
rect 6227 7157 6236 7191
rect 6184 7148 6236 7157
rect 7012 7191 7064 7200
rect 7012 7157 7021 7191
rect 7021 7157 7055 7191
rect 7055 7157 7064 7191
rect 7012 7148 7064 7157
rect 7380 7191 7432 7200
rect 7380 7157 7389 7191
rect 7389 7157 7423 7191
rect 7423 7157 7432 7191
rect 7380 7148 7432 7157
rect 7748 7148 7800 7200
rect 11888 7395 11940 7404
rect 11888 7361 11897 7395
rect 11897 7361 11931 7395
rect 11931 7361 11940 7395
rect 11888 7352 11940 7361
rect 12164 7395 12216 7404
rect 12164 7361 12173 7395
rect 12173 7361 12207 7395
rect 12207 7361 12216 7395
rect 12164 7352 12216 7361
rect 12440 7395 12492 7404
rect 12440 7361 12449 7395
rect 12449 7361 12483 7395
rect 12483 7361 12492 7395
rect 12440 7352 12492 7361
rect 13912 7420 13964 7472
rect 14464 7395 14516 7404
rect 14464 7361 14483 7395
rect 14483 7361 14516 7395
rect 14464 7352 14516 7361
rect 14556 7395 14608 7404
rect 14556 7361 14565 7395
rect 14565 7361 14599 7395
rect 14599 7361 14608 7395
rect 14556 7352 14608 7361
rect 16304 7352 16356 7404
rect 17132 7463 17184 7472
rect 17132 7429 17141 7463
rect 17141 7429 17175 7463
rect 17175 7429 17184 7463
rect 17132 7420 17184 7429
rect 19524 7420 19576 7472
rect 20260 7531 20312 7540
rect 20260 7497 20269 7531
rect 20269 7497 20303 7531
rect 20303 7497 20312 7531
rect 20260 7488 20312 7497
rect 9312 7216 9364 7268
rect 10968 7216 11020 7268
rect 16396 7284 16448 7336
rect 19616 7352 19668 7404
rect 21640 7488 21692 7540
rect 22928 7531 22980 7540
rect 22928 7497 22937 7531
rect 22937 7497 22971 7531
rect 22971 7497 22980 7531
rect 22928 7488 22980 7497
rect 24216 7531 24268 7540
rect 24216 7497 24225 7531
rect 24225 7497 24259 7531
rect 24259 7497 24268 7531
rect 24216 7488 24268 7497
rect 25136 7531 25188 7540
rect 25136 7497 25145 7531
rect 25145 7497 25179 7531
rect 25179 7497 25188 7531
rect 25136 7488 25188 7497
rect 25320 7531 25372 7540
rect 25320 7497 25329 7531
rect 25329 7497 25363 7531
rect 25363 7497 25372 7531
rect 25320 7488 25372 7497
rect 31484 7531 31536 7540
rect 31484 7497 31493 7531
rect 31493 7497 31527 7531
rect 31527 7497 31536 7531
rect 31484 7488 31536 7497
rect 20904 7395 20956 7404
rect 20904 7361 20913 7395
rect 20913 7361 20947 7395
rect 20947 7361 20956 7395
rect 20904 7352 20956 7361
rect 25688 7420 25740 7472
rect 24308 7352 24360 7404
rect 23940 7284 23992 7336
rect 24032 7284 24084 7336
rect 25872 7352 25924 7404
rect 31300 7395 31352 7404
rect 31300 7361 31309 7395
rect 31309 7361 31343 7395
rect 31343 7361 31352 7395
rect 31300 7352 31352 7361
rect 15384 7216 15436 7268
rect 15476 7216 15528 7268
rect 9220 7191 9272 7200
rect 9220 7157 9229 7191
rect 9229 7157 9263 7191
rect 9263 7157 9272 7191
rect 9220 7148 9272 7157
rect 9496 7191 9548 7200
rect 9496 7157 9505 7191
rect 9505 7157 9539 7191
rect 9539 7157 9548 7191
rect 9496 7148 9548 7157
rect 12072 7191 12124 7200
rect 12072 7157 12081 7191
rect 12081 7157 12115 7191
rect 12115 7157 12124 7191
rect 12072 7148 12124 7157
rect 12348 7191 12400 7200
rect 12348 7157 12357 7191
rect 12357 7157 12391 7191
rect 12391 7157 12400 7191
rect 12348 7148 12400 7157
rect 12532 7148 12584 7200
rect 12716 7191 12768 7200
rect 12716 7157 12725 7191
rect 12725 7157 12759 7191
rect 12759 7157 12768 7191
rect 12716 7148 12768 7157
rect 13084 7191 13136 7200
rect 13084 7157 13093 7191
rect 13093 7157 13127 7191
rect 13127 7157 13136 7191
rect 13084 7148 13136 7157
rect 14188 7191 14240 7200
rect 14188 7157 14197 7191
rect 14197 7157 14231 7191
rect 14231 7157 14240 7191
rect 14188 7148 14240 7157
rect 14280 7191 14332 7200
rect 14280 7157 14289 7191
rect 14289 7157 14323 7191
rect 14323 7157 14332 7191
rect 14280 7148 14332 7157
rect 14924 7191 14976 7200
rect 14924 7157 14933 7191
rect 14933 7157 14967 7191
rect 14967 7157 14976 7191
rect 14924 7148 14976 7157
rect 16856 7191 16908 7200
rect 16856 7157 16865 7191
rect 16865 7157 16899 7191
rect 16899 7157 16908 7191
rect 16856 7148 16908 7157
rect 17500 7191 17552 7200
rect 17500 7157 17509 7191
rect 17509 7157 17543 7191
rect 17543 7157 17552 7191
rect 17500 7148 17552 7157
rect 17868 7148 17920 7200
rect 32772 7148 32824 7200
rect 1950 7046 2002 7098
rect 2014 7046 2066 7098
rect 2078 7046 2130 7098
rect 2142 7046 2194 7098
rect 2206 7046 2258 7098
rect 7950 7046 8002 7098
rect 8014 7046 8066 7098
rect 8078 7046 8130 7098
rect 8142 7046 8194 7098
rect 8206 7046 8258 7098
rect 13950 7046 14002 7098
rect 14014 7046 14066 7098
rect 14078 7046 14130 7098
rect 14142 7046 14194 7098
rect 14206 7046 14258 7098
rect 19950 7046 20002 7098
rect 20014 7046 20066 7098
rect 20078 7046 20130 7098
rect 20142 7046 20194 7098
rect 20206 7046 20258 7098
rect 25950 7046 26002 7098
rect 26014 7046 26066 7098
rect 26078 7046 26130 7098
rect 26142 7046 26194 7098
rect 26206 7046 26258 7098
rect 31950 7046 32002 7098
rect 32014 7046 32066 7098
rect 32078 7046 32130 7098
rect 32142 7046 32194 7098
rect 32206 7046 32258 7098
rect 4712 6944 4764 6996
rect 7472 6944 7524 6996
rect 12348 6944 12400 6996
rect 30840 6944 30892 6996
rect 7104 6876 7156 6928
rect 7748 6876 7800 6928
rect 9220 6876 9272 6928
rect 16304 6876 16356 6928
rect 20904 6876 20956 6928
rect 24584 6876 24636 6928
rect 9312 6808 9364 6860
rect 17040 6808 17092 6860
rect 5816 6740 5868 6792
rect 4712 6672 4764 6724
rect 8300 6740 8352 6792
rect 6368 6672 6420 6724
rect 5908 6647 5960 6656
rect 5908 6613 5917 6647
rect 5917 6613 5951 6647
rect 5951 6613 5960 6647
rect 5908 6604 5960 6613
rect 8208 6647 8260 6656
rect 8208 6613 8217 6647
rect 8217 6613 8251 6647
rect 8251 6613 8260 6647
rect 8208 6604 8260 6613
rect 15568 6740 15620 6792
rect 16488 6740 16540 6792
rect 17224 6783 17276 6792
rect 17224 6749 17233 6783
rect 17233 6749 17267 6783
rect 17267 6749 17276 6783
rect 17224 6740 17276 6749
rect 26332 6740 26384 6792
rect 31576 6783 31628 6792
rect 31576 6749 31585 6783
rect 31585 6749 31619 6783
rect 31619 6749 31628 6783
rect 31576 6740 31628 6749
rect 31668 6740 31720 6792
rect 9496 6672 9548 6724
rect 31484 6672 31536 6724
rect 16120 6604 16172 6656
rect 16948 6604 17000 6656
rect 17224 6604 17276 6656
rect 19248 6604 19300 6656
rect 19340 6647 19392 6656
rect 19340 6613 19349 6647
rect 19349 6613 19383 6647
rect 19383 6613 19392 6647
rect 19340 6604 19392 6613
rect 19708 6647 19760 6656
rect 19708 6613 19717 6647
rect 19717 6613 19751 6647
rect 19751 6613 19760 6647
rect 19708 6604 19760 6613
rect 24952 6604 25004 6656
rect 31392 6647 31444 6656
rect 31392 6613 31401 6647
rect 31401 6613 31435 6647
rect 31435 6613 31444 6647
rect 31392 6604 31444 6613
rect 31760 6647 31812 6656
rect 31760 6613 31769 6647
rect 31769 6613 31803 6647
rect 31803 6613 31812 6647
rect 31760 6604 31812 6613
rect 32312 6604 32364 6656
rect 3010 6502 3062 6554
rect 3074 6502 3126 6554
rect 3138 6502 3190 6554
rect 3202 6502 3254 6554
rect 3266 6502 3318 6554
rect 9010 6502 9062 6554
rect 9074 6502 9126 6554
rect 9138 6502 9190 6554
rect 9202 6502 9254 6554
rect 9266 6502 9318 6554
rect 15010 6502 15062 6554
rect 15074 6502 15126 6554
rect 15138 6502 15190 6554
rect 15202 6502 15254 6554
rect 15266 6502 15318 6554
rect 21010 6502 21062 6554
rect 21074 6502 21126 6554
rect 21138 6502 21190 6554
rect 21202 6502 21254 6554
rect 21266 6502 21318 6554
rect 27010 6502 27062 6554
rect 27074 6502 27126 6554
rect 27138 6502 27190 6554
rect 27202 6502 27254 6554
rect 27266 6502 27318 6554
rect 8208 6400 8260 6452
rect 14740 6400 14792 6452
rect 19708 6400 19760 6452
rect 27620 6400 27672 6452
rect 31852 6443 31904 6452
rect 31852 6409 31861 6443
rect 31861 6409 31895 6443
rect 31895 6409 31904 6443
rect 31852 6400 31904 6409
rect 17040 6332 17092 6384
rect 31576 6332 31628 6384
rect 4436 6264 4488 6316
rect 8576 6264 8628 6316
rect 5908 6196 5960 6248
rect 13360 6196 13412 6248
rect 14464 6196 14516 6248
rect 30380 6264 30432 6316
rect 31484 6264 31536 6316
rect 18788 6128 18840 6180
rect 22836 6196 22888 6248
rect 25136 6128 25188 6180
rect 9588 6060 9640 6112
rect 17776 6060 17828 6112
rect 20904 6060 20956 6112
rect 31484 6103 31536 6112
rect 31484 6069 31493 6103
rect 31493 6069 31527 6103
rect 31527 6069 31536 6103
rect 31484 6060 31536 6069
rect 31852 6060 31904 6112
rect 1950 5958 2002 6010
rect 2014 5958 2066 6010
rect 2078 5958 2130 6010
rect 2142 5958 2194 6010
rect 2206 5958 2258 6010
rect 7950 5958 8002 6010
rect 8014 5958 8066 6010
rect 8078 5958 8130 6010
rect 8142 5958 8194 6010
rect 8206 5958 8258 6010
rect 13950 5958 14002 6010
rect 14014 5958 14066 6010
rect 14078 5958 14130 6010
rect 14142 5958 14194 6010
rect 14206 5958 14258 6010
rect 19950 5958 20002 6010
rect 20014 5958 20066 6010
rect 20078 5958 20130 6010
rect 20142 5958 20194 6010
rect 20206 5958 20258 6010
rect 25950 5958 26002 6010
rect 26014 5958 26066 6010
rect 26078 5958 26130 6010
rect 26142 5958 26194 6010
rect 26206 5958 26258 6010
rect 31950 5958 32002 6010
rect 32014 5958 32066 6010
rect 32078 5958 32130 6010
rect 32142 5958 32194 6010
rect 32206 5958 32258 6010
rect 12072 5856 12124 5908
rect 31208 5856 31260 5908
rect 15384 5788 15436 5840
rect 13084 5720 13136 5772
rect 30472 5788 30524 5840
rect 32036 5788 32088 5840
rect 32128 5831 32180 5840
rect 32128 5797 32137 5831
rect 32137 5797 32171 5831
rect 32171 5797 32180 5831
rect 32128 5788 32180 5797
rect 5540 5652 5592 5704
rect 8852 5652 8904 5704
rect 16764 5584 16816 5636
rect 20536 5584 20588 5636
rect 7380 5516 7432 5568
rect 8392 5516 8444 5568
rect 17960 5516 18012 5568
rect 18052 5559 18104 5568
rect 18052 5525 18061 5559
rect 18061 5525 18095 5559
rect 18095 5525 18104 5559
rect 18052 5516 18104 5525
rect 19800 5516 19852 5568
rect 20352 5516 20404 5568
rect 26056 5516 26108 5568
rect 29276 5652 29328 5704
rect 29552 5652 29604 5704
rect 31208 5695 31260 5704
rect 31208 5661 31217 5695
rect 31217 5661 31251 5695
rect 31251 5661 31260 5695
rect 31208 5652 31260 5661
rect 26792 5516 26844 5568
rect 31668 5516 31720 5568
rect 31760 5559 31812 5568
rect 31760 5525 31769 5559
rect 31769 5525 31803 5559
rect 31803 5525 31812 5559
rect 31760 5516 31812 5525
rect 3010 5414 3062 5466
rect 3074 5414 3126 5466
rect 3138 5414 3190 5466
rect 3202 5414 3254 5466
rect 3266 5414 3318 5466
rect 9010 5414 9062 5466
rect 9074 5414 9126 5466
rect 9138 5414 9190 5466
rect 9202 5414 9254 5466
rect 9266 5414 9318 5466
rect 15010 5414 15062 5466
rect 15074 5414 15126 5466
rect 15138 5414 15190 5466
rect 15202 5414 15254 5466
rect 15266 5414 15318 5466
rect 21010 5414 21062 5466
rect 21074 5414 21126 5466
rect 21138 5414 21190 5466
rect 21202 5414 21254 5466
rect 21266 5414 21318 5466
rect 27010 5414 27062 5466
rect 27074 5414 27126 5466
rect 27138 5414 27190 5466
rect 27202 5414 27254 5466
rect 27266 5414 27318 5466
rect 12532 5312 12584 5364
rect 18052 5312 18104 5364
rect 23388 5312 23440 5364
rect 29000 5312 29052 5364
rect 19432 5244 19484 5296
rect 4160 5176 4212 5228
rect 4988 5108 5040 5160
rect 26516 5176 26568 5228
rect 29092 5176 29144 5228
rect 26240 5108 26292 5160
rect 27344 5108 27396 5160
rect 27620 5108 27672 5160
rect 9496 4972 9548 5024
rect 13636 4972 13688 5024
rect 15476 4972 15528 5024
rect 19432 4972 19484 5024
rect 23020 4972 23072 5024
rect 23480 5015 23532 5024
rect 23480 4981 23489 5015
rect 23489 4981 23523 5015
rect 23523 4981 23532 5015
rect 23480 4972 23532 4981
rect 31484 5015 31536 5024
rect 31484 4981 31493 5015
rect 31493 4981 31527 5015
rect 31527 4981 31536 5015
rect 31484 4972 31536 4981
rect 32864 4972 32916 5024
rect 1950 4870 2002 4922
rect 2014 4870 2066 4922
rect 2078 4870 2130 4922
rect 2142 4870 2194 4922
rect 2206 4870 2258 4922
rect 7950 4870 8002 4922
rect 8014 4870 8066 4922
rect 8078 4870 8130 4922
rect 8142 4870 8194 4922
rect 8206 4870 8258 4922
rect 13950 4870 14002 4922
rect 14014 4870 14066 4922
rect 14078 4870 14130 4922
rect 14142 4870 14194 4922
rect 14206 4870 14258 4922
rect 19950 4870 20002 4922
rect 20014 4870 20066 4922
rect 20078 4870 20130 4922
rect 20142 4870 20194 4922
rect 20206 4870 20258 4922
rect 25950 4870 26002 4922
rect 26014 4870 26066 4922
rect 26078 4870 26130 4922
rect 26142 4870 26194 4922
rect 26206 4870 26258 4922
rect 31950 4870 32002 4922
rect 32014 4870 32066 4922
rect 32078 4870 32130 4922
rect 32142 4870 32194 4922
rect 32206 4870 32258 4922
rect 14924 4768 14976 4820
rect 25044 4811 25096 4820
rect 25044 4777 25053 4811
rect 25053 4777 25087 4811
rect 25087 4777 25096 4811
rect 25044 4768 25096 4777
rect 12808 4700 12860 4752
rect 15384 4700 15436 4752
rect 11888 4632 11940 4684
rect 5264 4564 5316 4616
rect 6644 4564 6696 4616
rect 23480 4632 23532 4684
rect 6920 4496 6972 4548
rect 7104 4428 7156 4480
rect 7196 4428 7248 4480
rect 13084 4428 13136 4480
rect 31852 4564 31904 4616
rect 20352 4428 20404 4480
rect 28724 4496 28776 4548
rect 31300 4428 31352 4480
rect 31760 4471 31812 4480
rect 31760 4437 31769 4471
rect 31769 4437 31803 4471
rect 31803 4437 31812 4471
rect 31760 4428 31812 4437
rect 32128 4471 32180 4480
rect 32128 4437 32137 4471
rect 32137 4437 32171 4471
rect 32171 4437 32180 4471
rect 32128 4428 32180 4437
rect 3010 4326 3062 4378
rect 3074 4326 3126 4378
rect 3138 4326 3190 4378
rect 3202 4326 3254 4378
rect 3266 4326 3318 4378
rect 9010 4326 9062 4378
rect 9074 4326 9126 4378
rect 9138 4326 9190 4378
rect 9202 4326 9254 4378
rect 9266 4326 9318 4378
rect 15010 4326 15062 4378
rect 15074 4326 15126 4378
rect 15138 4326 15190 4378
rect 15202 4326 15254 4378
rect 15266 4326 15318 4378
rect 21010 4326 21062 4378
rect 21074 4326 21126 4378
rect 21138 4326 21190 4378
rect 21202 4326 21254 4378
rect 21266 4326 21318 4378
rect 27010 4326 27062 4378
rect 27074 4326 27126 4378
rect 27138 4326 27190 4378
rect 27202 4326 27254 4378
rect 27266 4326 27318 4378
rect 7104 4224 7156 4276
rect 10140 4224 10192 4276
rect 12440 4131 12492 4140
rect 12440 4097 12449 4131
rect 12449 4097 12483 4131
rect 12483 4097 12492 4131
rect 12440 4088 12492 4097
rect 12992 4088 13044 4140
rect 12900 4020 12952 4072
rect 12716 3952 12768 4004
rect 13544 4131 13596 4140
rect 13544 4097 13553 4131
rect 13553 4097 13587 4131
rect 13587 4097 13596 4131
rect 13544 4088 13596 4097
rect 13912 4088 13964 4140
rect 14464 4131 14516 4140
rect 14464 4097 14473 4131
rect 14473 4097 14507 4131
rect 14507 4097 14516 4131
rect 14464 4088 14516 4097
rect 14556 4088 14608 4140
rect 14832 4088 14884 4140
rect 15200 4088 15252 4140
rect 16672 4131 16724 4140
rect 16672 4097 16681 4131
rect 16681 4097 16715 4131
rect 16715 4097 16724 4131
rect 16672 4088 16724 4097
rect 17132 4131 17184 4140
rect 17132 4097 17141 4131
rect 17141 4097 17175 4131
rect 17175 4097 17184 4131
rect 17132 4088 17184 4097
rect 18052 4131 18104 4140
rect 18052 4097 18061 4131
rect 18061 4097 18095 4131
rect 18095 4097 18104 4131
rect 18052 4088 18104 4097
rect 12348 3927 12400 3936
rect 12348 3893 12357 3927
rect 12357 3893 12391 3927
rect 12391 3893 12400 3927
rect 12348 3884 12400 3893
rect 12624 3927 12676 3936
rect 12624 3893 12633 3927
rect 12633 3893 12667 3927
rect 12667 3893 12676 3927
rect 12624 3884 12676 3893
rect 18512 3952 18564 4004
rect 13728 3927 13780 3936
rect 13728 3893 13737 3927
rect 13737 3893 13771 3927
rect 13771 3893 13780 3927
rect 13728 3884 13780 3893
rect 14280 3884 14332 3936
rect 14372 3927 14424 3936
rect 14372 3893 14381 3927
rect 14381 3893 14415 3927
rect 14415 3893 14424 3927
rect 14372 3884 14424 3893
rect 14648 3927 14700 3936
rect 14648 3893 14657 3927
rect 14657 3893 14691 3927
rect 14691 3893 14700 3927
rect 14648 3884 14700 3893
rect 15292 3927 15344 3936
rect 15292 3893 15301 3927
rect 15301 3893 15335 3927
rect 15335 3893 15344 3927
rect 15292 3884 15344 3893
rect 15936 3927 15988 3936
rect 15936 3893 15945 3927
rect 15945 3893 15979 3927
rect 15979 3893 15988 3927
rect 15936 3884 15988 3893
rect 16856 3927 16908 3936
rect 16856 3893 16865 3927
rect 16865 3893 16899 3927
rect 16899 3893 16908 3927
rect 16856 3884 16908 3893
rect 17316 3927 17368 3936
rect 17316 3893 17325 3927
rect 17325 3893 17359 3927
rect 17359 3893 17368 3927
rect 17316 3884 17368 3893
rect 17408 3927 17460 3936
rect 17408 3893 17417 3927
rect 17417 3893 17451 3927
rect 17451 3893 17460 3927
rect 17408 3884 17460 3893
rect 18696 3884 18748 3936
rect 18972 4063 19024 4072
rect 18972 4029 18981 4063
rect 18981 4029 19015 4063
rect 19015 4029 19024 4063
rect 18972 4020 19024 4029
rect 22008 4088 22060 4140
rect 22376 4131 22428 4140
rect 22376 4097 22385 4131
rect 22385 4097 22419 4131
rect 22419 4097 22428 4131
rect 22376 4088 22428 4097
rect 23296 4131 23348 4140
rect 23296 4097 23305 4131
rect 23305 4097 23339 4131
rect 23339 4097 23348 4131
rect 23296 4088 23348 4097
rect 28448 4088 28500 4140
rect 31300 4131 31352 4140
rect 31300 4097 31309 4131
rect 31309 4097 31343 4131
rect 31343 4097 31352 4131
rect 31300 4088 31352 4097
rect 18880 3952 18932 4004
rect 28172 4020 28224 4072
rect 29000 4020 29052 4072
rect 20904 3952 20956 4004
rect 22192 3995 22244 4004
rect 22192 3961 22201 3995
rect 22201 3961 22235 3995
rect 22235 3961 22244 3995
rect 22192 3952 22244 3961
rect 23112 3995 23164 4004
rect 23112 3961 23121 3995
rect 23121 3961 23155 3995
rect 23155 3961 23164 3995
rect 23112 3952 23164 3961
rect 23664 3995 23716 4004
rect 23664 3961 23673 3995
rect 23673 3961 23707 3995
rect 23707 3961 23716 3995
rect 23664 3952 23716 3961
rect 26424 3952 26476 4004
rect 19800 3884 19852 3936
rect 31300 3884 31352 3936
rect 31484 3927 31536 3936
rect 31484 3893 31493 3927
rect 31493 3893 31527 3927
rect 31527 3893 31536 3927
rect 31484 3884 31536 3893
rect 32864 3884 32916 3936
rect 1950 3782 2002 3834
rect 2014 3782 2066 3834
rect 2078 3782 2130 3834
rect 2142 3782 2194 3834
rect 2206 3782 2258 3834
rect 7950 3782 8002 3834
rect 8014 3782 8066 3834
rect 8078 3782 8130 3834
rect 8142 3782 8194 3834
rect 8206 3782 8258 3834
rect 13950 3782 14002 3834
rect 14014 3782 14066 3834
rect 14078 3782 14130 3834
rect 14142 3782 14194 3834
rect 14206 3782 14258 3834
rect 19950 3782 20002 3834
rect 20014 3782 20066 3834
rect 20078 3782 20130 3834
rect 20142 3782 20194 3834
rect 20206 3782 20258 3834
rect 25950 3782 26002 3834
rect 26014 3782 26066 3834
rect 26078 3782 26130 3834
rect 26142 3782 26194 3834
rect 26206 3782 26258 3834
rect 31950 3782 32002 3834
rect 32014 3782 32066 3834
rect 32078 3782 32130 3834
rect 32142 3782 32194 3834
rect 32206 3782 32258 3834
rect 9404 3680 9456 3732
rect 13544 3680 13596 3732
rect 13728 3680 13780 3732
rect 15476 3680 15528 3732
rect 15936 3680 15988 3732
rect 17224 3680 17276 3732
rect 17316 3680 17368 3732
rect 22744 3680 22796 3732
rect 23296 3680 23348 3732
rect 27896 3680 27948 3732
rect 12624 3612 12676 3664
rect 19892 3612 19944 3664
rect 12164 3544 12216 3596
rect 13728 3544 13780 3596
rect 14280 3544 14332 3596
rect 17500 3544 17552 3596
rect 21456 3612 21508 3664
rect 24124 3612 24176 3664
rect 13820 3476 13872 3528
rect 14188 3476 14240 3528
rect 15108 3476 15160 3528
rect 15292 3476 15344 3528
rect 19340 3476 19392 3528
rect 12532 3408 12584 3460
rect 14464 3408 14516 3460
rect 14648 3408 14700 3460
rect 17868 3408 17920 3460
rect 19524 3408 19576 3460
rect 15936 3340 15988 3392
rect 17224 3340 17276 3392
rect 19156 3340 19208 3392
rect 22284 3544 22336 3596
rect 22376 3544 22428 3596
rect 27620 3544 27672 3596
rect 20720 3476 20772 3528
rect 21732 3519 21784 3528
rect 21732 3485 21741 3519
rect 21741 3485 21775 3519
rect 21775 3485 21784 3519
rect 21732 3476 21784 3485
rect 20352 3408 20404 3460
rect 21364 3408 21416 3460
rect 20260 3383 20312 3392
rect 20260 3349 20269 3383
rect 20269 3349 20303 3383
rect 20303 3349 20312 3383
rect 20260 3340 20312 3349
rect 20444 3383 20496 3392
rect 20444 3349 20453 3383
rect 20453 3349 20487 3383
rect 20487 3349 20496 3383
rect 20444 3340 20496 3349
rect 20812 3383 20864 3392
rect 20812 3349 20821 3383
rect 20821 3349 20855 3383
rect 20855 3349 20864 3383
rect 20812 3340 20864 3349
rect 23940 3408 23992 3460
rect 25228 3451 25280 3460
rect 25228 3417 25237 3451
rect 25237 3417 25271 3451
rect 25271 3417 25280 3451
rect 25228 3408 25280 3417
rect 25780 3383 25832 3392
rect 25780 3349 25789 3383
rect 25789 3349 25823 3383
rect 25823 3349 25832 3383
rect 25780 3340 25832 3349
rect 26240 3383 26292 3392
rect 26240 3349 26249 3383
rect 26249 3349 26283 3383
rect 26283 3349 26292 3383
rect 26240 3340 26292 3349
rect 31668 3340 31720 3392
rect 31760 3383 31812 3392
rect 31760 3349 31769 3383
rect 31769 3349 31803 3383
rect 31803 3349 31812 3383
rect 31760 3340 31812 3349
rect 32128 3383 32180 3392
rect 32128 3349 32137 3383
rect 32137 3349 32171 3383
rect 32171 3349 32180 3383
rect 32128 3340 32180 3349
rect 3010 3238 3062 3290
rect 3074 3238 3126 3290
rect 3138 3238 3190 3290
rect 3202 3238 3254 3290
rect 3266 3238 3318 3290
rect 9010 3238 9062 3290
rect 9074 3238 9126 3290
rect 9138 3238 9190 3290
rect 9202 3238 9254 3290
rect 9266 3238 9318 3290
rect 15010 3238 15062 3290
rect 15074 3238 15126 3290
rect 15138 3238 15190 3290
rect 15202 3238 15254 3290
rect 15266 3238 15318 3290
rect 21010 3238 21062 3290
rect 21074 3238 21126 3290
rect 21138 3238 21190 3290
rect 21202 3238 21254 3290
rect 21266 3238 21318 3290
rect 27010 3238 27062 3290
rect 27074 3238 27126 3290
rect 27138 3238 27190 3290
rect 27202 3238 27254 3290
rect 27266 3238 27318 3290
rect 14372 3136 14424 3188
rect 20628 3136 20680 3188
rect 20812 3136 20864 3188
rect 30932 3136 30984 3188
rect 11612 3068 11664 3120
rect 14832 3068 14884 3120
rect 18512 3068 18564 3120
rect 14740 3000 14792 3052
rect 15384 3000 15436 3052
rect 16120 3043 16172 3052
rect 16120 3009 16129 3043
rect 16129 3009 16163 3043
rect 16163 3009 16172 3043
rect 16120 3000 16172 3009
rect 19432 3043 19484 3052
rect 19432 3009 19441 3043
rect 19441 3009 19475 3043
rect 19475 3009 19484 3043
rect 19432 3000 19484 3009
rect 20260 3068 20312 3120
rect 20904 3043 20956 3052
rect 20904 3009 20913 3043
rect 20913 3009 20947 3043
rect 20947 3009 20956 3043
rect 20904 3000 20956 3009
rect 21364 3000 21416 3052
rect 22744 3043 22796 3052
rect 22744 3009 22753 3043
rect 22753 3009 22787 3043
rect 22787 3009 22796 3043
rect 22744 3000 22796 3009
rect 12348 2932 12400 2984
rect 19708 2932 19760 2984
rect 19800 2932 19852 2984
rect 31300 3043 31352 3052
rect 31300 3009 31309 3043
rect 31309 3009 31343 3043
rect 31343 3009 31352 3043
rect 31300 3000 31352 3009
rect 31668 3043 31720 3052
rect 31668 3009 31677 3043
rect 31677 3009 31711 3043
rect 31711 3009 31720 3043
rect 31668 3000 31720 3009
rect 12900 2864 12952 2916
rect 13544 2864 13596 2916
rect 16856 2864 16908 2916
rect 19892 2864 19944 2916
rect 20536 2864 20588 2916
rect 21456 2864 21508 2916
rect 22376 2864 22428 2916
rect 12440 2796 12492 2848
rect 13268 2796 13320 2848
rect 14372 2796 14424 2848
rect 15384 2796 15436 2848
rect 16028 2796 16080 2848
rect 17776 2796 17828 2848
rect 18512 2796 18564 2848
rect 19340 2796 19392 2848
rect 19800 2796 19852 2848
rect 20444 2796 20496 2848
rect 20812 2796 20864 2848
rect 21548 2796 21600 2848
rect 22652 2796 22704 2848
rect 23204 2796 23256 2848
rect 23756 2796 23808 2848
rect 31760 2796 31812 2848
rect 32864 2796 32916 2848
rect 1950 2694 2002 2746
rect 2014 2694 2066 2746
rect 2078 2694 2130 2746
rect 2142 2694 2194 2746
rect 2206 2694 2258 2746
rect 7950 2694 8002 2746
rect 8014 2694 8066 2746
rect 8078 2694 8130 2746
rect 8142 2694 8194 2746
rect 8206 2694 8258 2746
rect 13950 2694 14002 2746
rect 14014 2694 14066 2746
rect 14078 2694 14130 2746
rect 14142 2694 14194 2746
rect 14206 2694 14258 2746
rect 19950 2694 20002 2746
rect 20014 2694 20066 2746
rect 20078 2694 20130 2746
rect 20142 2694 20194 2746
rect 20206 2694 20258 2746
rect 25950 2694 26002 2746
rect 26014 2694 26066 2746
rect 26078 2694 26130 2746
rect 26142 2694 26194 2746
rect 26206 2694 26258 2746
rect 31950 2694 32002 2746
rect 32014 2694 32066 2746
rect 32078 2694 32130 2746
rect 32142 2694 32194 2746
rect 32206 2694 32258 2746
rect 9496 2592 9548 2644
rect 14188 2592 14240 2644
rect 17684 2592 17736 2644
rect 18880 2592 18932 2644
rect 19524 2592 19576 2644
rect 13176 2524 13228 2576
rect 9588 2456 9640 2508
rect 15476 2524 15528 2576
rect 18236 2524 18288 2576
rect 19064 2524 19116 2576
rect 19432 2524 19484 2576
rect 13636 2431 13688 2440
rect 13636 2397 13645 2431
rect 13645 2397 13679 2431
rect 13679 2397 13688 2431
rect 13636 2388 13688 2397
rect 14464 2388 14516 2440
rect 14924 2388 14976 2440
rect 12808 2320 12860 2372
rect 16212 2431 16264 2440
rect 16212 2397 16221 2431
rect 16221 2397 16255 2431
rect 16255 2397 16264 2431
rect 16212 2388 16264 2397
rect 16764 2431 16816 2440
rect 16764 2397 16773 2431
rect 16773 2397 16807 2431
rect 16807 2397 16816 2431
rect 16764 2388 16816 2397
rect 16948 2388 17000 2440
rect 17500 2431 17552 2440
rect 17500 2397 17509 2431
rect 17509 2397 17543 2431
rect 17543 2397 17552 2431
rect 17500 2388 17552 2397
rect 17960 2388 18012 2440
rect 18512 2388 18564 2440
rect 15568 2320 15620 2372
rect 19432 2388 19484 2440
rect 21456 2592 21508 2644
rect 22468 2592 22520 2644
rect 19892 2524 19944 2576
rect 21824 2524 21876 2576
rect 22928 2524 22980 2576
rect 24124 2524 24176 2576
rect 20536 2456 20588 2508
rect 19984 2431 20036 2440
rect 19984 2397 19993 2431
rect 19993 2397 20027 2431
rect 20027 2397 20036 2431
rect 19984 2388 20036 2397
rect 20352 2431 20404 2440
rect 20352 2397 20361 2431
rect 20361 2397 20395 2431
rect 20395 2397 20404 2431
rect 20352 2388 20404 2397
rect 22284 2456 22336 2508
rect 21640 2388 21692 2440
rect 20536 2320 20588 2372
rect 20628 2320 20680 2372
rect 22376 2388 22428 2440
rect 22744 2388 22796 2440
rect 23296 2431 23348 2440
rect 23296 2397 23305 2431
rect 23305 2397 23339 2431
rect 23339 2397 23348 2431
rect 23296 2388 23348 2397
rect 23664 2431 23716 2440
rect 23664 2397 23673 2431
rect 23673 2397 23707 2431
rect 23707 2397 23716 2431
rect 23664 2388 23716 2397
rect 23940 2456 23992 2508
rect 30932 2431 30984 2440
rect 30932 2397 30941 2431
rect 30941 2397 30975 2431
rect 30975 2397 30984 2431
rect 30932 2388 30984 2397
rect 31300 2431 31352 2440
rect 31300 2397 31309 2431
rect 31309 2397 31343 2431
rect 31343 2397 31352 2431
rect 31300 2388 31352 2397
rect 14096 2252 14148 2304
rect 14188 2252 14240 2304
rect 14464 2252 14516 2304
rect 14648 2252 14700 2304
rect 14924 2295 14976 2304
rect 14924 2261 14933 2295
rect 14933 2261 14967 2295
rect 14967 2261 14976 2295
rect 14924 2252 14976 2261
rect 15476 2252 15528 2304
rect 15752 2252 15804 2304
rect 16304 2252 16356 2304
rect 16580 2252 16632 2304
rect 16856 2252 16908 2304
rect 17132 2252 17184 2304
rect 17408 2252 17460 2304
rect 17960 2252 18012 2304
rect 18512 2252 18564 2304
rect 19616 2252 19668 2304
rect 19708 2252 19760 2304
rect 20168 2295 20220 2304
rect 20168 2261 20177 2295
rect 20177 2261 20211 2295
rect 20211 2261 20220 2295
rect 20168 2252 20220 2261
rect 20260 2252 20312 2304
rect 21364 2252 21416 2304
rect 22100 2252 22152 2304
rect 23572 2252 23624 2304
rect 30748 2295 30800 2304
rect 30748 2261 30757 2295
rect 30757 2261 30791 2295
rect 30791 2261 30800 2295
rect 30748 2252 30800 2261
rect 31116 2295 31168 2304
rect 31116 2261 31125 2295
rect 31125 2261 31159 2295
rect 31159 2261 31168 2295
rect 31116 2252 31168 2261
rect 31484 2295 31536 2304
rect 31484 2261 31493 2295
rect 31493 2261 31527 2295
rect 31527 2261 31536 2295
rect 31484 2252 31536 2261
rect 31852 2295 31904 2304
rect 31852 2261 31861 2295
rect 31861 2261 31895 2295
rect 31895 2261 31904 2295
rect 31852 2252 31904 2261
rect 3010 2150 3062 2202
rect 3074 2150 3126 2202
rect 3138 2150 3190 2202
rect 3202 2150 3254 2202
rect 3266 2150 3318 2202
rect 9010 2150 9062 2202
rect 9074 2150 9126 2202
rect 9138 2150 9190 2202
rect 9202 2150 9254 2202
rect 9266 2150 9318 2202
rect 15010 2150 15062 2202
rect 15074 2150 15126 2202
rect 15138 2150 15190 2202
rect 15202 2150 15254 2202
rect 15266 2150 15318 2202
rect 21010 2150 21062 2202
rect 21074 2150 21126 2202
rect 21138 2150 21190 2202
rect 21202 2150 21254 2202
rect 21266 2150 21318 2202
rect 27010 2150 27062 2202
rect 27074 2150 27126 2202
rect 27138 2150 27190 2202
rect 27202 2150 27254 2202
rect 27266 2150 27318 2202
rect 11336 2048 11388 2100
rect 14280 2048 14332 2100
rect 17868 2048 17920 2100
rect 21640 2048 21692 2100
rect 22008 2048 22060 2100
rect 23664 2048 23716 2100
rect 9680 1980 9732 2032
rect 6184 1912 6236 1964
rect 18880 1980 18932 2032
rect 18972 1980 19024 2032
rect 19708 1980 19760 2032
rect 19800 1980 19852 2032
rect 23296 1980 23348 2032
rect 15936 1912 15988 1964
rect 20352 1912 20404 1964
rect 19984 1844 20036 1896
rect 8392 1776 8444 1828
rect 19432 1776 19484 1828
rect 9956 1708 10008 1760
rect 19064 1708 19116 1760
rect 19156 1708 19208 1760
rect 22744 1844 22796 1896
rect 10140 1640 10192 1692
rect 16948 1640 17000 1692
rect 18696 1640 18748 1692
rect 31300 1640 31352 1692
rect 13360 1572 13412 1624
rect 16212 1572 16264 1624
rect 19064 1368 19116 1420
rect 20168 1368 20220 1420
rect 9496 1300 9548 1352
rect 14556 1300 14608 1352
rect 19524 1300 19576 1352
rect 25412 1300 25464 1352
rect 11060 1232 11112 1284
rect 16672 1232 16724 1284
rect 22836 1096 22888 1148
rect 27068 1096 27120 1148
<< metal2 >>
rect 1214 11194 1270 11250
rect 2778 11194 2834 11250
rect 4342 11194 4398 11250
rect 5906 11194 5962 11250
rect 7470 11194 7526 11250
rect 9034 11194 9090 11250
rect 10598 11194 10654 11250
rect 12162 11194 12218 11250
rect 13726 11194 13782 11250
rect 15290 11194 15346 11250
rect 16854 11194 16910 11250
rect 18418 11194 18474 11250
rect 19982 11194 20038 11250
rect 21546 11194 21602 11250
rect 23110 11194 23166 11250
rect 24674 11194 24730 11250
rect 26238 11194 26294 11250
rect 27802 11194 27858 11250
rect 29366 11194 29422 11250
rect 30930 11194 30986 11250
rect 32494 11194 32550 11250
rect 1228 8634 1256 11194
rect 2792 8634 2820 11194
rect 3010 8732 3318 8741
rect 3010 8730 3016 8732
rect 3072 8730 3096 8732
rect 3152 8730 3176 8732
rect 3232 8730 3256 8732
rect 3312 8730 3318 8732
rect 3072 8678 3074 8730
rect 3254 8678 3256 8730
rect 3010 8676 3016 8678
rect 3072 8676 3096 8678
rect 3152 8676 3176 8678
rect 3232 8676 3256 8678
rect 3312 8676 3318 8678
rect 2870 8664 2926 8673
rect 3010 8667 3318 8676
rect 1216 8628 1268 8634
rect 1216 8570 1268 8576
rect 2780 8628 2832 8634
rect 4356 8634 4384 11194
rect 4802 9344 4858 9353
rect 4802 9279 4858 9288
rect 4712 8832 4764 8838
rect 4712 8774 4764 8780
rect 4724 8634 4752 8774
rect 2870 8599 2926 8608
rect 4344 8628 4396 8634
rect 2780 8570 2832 8576
rect 1582 8528 1638 8537
rect 1582 8463 1584 8472
rect 1636 8463 1638 8472
rect 1584 8434 1636 8440
rect 2884 8401 2912 8599
rect 4344 8570 4396 8576
rect 4712 8628 4764 8634
rect 4712 8570 4764 8576
rect 2870 8392 2926 8401
rect 2870 8327 2926 8336
rect 1950 8188 2258 8197
rect 1950 8186 1956 8188
rect 2012 8186 2036 8188
rect 2092 8186 2116 8188
rect 2172 8186 2196 8188
rect 2252 8186 2258 8188
rect 2012 8134 2014 8186
rect 2194 8134 2196 8186
rect 1950 8132 1956 8134
rect 2012 8132 2036 8134
rect 2092 8132 2116 8134
rect 2172 8132 2196 8134
rect 2252 8132 2258 8134
rect 1950 8123 2258 8132
rect 3010 7644 3318 7653
rect 3010 7642 3016 7644
rect 3072 7642 3096 7644
rect 3152 7642 3176 7644
rect 3232 7642 3256 7644
rect 3312 7642 3318 7644
rect 3072 7590 3074 7642
rect 3254 7590 3256 7642
rect 3010 7588 3016 7590
rect 3072 7588 3096 7590
rect 3152 7588 3176 7590
rect 3232 7588 3256 7590
rect 3312 7588 3318 7590
rect 3010 7579 3318 7588
rect 4816 7410 4844 9279
rect 4988 8968 5040 8974
rect 4988 8910 5040 8916
rect 5000 8430 5028 8910
rect 5920 8634 5948 11194
rect 7378 8936 7434 8945
rect 7378 8871 7434 8880
rect 5908 8628 5960 8634
rect 5908 8570 5960 8576
rect 4988 8424 5040 8430
rect 4988 8366 5040 8372
rect 4896 8016 4948 8022
rect 4896 7958 4948 7964
rect 7012 8016 7064 8022
rect 7012 7958 7064 7964
rect 4908 7546 4936 7958
rect 6826 7848 6882 7857
rect 6826 7783 6882 7792
rect 5632 7744 5684 7750
rect 5632 7686 5684 7692
rect 4896 7540 4948 7546
rect 4896 7482 4948 7488
rect 5540 7472 5592 7478
rect 5540 7414 5592 7420
rect 4712 7404 4764 7410
rect 4712 7346 4764 7352
rect 4804 7404 4856 7410
rect 4804 7346 4856 7352
rect 1950 7100 2258 7109
rect 1950 7098 1956 7100
rect 2012 7098 2036 7100
rect 2092 7098 2116 7100
rect 2172 7098 2196 7100
rect 2252 7098 2258 7100
rect 2012 7046 2014 7098
rect 2194 7046 2196 7098
rect 1950 7044 1956 7046
rect 2012 7044 2036 7046
rect 2092 7044 2116 7046
rect 2172 7044 2196 7046
rect 2252 7044 2258 7046
rect 1950 7035 2258 7044
rect 4724 7002 4752 7346
rect 5552 7313 5580 7414
rect 5538 7304 5594 7313
rect 5538 7239 5594 7248
rect 4712 6996 4764 7002
rect 4712 6938 4764 6944
rect 5644 6914 5672 7686
rect 6092 7540 6144 7546
rect 6092 7482 6144 7488
rect 5906 7304 5962 7313
rect 5906 7239 5908 7248
rect 5960 7239 5962 7248
rect 5908 7210 5960 7216
rect 5552 6886 5672 6914
rect 4712 6724 4764 6730
rect 4712 6666 4764 6672
rect 3010 6556 3318 6565
rect 3010 6554 3016 6556
rect 3072 6554 3096 6556
rect 3152 6554 3176 6556
rect 3232 6554 3256 6556
rect 3312 6554 3318 6556
rect 3072 6502 3074 6554
rect 3254 6502 3256 6554
rect 3010 6500 3016 6502
rect 3072 6500 3096 6502
rect 3152 6500 3176 6502
rect 3232 6500 3256 6502
rect 3312 6500 3318 6502
rect 3010 6491 3318 6500
rect 4436 6316 4488 6322
rect 4436 6258 4488 6264
rect 1950 6012 2258 6021
rect 1950 6010 1956 6012
rect 2012 6010 2036 6012
rect 2092 6010 2116 6012
rect 2172 6010 2196 6012
rect 2252 6010 2258 6012
rect 2012 5958 2014 6010
rect 2194 5958 2196 6010
rect 1950 5956 1956 5958
rect 2012 5956 2036 5958
rect 2092 5956 2116 5958
rect 2172 5956 2196 5958
rect 2252 5956 2258 5958
rect 1950 5947 2258 5956
rect 3010 5468 3318 5477
rect 3010 5466 3016 5468
rect 3072 5466 3096 5468
rect 3152 5466 3176 5468
rect 3232 5466 3256 5468
rect 3312 5466 3318 5468
rect 3072 5414 3074 5466
rect 3254 5414 3256 5466
rect 3010 5412 3016 5414
rect 3072 5412 3096 5414
rect 3152 5412 3176 5414
rect 3232 5412 3256 5414
rect 3312 5412 3318 5414
rect 3010 5403 3318 5412
rect 4160 5228 4212 5234
rect 4160 5170 4212 5176
rect 1950 4924 2258 4933
rect 1950 4922 1956 4924
rect 2012 4922 2036 4924
rect 2092 4922 2116 4924
rect 2172 4922 2196 4924
rect 2252 4922 2258 4924
rect 2012 4870 2014 4922
rect 2194 4870 2196 4922
rect 1950 4868 1956 4870
rect 2012 4868 2036 4870
rect 2092 4868 2116 4870
rect 2172 4868 2196 4870
rect 2252 4868 2258 4870
rect 1950 4859 2258 4868
rect 3010 4380 3318 4389
rect 3010 4378 3016 4380
rect 3072 4378 3096 4380
rect 3152 4378 3176 4380
rect 3232 4378 3256 4380
rect 3312 4378 3318 4380
rect 3072 4326 3074 4378
rect 3254 4326 3256 4378
rect 3010 4324 3016 4326
rect 3072 4324 3096 4326
rect 3152 4324 3176 4326
rect 3232 4324 3256 4326
rect 3312 4324 3318 4326
rect 3010 4315 3318 4324
rect 1950 3836 2258 3845
rect 1950 3834 1956 3836
rect 2012 3834 2036 3836
rect 2092 3834 2116 3836
rect 2172 3834 2196 3836
rect 2252 3834 2258 3836
rect 2012 3782 2014 3834
rect 2194 3782 2196 3834
rect 1950 3780 1956 3782
rect 2012 3780 2036 3782
rect 2092 3780 2116 3782
rect 2172 3780 2196 3782
rect 2252 3780 2258 3782
rect 1950 3771 2258 3780
rect 3010 3292 3318 3301
rect 3010 3290 3016 3292
rect 3072 3290 3096 3292
rect 3152 3290 3176 3292
rect 3232 3290 3256 3292
rect 3312 3290 3318 3292
rect 3072 3238 3074 3290
rect 3254 3238 3256 3290
rect 3010 3236 3016 3238
rect 3072 3236 3096 3238
rect 3152 3236 3176 3238
rect 3232 3236 3256 3238
rect 3312 3236 3318 3238
rect 3010 3227 3318 3236
rect 1950 2748 2258 2757
rect 1950 2746 1956 2748
rect 2012 2746 2036 2748
rect 2092 2746 2116 2748
rect 2172 2746 2196 2748
rect 2252 2746 2258 2748
rect 2012 2694 2014 2746
rect 2194 2694 2196 2746
rect 1950 2692 1956 2694
rect 2012 2692 2036 2694
rect 2092 2692 2116 2694
rect 2172 2692 2196 2694
rect 2252 2692 2258 2694
rect 1950 2683 2258 2692
rect 2870 2272 2926 2281
rect 2870 2207 2926 2216
rect 2884 1873 2912 2207
rect 3010 2204 3318 2213
rect 3010 2202 3016 2204
rect 3072 2202 3096 2204
rect 3152 2202 3176 2204
rect 3232 2202 3256 2204
rect 3312 2202 3318 2204
rect 3072 2150 3074 2202
rect 3254 2150 3256 2202
rect 3010 2148 3016 2150
rect 3072 2148 3096 2150
rect 3152 2148 3176 2150
rect 3232 2148 3256 2150
rect 3312 2148 3318 2150
rect 3010 2139 3318 2148
rect 2870 1864 2926 1873
rect 2870 1799 2926 1808
rect 4172 56 4200 5170
rect 4448 56 4476 6258
rect 4724 56 4752 6666
rect 5552 6361 5580 6886
rect 5816 6792 5868 6798
rect 5816 6734 5868 6740
rect 5538 6352 5594 6361
rect 5538 6287 5594 6296
rect 5540 5704 5592 5710
rect 5540 5646 5592 5652
rect 4988 5160 5040 5166
rect 4988 5102 5040 5108
rect 5000 56 5028 5102
rect 5264 4616 5316 4622
rect 5264 4558 5316 4564
rect 5276 56 5304 4558
rect 5552 56 5580 5646
rect 5828 56 5856 6734
rect 5908 6656 5960 6662
rect 5908 6598 5960 6604
rect 5920 6254 5948 6598
rect 5908 6248 5960 6254
rect 5908 6190 5960 6196
rect 6104 56 6132 7482
rect 6840 7410 6868 7783
rect 6828 7404 6880 7410
rect 6828 7346 6880 7352
rect 6276 7268 6328 7274
rect 6276 7210 6328 7216
rect 6184 7200 6236 7206
rect 6184 7142 6236 7148
rect 6196 1970 6224 7142
rect 6288 6905 6316 7210
rect 7024 7206 7052 7958
rect 7392 7818 7420 8871
rect 7484 8634 7512 11194
rect 7746 9616 7802 9625
rect 7746 9551 7802 9560
rect 7472 8628 7524 8634
rect 7472 8570 7524 8576
rect 7654 8256 7710 8265
rect 7654 8191 7710 8200
rect 7668 7954 7696 8191
rect 7656 7948 7708 7954
rect 7656 7890 7708 7896
rect 7564 7880 7616 7886
rect 7564 7822 7616 7828
rect 7380 7812 7432 7818
rect 7380 7754 7432 7760
rect 7576 7546 7604 7822
rect 7564 7540 7616 7546
rect 7564 7482 7616 7488
rect 7104 7336 7156 7342
rect 7104 7278 7156 7284
rect 7012 7200 7064 7206
rect 7012 7142 7064 7148
rect 7116 6934 7144 7278
rect 7760 7206 7788 9551
rect 9048 9466 9076 11194
rect 8864 9438 9076 9466
rect 8864 8634 8892 9438
rect 9404 9240 9456 9246
rect 9404 9182 9456 9188
rect 9010 8732 9318 8741
rect 9010 8730 9016 8732
rect 9072 8730 9096 8732
rect 9152 8730 9176 8732
rect 9232 8730 9256 8732
rect 9312 8730 9318 8732
rect 9072 8678 9074 8730
rect 9254 8678 9256 8730
rect 9010 8676 9016 8678
rect 9072 8676 9096 8678
rect 9152 8676 9176 8678
rect 9232 8676 9256 8678
rect 9312 8676 9318 8678
rect 9010 8667 9318 8676
rect 8852 8628 8904 8634
rect 8852 8570 8904 8576
rect 9416 8498 9444 9182
rect 10612 8634 10640 11194
rect 10968 8900 11020 8906
rect 10968 8842 11020 8848
rect 10600 8628 10652 8634
rect 10600 8570 10652 8576
rect 10980 8498 11008 8842
rect 12176 8634 12204 11194
rect 12532 9172 12584 9178
rect 12532 9114 12584 9120
rect 12438 9072 12494 9081
rect 12438 9007 12494 9016
rect 12072 8628 12124 8634
rect 12072 8570 12124 8576
rect 12164 8628 12216 8634
rect 12164 8570 12216 8576
rect 9404 8492 9456 8498
rect 9404 8434 9456 8440
rect 10968 8492 11020 8498
rect 10968 8434 11020 8440
rect 7950 8188 8258 8197
rect 7950 8186 7956 8188
rect 8012 8186 8036 8188
rect 8092 8186 8116 8188
rect 8172 8186 8196 8188
rect 8252 8186 8258 8188
rect 8012 8134 8014 8186
rect 8194 8134 8196 8186
rect 7950 8132 7956 8134
rect 8012 8132 8036 8134
rect 8092 8132 8116 8134
rect 8172 8132 8196 8134
rect 8252 8132 8258 8134
rect 7950 8123 8258 8132
rect 12084 7750 12112 8570
rect 12164 7812 12216 7818
rect 12164 7754 12216 7760
rect 8116 7744 8168 7750
rect 8116 7686 8168 7692
rect 12072 7744 12124 7750
rect 12072 7686 12124 7692
rect 8128 7478 8156 7686
rect 9010 7644 9318 7653
rect 9010 7642 9016 7644
rect 9072 7642 9096 7644
rect 9152 7642 9176 7644
rect 9232 7642 9256 7644
rect 9312 7642 9318 7644
rect 9072 7590 9074 7642
rect 9254 7590 9256 7642
rect 9010 7588 9016 7590
rect 9072 7588 9096 7590
rect 9152 7588 9176 7590
rect 9232 7588 9256 7590
rect 9312 7588 9318 7590
rect 9010 7579 9318 7588
rect 8116 7472 8168 7478
rect 8116 7414 8168 7420
rect 12176 7410 12204 7754
rect 12452 7410 12480 9007
rect 12544 8498 12572 9114
rect 12624 9104 12676 9110
rect 12624 9046 12676 9052
rect 12532 8492 12584 8498
rect 12532 8434 12584 8440
rect 12636 7698 12664 9046
rect 13740 8634 13768 11194
rect 14280 9308 14332 9314
rect 14280 9250 14332 9256
rect 13728 8628 13780 8634
rect 13728 8570 13780 8576
rect 13950 8188 14258 8197
rect 13950 8186 13956 8188
rect 14012 8186 14036 8188
rect 14092 8186 14116 8188
rect 14172 8186 14196 8188
rect 14252 8186 14258 8188
rect 14012 8134 14014 8186
rect 14194 8134 14196 8186
rect 13950 8132 13956 8134
rect 14012 8132 14036 8134
rect 14092 8132 14116 8134
rect 14172 8132 14196 8134
rect 14252 8132 14258 8134
rect 13950 8123 14258 8132
rect 14292 7970 14320 9250
rect 14372 8832 14424 8838
rect 15304 8820 15332 11194
rect 16764 9444 16816 9450
rect 16764 9386 16816 9392
rect 16776 8838 16804 9386
rect 16764 8832 16816 8838
rect 15304 8792 15424 8820
rect 14372 8774 14424 8780
rect 14384 8498 14412 8774
rect 15010 8732 15318 8741
rect 15010 8730 15016 8732
rect 15072 8730 15096 8732
rect 15152 8730 15176 8732
rect 15232 8730 15256 8732
rect 15312 8730 15318 8732
rect 15072 8678 15074 8730
rect 15254 8678 15256 8730
rect 15010 8676 15016 8678
rect 15072 8676 15096 8678
rect 15152 8676 15176 8678
rect 15232 8676 15256 8678
rect 15312 8676 15318 8678
rect 15010 8667 15318 8676
rect 15396 8634 15424 8792
rect 16764 8774 16816 8780
rect 16868 8634 16896 11194
rect 17130 9888 17186 9897
rect 17130 9823 17186 9832
rect 17040 8900 17092 8906
rect 17040 8842 17092 8848
rect 15384 8628 15436 8634
rect 15384 8570 15436 8576
rect 16856 8628 16908 8634
rect 16856 8570 16908 8576
rect 15672 8498 15884 8514
rect 14372 8492 14424 8498
rect 14372 8434 14424 8440
rect 15660 8492 15884 8498
rect 15712 8486 15884 8492
rect 15660 8434 15712 8440
rect 15856 8430 15884 8486
rect 17052 8430 17080 8842
rect 15844 8424 15896 8430
rect 15106 8392 15162 8401
rect 14924 8356 14976 8362
rect 15844 8366 15896 8372
rect 17040 8424 17092 8430
rect 17040 8366 17092 8372
rect 15106 8327 15162 8336
rect 14924 8298 14976 8304
rect 13360 7948 13412 7954
rect 13360 7890 13412 7896
rect 14200 7942 14320 7970
rect 14554 7984 14610 7993
rect 12544 7670 12664 7698
rect 11888 7404 11940 7410
rect 11888 7346 11940 7352
rect 12164 7404 12216 7410
rect 12164 7346 12216 7352
rect 12440 7404 12492 7410
rect 12440 7346 12492 7352
rect 7840 7336 7892 7342
rect 7840 7278 7892 7284
rect 7380 7200 7432 7206
rect 7380 7142 7432 7148
rect 7748 7200 7800 7206
rect 7748 7142 7800 7148
rect 7104 6928 7156 6934
rect 6274 6896 6330 6905
rect 7104 6870 7156 6876
rect 6274 6831 6330 6840
rect 6368 6724 6420 6730
rect 6368 6666 6420 6672
rect 6184 1964 6236 1970
rect 6184 1906 6236 1912
rect 6380 56 6408 6666
rect 7392 5574 7420 7142
rect 7472 6996 7524 7002
rect 7472 6938 7524 6944
rect 7380 5568 7432 5574
rect 7380 5510 7432 5516
rect 6644 4616 6696 4622
rect 6644 4558 6696 4564
rect 6656 56 6684 4558
rect 6920 4548 6972 4554
rect 6920 4490 6972 4496
rect 6932 56 6960 4490
rect 7104 4480 7156 4486
rect 7104 4422 7156 4428
rect 7196 4480 7248 4486
rect 7196 4422 7248 4428
rect 7116 4282 7144 4422
rect 7104 4276 7156 4282
rect 7104 4218 7156 4224
rect 7208 56 7236 4422
rect 7484 56 7512 6938
rect 7748 6928 7800 6934
rect 7748 6870 7800 6876
rect 7760 56 7788 6870
rect 4158 0 4214 56
rect 4434 0 4490 56
rect 4710 0 4766 56
rect 4986 0 5042 56
rect 5262 0 5318 56
rect 5538 0 5594 56
rect 5814 0 5870 56
rect 6090 0 6146 56
rect 6366 0 6422 56
rect 6642 0 6698 56
rect 6918 0 6974 56
rect 7194 0 7250 56
rect 7470 0 7526 56
rect 7746 0 7802 56
rect 7852 42 7880 7278
rect 9312 7268 9364 7274
rect 9312 7210 9364 7216
rect 10968 7268 11020 7274
rect 10968 7210 11020 7216
rect 9220 7200 9272 7206
rect 9220 7142 9272 7148
rect 7950 7100 8258 7109
rect 7950 7098 7956 7100
rect 8012 7098 8036 7100
rect 8092 7098 8116 7100
rect 8172 7098 8196 7100
rect 8252 7098 8258 7100
rect 8012 7046 8014 7098
rect 8194 7046 8196 7098
rect 7950 7044 7956 7046
rect 8012 7044 8036 7046
rect 8092 7044 8116 7046
rect 8172 7044 8196 7046
rect 8252 7044 8258 7046
rect 7950 7035 8258 7044
rect 9232 6934 9260 7142
rect 9220 6928 9272 6934
rect 9220 6870 9272 6876
rect 9324 6866 9352 7210
rect 9496 7200 9548 7206
rect 9496 7142 9548 7148
rect 9312 6860 9364 6866
rect 9312 6802 9364 6808
rect 8300 6792 8352 6798
rect 8300 6734 8352 6740
rect 8208 6656 8260 6662
rect 8208 6598 8260 6604
rect 8220 6458 8248 6598
rect 8208 6452 8260 6458
rect 8208 6394 8260 6400
rect 7950 6012 8258 6021
rect 7950 6010 7956 6012
rect 8012 6010 8036 6012
rect 8092 6010 8116 6012
rect 8172 6010 8196 6012
rect 8252 6010 8258 6012
rect 8012 5958 8014 6010
rect 8194 5958 8196 6010
rect 7950 5956 7956 5958
rect 8012 5956 8036 5958
rect 8092 5956 8116 5958
rect 8172 5956 8196 5958
rect 8252 5956 8258 5958
rect 7950 5947 8258 5956
rect 7950 4924 8258 4933
rect 7950 4922 7956 4924
rect 8012 4922 8036 4924
rect 8092 4922 8116 4924
rect 8172 4922 8196 4924
rect 8252 4922 8258 4924
rect 8012 4870 8014 4922
rect 8194 4870 8196 4922
rect 7950 4868 7956 4870
rect 8012 4868 8036 4870
rect 8092 4868 8116 4870
rect 8172 4868 8196 4870
rect 8252 4868 8258 4870
rect 7950 4859 8258 4868
rect 7950 3836 8258 3845
rect 7950 3834 7956 3836
rect 8012 3834 8036 3836
rect 8092 3834 8116 3836
rect 8172 3834 8196 3836
rect 8252 3834 8258 3836
rect 8012 3782 8014 3834
rect 8194 3782 8196 3834
rect 7950 3780 7956 3782
rect 8012 3780 8036 3782
rect 8092 3780 8116 3782
rect 8172 3780 8196 3782
rect 8252 3780 8258 3782
rect 7950 3771 8258 3780
rect 7950 2748 8258 2757
rect 7950 2746 7956 2748
rect 8012 2746 8036 2748
rect 8092 2746 8116 2748
rect 8172 2746 8196 2748
rect 8252 2746 8258 2748
rect 8012 2694 8014 2746
rect 8194 2694 8196 2746
rect 7950 2692 7956 2694
rect 8012 2692 8036 2694
rect 8092 2692 8116 2694
rect 8172 2692 8196 2694
rect 8252 2692 8258 2694
rect 7950 2683 8258 2692
rect 7944 56 8064 82
rect 8312 56 8340 6734
rect 9508 6730 9536 7142
rect 10980 6769 11008 7210
rect 10966 6760 11022 6769
rect 9496 6724 9548 6730
rect 10966 6695 11022 6704
rect 9496 6666 9548 6672
rect 9010 6556 9318 6565
rect 9010 6554 9016 6556
rect 9072 6554 9096 6556
rect 9152 6554 9176 6556
rect 9232 6554 9256 6556
rect 9312 6554 9318 6556
rect 9072 6502 9074 6554
rect 9254 6502 9256 6554
rect 9010 6500 9016 6502
rect 9072 6500 9096 6502
rect 9152 6500 9176 6502
rect 9232 6500 9256 6502
rect 9312 6500 9318 6502
rect 9010 6491 9318 6500
rect 8576 6316 8628 6322
rect 8576 6258 8628 6264
rect 8392 5568 8444 5574
rect 8392 5510 8444 5516
rect 8404 1834 8432 5510
rect 8392 1828 8444 1834
rect 8392 1770 8444 1776
rect 8588 56 8616 6258
rect 9588 6112 9640 6118
rect 9588 6054 9640 6060
rect 8852 5704 8904 5710
rect 8852 5646 8904 5652
rect 8864 56 8892 5646
rect 9010 5468 9318 5477
rect 9010 5466 9016 5468
rect 9072 5466 9096 5468
rect 9152 5466 9176 5468
rect 9232 5466 9256 5468
rect 9312 5466 9318 5468
rect 9072 5414 9074 5466
rect 9254 5414 9256 5466
rect 9010 5412 9016 5414
rect 9072 5412 9096 5414
rect 9152 5412 9176 5414
rect 9232 5412 9256 5414
rect 9312 5412 9318 5414
rect 9010 5403 9318 5412
rect 9496 5024 9548 5030
rect 9496 4966 9548 4972
rect 9010 4380 9318 4389
rect 9010 4378 9016 4380
rect 9072 4378 9096 4380
rect 9152 4378 9176 4380
rect 9232 4378 9256 4380
rect 9312 4378 9318 4380
rect 9072 4326 9074 4378
rect 9254 4326 9256 4378
rect 9010 4324 9016 4326
rect 9072 4324 9096 4326
rect 9152 4324 9176 4326
rect 9232 4324 9256 4326
rect 9312 4324 9318 4326
rect 9010 4315 9318 4324
rect 9404 3732 9456 3738
rect 9404 3674 9456 3680
rect 9010 3292 9318 3301
rect 9010 3290 9016 3292
rect 9072 3290 9096 3292
rect 9152 3290 9176 3292
rect 9232 3290 9256 3292
rect 9312 3290 9318 3292
rect 9072 3238 9074 3290
rect 9254 3238 9256 3290
rect 9010 3236 9016 3238
rect 9072 3236 9096 3238
rect 9152 3236 9176 3238
rect 9232 3236 9256 3238
rect 9312 3236 9318 3238
rect 9010 3227 9318 3236
rect 9010 2204 9318 2213
rect 9010 2202 9016 2204
rect 9072 2202 9096 2204
rect 9152 2202 9176 2204
rect 9232 2202 9256 2204
rect 9312 2202 9318 2204
rect 9072 2150 9074 2202
rect 9254 2150 9256 2202
rect 9010 2148 9016 2150
rect 9072 2148 9096 2150
rect 9152 2148 9176 2150
rect 9232 2148 9256 2150
rect 9312 2148 9318 2150
rect 9010 2139 9318 2148
rect 9416 218 9444 3674
rect 9508 2650 9536 4966
rect 9496 2644 9548 2650
rect 9496 2586 9548 2592
rect 9600 2514 9628 6054
rect 11900 5273 11928 7346
rect 12544 7206 12572 7670
rect 13372 7546 13400 7890
rect 12624 7540 12676 7546
rect 12624 7482 12676 7488
rect 13360 7540 13412 7546
rect 13360 7482 13412 7488
rect 13728 7540 13780 7546
rect 13728 7482 13780 7488
rect 12072 7200 12124 7206
rect 12072 7142 12124 7148
rect 12348 7200 12400 7206
rect 12348 7142 12400 7148
rect 12532 7200 12584 7206
rect 12532 7142 12584 7148
rect 12084 5914 12112 7142
rect 12360 7002 12388 7142
rect 12348 6996 12400 7002
rect 12348 6938 12400 6944
rect 12072 5908 12124 5914
rect 12072 5850 12124 5856
rect 12636 5386 12664 7482
rect 12716 7200 12768 7206
rect 12716 7142 12768 7148
rect 13084 7200 13136 7206
rect 13084 7142 13136 7148
rect 12728 5545 12756 7142
rect 13096 5778 13124 7142
rect 13360 6248 13412 6254
rect 13360 6190 13412 6196
rect 13084 5772 13136 5778
rect 13084 5714 13136 5720
rect 12714 5536 12770 5545
rect 12714 5471 12770 5480
rect 12532 5364 12584 5370
rect 12636 5358 12940 5386
rect 12532 5306 12584 5312
rect 11886 5264 11942 5273
rect 11886 5199 11942 5208
rect 11888 4684 11940 4690
rect 11888 4626 11940 4632
rect 10140 4276 10192 4282
rect 10140 4218 10192 4224
rect 9588 2508 9640 2514
rect 9588 2450 9640 2456
rect 9680 2032 9732 2038
rect 9680 1974 9732 1980
rect 9496 1352 9548 1358
rect 9496 1294 9548 1300
rect 9324 190 9444 218
rect 9140 56 9260 82
rect 7944 54 8078 56
rect 7944 42 7972 54
rect 7852 14 7972 42
rect 8022 0 8078 54
rect 8298 0 8354 56
rect 8574 0 8630 56
rect 8850 0 8906 56
rect 9126 54 9260 56
rect 9126 0 9182 54
rect 9232 42 9260 54
rect 9324 42 9352 190
rect 9508 82 9536 1294
rect 9416 56 9536 82
rect 9692 56 9720 1974
rect 9956 1760 10008 1766
rect 9956 1702 10008 1708
rect 9968 56 9996 1702
rect 10152 1698 10180 4218
rect 11612 3120 11664 3126
rect 11612 3062 11664 3068
rect 10782 2408 10838 2417
rect 10782 2343 10838 2352
rect 10140 1692 10192 1698
rect 10140 1634 10192 1640
rect 10506 1320 10562 1329
rect 10506 1255 10562 1264
rect 10230 1184 10286 1193
rect 10230 1119 10286 1128
rect 10244 56 10272 1119
rect 10520 56 10548 1255
rect 10796 56 10824 2343
rect 11336 2100 11388 2106
rect 11336 2042 11388 2048
rect 11060 1284 11112 1290
rect 11060 1226 11112 1232
rect 11072 56 11100 1226
rect 11348 56 11376 2042
rect 11624 56 11652 3062
rect 11900 56 11928 4626
rect 12440 4140 12492 4146
rect 12440 4082 12492 4088
rect 12348 3936 12400 3942
rect 12348 3878 12400 3884
rect 12164 3596 12216 3602
rect 12164 3538 12216 3544
rect 12176 56 12204 3538
rect 12360 2990 12388 3878
rect 12348 2984 12400 2990
rect 12348 2926 12400 2932
rect 12452 2854 12480 4082
rect 12544 4049 12572 5306
rect 12808 4752 12860 4758
rect 12808 4694 12860 4700
rect 12530 4040 12586 4049
rect 12530 3975 12586 3984
rect 12716 4004 12768 4010
rect 12716 3946 12768 3952
rect 12624 3936 12676 3942
rect 12624 3878 12676 3884
rect 12636 3670 12664 3878
rect 12624 3664 12676 3670
rect 12624 3606 12676 3612
rect 12532 3460 12584 3466
rect 12532 3402 12584 3408
rect 12440 2848 12492 2854
rect 12440 2790 12492 2796
rect 12544 1442 12572 3402
rect 12452 1414 12572 1442
rect 12452 56 12480 1414
rect 12728 56 12756 3946
rect 12820 2378 12848 4694
rect 12912 4604 12940 5358
rect 12912 4576 13216 4604
rect 13084 4480 13136 4486
rect 13084 4422 13136 4428
rect 12992 4140 13044 4146
rect 12992 4082 13044 4088
rect 12900 4072 12952 4078
rect 12900 4014 12952 4020
rect 12912 2922 12940 4014
rect 12900 2916 12952 2922
rect 12900 2858 12952 2864
rect 12808 2372 12860 2378
rect 12808 2314 12860 2320
rect 13004 56 13032 4082
rect 13096 3641 13124 4422
rect 13082 3632 13138 3641
rect 13082 3567 13138 3576
rect 13188 2582 13216 4576
rect 13268 2848 13320 2854
rect 13268 2790 13320 2796
rect 13176 2576 13228 2582
rect 13176 2518 13228 2524
rect 13280 56 13308 2790
rect 13372 1630 13400 6190
rect 13740 5817 13768 7482
rect 13912 7472 13964 7478
rect 13910 7440 13912 7449
rect 13964 7440 13966 7449
rect 13910 7375 13966 7384
rect 14200 7206 14228 7942
rect 14554 7919 14610 7928
rect 14280 7744 14332 7750
rect 14280 7686 14332 7692
rect 14292 7206 14320 7686
rect 14568 7410 14596 7919
rect 14464 7404 14516 7410
rect 14464 7346 14516 7352
rect 14556 7404 14608 7410
rect 14556 7346 14608 7352
rect 14188 7200 14240 7206
rect 14188 7142 14240 7148
rect 14280 7200 14332 7206
rect 14280 7142 14332 7148
rect 13950 7100 14258 7109
rect 13950 7098 13956 7100
rect 14012 7098 14036 7100
rect 14092 7098 14116 7100
rect 14172 7098 14196 7100
rect 14252 7098 14258 7100
rect 14012 7046 14014 7098
rect 14194 7046 14196 7098
rect 13950 7044 13956 7046
rect 14012 7044 14036 7046
rect 14092 7044 14116 7046
rect 14172 7044 14196 7046
rect 14252 7044 14258 7046
rect 13950 7035 14258 7044
rect 14476 6254 14504 7346
rect 14936 7206 14964 8298
rect 15120 7732 15148 8327
rect 15568 8084 15620 8090
rect 15568 8026 15620 8032
rect 15476 7880 15528 7886
rect 15476 7822 15528 7828
rect 15120 7704 15424 7732
rect 15010 7644 15318 7653
rect 15010 7642 15016 7644
rect 15072 7642 15096 7644
rect 15152 7642 15176 7644
rect 15232 7642 15256 7644
rect 15312 7642 15318 7644
rect 15072 7590 15074 7642
rect 15254 7590 15256 7642
rect 15010 7588 15016 7590
rect 15072 7588 15096 7590
rect 15152 7588 15176 7590
rect 15232 7588 15256 7590
rect 15312 7588 15318 7590
rect 15010 7579 15318 7588
rect 15396 7546 15424 7704
rect 15384 7540 15436 7546
rect 15384 7482 15436 7488
rect 15488 7274 15516 7822
rect 15384 7268 15436 7274
rect 15384 7210 15436 7216
rect 15476 7268 15528 7274
rect 15476 7210 15528 7216
rect 14924 7200 14976 7206
rect 14924 7142 14976 7148
rect 15010 6556 15318 6565
rect 15010 6554 15016 6556
rect 15072 6554 15096 6556
rect 15152 6554 15176 6556
rect 15232 6554 15256 6556
rect 15312 6554 15318 6556
rect 15072 6502 15074 6554
rect 15254 6502 15256 6554
rect 15010 6500 15016 6502
rect 15072 6500 15096 6502
rect 15152 6500 15176 6502
rect 15232 6500 15256 6502
rect 15312 6500 15318 6502
rect 15010 6491 15318 6500
rect 14740 6452 14792 6458
rect 14740 6394 14792 6400
rect 14464 6248 14516 6254
rect 14464 6190 14516 6196
rect 13950 6012 14258 6021
rect 13950 6010 13956 6012
rect 14012 6010 14036 6012
rect 14092 6010 14116 6012
rect 14172 6010 14196 6012
rect 14252 6010 14258 6012
rect 14012 5958 14014 6010
rect 14194 5958 14196 6010
rect 13950 5956 13956 5958
rect 14012 5956 14036 5958
rect 14092 5956 14116 5958
rect 14172 5956 14196 5958
rect 14252 5956 14258 5958
rect 13950 5947 14258 5956
rect 13726 5808 13782 5817
rect 13726 5743 13782 5752
rect 13636 5024 13688 5030
rect 13636 4966 13688 4972
rect 13544 4140 13596 4146
rect 13544 4082 13596 4088
rect 13556 3738 13584 4082
rect 13544 3732 13596 3738
rect 13544 3674 13596 3680
rect 13544 2916 13596 2922
rect 13544 2858 13596 2864
rect 13360 1624 13412 1630
rect 13360 1566 13412 1572
rect 13556 56 13584 2858
rect 13648 2446 13676 4966
rect 13950 4924 14258 4933
rect 13950 4922 13956 4924
rect 14012 4922 14036 4924
rect 14092 4922 14116 4924
rect 14172 4922 14196 4924
rect 14252 4922 14258 4924
rect 14012 4870 14014 4922
rect 14194 4870 14196 4922
rect 13950 4868 13956 4870
rect 14012 4868 14036 4870
rect 14092 4868 14116 4870
rect 14172 4868 14196 4870
rect 14252 4868 14258 4870
rect 13950 4859 14258 4868
rect 13912 4140 13964 4146
rect 13912 4082 13964 4088
rect 14464 4140 14516 4146
rect 14464 4082 14516 4088
rect 14556 4140 14608 4146
rect 14556 4082 14608 4088
rect 13728 3936 13780 3942
rect 13924 3924 13952 4082
rect 13728 3878 13780 3884
rect 13832 3896 13952 3924
rect 14280 3936 14332 3942
rect 13740 3738 13768 3878
rect 13728 3732 13780 3738
rect 13728 3674 13780 3680
rect 13832 3618 13860 3896
rect 14280 3878 14332 3884
rect 14372 3936 14424 3942
rect 14372 3878 14424 3884
rect 13950 3836 14258 3845
rect 13950 3834 13956 3836
rect 14012 3834 14036 3836
rect 14092 3834 14116 3836
rect 14172 3834 14196 3836
rect 14252 3834 14258 3836
rect 14012 3782 14014 3834
rect 14194 3782 14196 3834
rect 13950 3780 13956 3782
rect 14012 3780 14036 3782
rect 14092 3780 14116 3782
rect 14172 3780 14196 3782
rect 14252 3780 14258 3782
rect 13950 3771 14258 3780
rect 13740 3602 13860 3618
rect 14292 3602 14320 3878
rect 13728 3596 13860 3602
rect 13780 3590 13860 3596
rect 14280 3596 14332 3602
rect 13728 3538 13780 3544
rect 14280 3538 14332 3544
rect 13820 3528 13872 3534
rect 13820 3470 13872 3476
rect 14188 3528 14240 3534
rect 14188 3470 14240 3476
rect 13636 2440 13688 2446
rect 13636 2382 13688 2388
rect 13832 56 13860 3470
rect 14200 2904 14228 3470
rect 14384 3194 14412 3878
rect 14476 3466 14504 4082
rect 14464 3460 14516 3466
rect 14464 3402 14516 3408
rect 14372 3188 14424 3194
rect 14372 3130 14424 3136
rect 14200 2876 14320 2904
rect 13950 2748 14258 2757
rect 13950 2746 13956 2748
rect 14012 2746 14036 2748
rect 14092 2746 14116 2748
rect 14172 2746 14196 2748
rect 14252 2746 14258 2748
rect 14012 2694 14014 2746
rect 14194 2694 14196 2746
rect 13950 2692 13956 2694
rect 14012 2692 14036 2694
rect 14092 2692 14116 2694
rect 14172 2692 14196 2694
rect 14252 2692 14258 2694
rect 13950 2683 14258 2692
rect 14188 2644 14240 2650
rect 14188 2586 14240 2592
rect 14200 2310 14228 2586
rect 14096 2304 14148 2310
rect 14096 2246 14148 2252
rect 14188 2304 14240 2310
rect 14188 2246 14240 2252
rect 14108 56 14136 2246
rect 14292 2106 14320 2876
rect 14372 2848 14424 2854
rect 14372 2790 14424 2796
rect 14280 2100 14332 2106
rect 14280 2042 14332 2048
rect 14384 56 14412 2790
rect 14464 2440 14516 2446
rect 14464 2382 14516 2388
rect 14476 2310 14504 2382
rect 14464 2304 14516 2310
rect 14464 2246 14516 2252
rect 14568 1358 14596 4082
rect 14648 3936 14700 3942
rect 14648 3878 14700 3884
rect 14660 3466 14688 3878
rect 14648 3460 14700 3466
rect 14648 3402 14700 3408
rect 14752 3058 14780 6394
rect 15396 5846 15424 7210
rect 15580 6914 15608 8026
rect 16396 7948 16448 7954
rect 16396 7890 16448 7896
rect 16408 7546 16436 7890
rect 16856 7744 16908 7750
rect 16856 7686 16908 7692
rect 16396 7540 16448 7546
rect 16396 7482 16448 7488
rect 16580 7540 16632 7546
rect 16580 7482 16632 7488
rect 16304 7404 16356 7410
rect 16304 7346 16356 7352
rect 16316 6934 16344 7346
rect 16396 7336 16448 7342
rect 16396 7278 16448 7284
rect 15488 6886 15608 6914
rect 16304 6928 16356 6934
rect 15384 5840 15436 5846
rect 15384 5782 15436 5788
rect 15010 5468 15318 5477
rect 15010 5466 15016 5468
rect 15072 5466 15096 5468
rect 15152 5466 15176 5468
rect 15232 5466 15256 5468
rect 15312 5466 15318 5468
rect 15072 5414 15074 5466
rect 15254 5414 15256 5466
rect 15010 5412 15016 5414
rect 15072 5412 15096 5414
rect 15152 5412 15176 5414
rect 15232 5412 15256 5414
rect 15312 5412 15318 5414
rect 15010 5403 15318 5412
rect 15488 5030 15516 6886
rect 16408 6914 16436 7278
rect 16408 6886 16528 6914
rect 16304 6870 16356 6876
rect 16500 6798 16528 6886
rect 15568 6792 15620 6798
rect 15568 6734 15620 6740
rect 16488 6792 16540 6798
rect 16488 6734 16540 6740
rect 15476 5024 15528 5030
rect 15476 4966 15528 4972
rect 14924 4820 14976 4826
rect 14924 4762 14976 4768
rect 14832 4140 14884 4146
rect 14832 4082 14884 4088
rect 14844 3126 14872 4082
rect 14832 3120 14884 3126
rect 14832 3062 14884 3068
rect 14740 3052 14792 3058
rect 14740 2994 14792 3000
rect 14936 2446 14964 4762
rect 15384 4752 15436 4758
rect 15384 4694 15436 4700
rect 15010 4380 15318 4389
rect 15010 4378 15016 4380
rect 15072 4378 15096 4380
rect 15152 4378 15176 4380
rect 15232 4378 15256 4380
rect 15312 4378 15318 4380
rect 15072 4326 15074 4378
rect 15254 4326 15256 4378
rect 15010 4324 15016 4326
rect 15072 4324 15096 4326
rect 15152 4324 15176 4326
rect 15232 4324 15256 4326
rect 15312 4324 15318 4326
rect 15010 4315 15318 4324
rect 15200 4140 15252 4146
rect 15120 4100 15200 4128
rect 15120 3534 15148 4100
rect 15200 4082 15252 4088
rect 15292 3936 15344 3942
rect 15292 3878 15344 3884
rect 15304 3534 15332 3878
rect 15108 3528 15160 3534
rect 15108 3470 15160 3476
rect 15292 3528 15344 3534
rect 15292 3470 15344 3476
rect 15010 3292 15318 3301
rect 15010 3290 15016 3292
rect 15072 3290 15096 3292
rect 15152 3290 15176 3292
rect 15232 3290 15256 3292
rect 15312 3290 15318 3292
rect 15072 3238 15074 3290
rect 15254 3238 15256 3290
rect 15010 3236 15016 3238
rect 15072 3236 15096 3238
rect 15152 3236 15176 3238
rect 15232 3236 15256 3238
rect 15312 3236 15318 3238
rect 15010 3227 15318 3236
rect 15396 3058 15424 4694
rect 15476 3732 15528 3738
rect 15476 3674 15528 3680
rect 15384 3052 15436 3058
rect 15384 2994 15436 3000
rect 15384 2848 15436 2854
rect 15384 2790 15436 2796
rect 14924 2440 14976 2446
rect 14924 2382 14976 2388
rect 14648 2304 14700 2310
rect 14648 2246 14700 2252
rect 14924 2304 14976 2310
rect 14924 2246 14976 2252
rect 14556 1352 14608 1358
rect 14556 1294 14608 1300
rect 14660 56 14688 2246
rect 14936 56 14964 2246
rect 15010 2204 15318 2213
rect 15010 2202 15016 2204
rect 15072 2202 15096 2204
rect 15152 2202 15176 2204
rect 15232 2202 15256 2204
rect 15312 2202 15318 2204
rect 15072 2150 15074 2202
rect 15254 2150 15256 2202
rect 15010 2148 15016 2150
rect 15072 2148 15096 2150
rect 15152 2148 15176 2150
rect 15232 2148 15256 2150
rect 15312 2148 15318 2150
rect 15010 2139 15318 2148
rect 15212 56 15332 82
rect 9232 14 9352 42
rect 9402 54 9536 56
rect 9402 0 9458 54
rect 9678 0 9734 56
rect 9954 0 10010 56
rect 10230 0 10286 56
rect 10506 0 10562 56
rect 10782 0 10838 56
rect 11058 0 11114 56
rect 11334 0 11390 56
rect 11610 0 11666 56
rect 11886 0 11942 56
rect 12162 0 12218 56
rect 12438 0 12494 56
rect 12714 0 12770 56
rect 12990 0 13046 56
rect 13266 0 13322 56
rect 13542 0 13598 56
rect 13818 0 13874 56
rect 14094 0 14150 56
rect 14370 0 14426 56
rect 14646 0 14702 56
rect 14922 0 14978 56
rect 15198 54 15332 56
rect 15198 0 15254 54
rect 15304 42 15332 54
rect 15396 42 15424 2790
rect 15488 2582 15516 3674
rect 15476 2576 15528 2582
rect 15476 2518 15528 2524
rect 15580 2378 15608 6734
rect 16120 6656 16172 6662
rect 16592 6644 16620 7482
rect 16868 7206 16896 7686
rect 17144 7478 17172 9823
rect 17316 9376 17368 9382
rect 17316 9318 17368 9324
rect 17328 9178 17356 9318
rect 17316 9172 17368 9178
rect 17316 9114 17368 9120
rect 17408 9172 17460 9178
rect 17408 9114 17460 9120
rect 17420 8974 17448 9114
rect 17868 9036 17920 9042
rect 17868 8978 17920 8984
rect 17408 8968 17460 8974
rect 17408 8910 17460 8916
rect 17500 8968 17552 8974
rect 17500 8910 17552 8916
rect 17132 7472 17184 7478
rect 17132 7414 17184 7420
rect 17512 7206 17540 8910
rect 17880 7206 17908 8978
rect 18432 8634 18460 11194
rect 19524 9240 19576 9246
rect 19524 9182 19576 9188
rect 18420 8628 18472 8634
rect 18420 8570 18472 8576
rect 19156 8560 19208 8566
rect 19156 8502 19208 8508
rect 18788 8492 18840 8498
rect 18788 8434 18840 8440
rect 18144 7880 18196 7886
rect 18144 7822 18196 7828
rect 18156 7546 18184 7822
rect 18144 7540 18196 7546
rect 18144 7482 18196 7488
rect 16856 7200 16908 7206
rect 16856 7142 16908 7148
rect 17500 7200 17552 7206
rect 17500 7142 17552 7148
rect 17868 7200 17920 7206
rect 17868 7142 17920 7148
rect 17040 6860 17092 6866
rect 17040 6802 17092 6808
rect 16120 6598 16172 6604
rect 16500 6616 16620 6644
rect 16948 6656 17000 6662
rect 15936 3936 15988 3942
rect 15936 3878 15988 3884
rect 15948 3738 15976 3878
rect 15936 3732 15988 3738
rect 15936 3674 15988 3680
rect 15936 3392 15988 3398
rect 15936 3334 15988 3340
rect 15568 2372 15620 2378
rect 15568 2314 15620 2320
rect 15476 2304 15528 2310
rect 15476 2246 15528 2252
rect 15752 2304 15804 2310
rect 15752 2246 15804 2252
rect 15488 56 15516 2246
rect 15764 56 15792 2246
rect 15948 1970 15976 3334
rect 16132 3058 16160 6598
rect 16500 6225 16528 6616
rect 16948 6598 17000 6604
rect 16486 6216 16542 6225
rect 16486 6151 16542 6160
rect 16764 5636 16816 5642
rect 16764 5578 16816 5584
rect 16672 4140 16724 4146
rect 16672 4082 16724 4088
rect 16120 3052 16172 3058
rect 16120 2994 16172 3000
rect 16028 2848 16080 2854
rect 16028 2790 16080 2796
rect 15936 1964 15988 1970
rect 15936 1906 15988 1912
rect 16040 56 16068 2790
rect 16212 2440 16264 2446
rect 16212 2382 16264 2388
rect 16224 1630 16252 2382
rect 16304 2304 16356 2310
rect 16304 2246 16356 2252
rect 16580 2304 16632 2310
rect 16580 2246 16632 2252
rect 16212 1624 16264 1630
rect 16212 1566 16264 1572
rect 16316 56 16344 2246
rect 16592 56 16620 2246
rect 16684 1290 16712 4082
rect 16776 2446 16804 5578
rect 16960 5137 16988 6598
rect 17052 6390 17080 6802
rect 17224 6792 17276 6798
rect 17224 6734 17276 6740
rect 17236 6662 17264 6734
rect 17224 6656 17276 6662
rect 17224 6598 17276 6604
rect 17040 6384 17092 6390
rect 17040 6326 17092 6332
rect 18800 6186 18828 8434
rect 19168 8022 19196 8502
rect 19156 8016 19208 8022
rect 19156 7958 19208 7964
rect 19536 7478 19564 9182
rect 19996 8634 20024 11194
rect 21010 8732 21318 8741
rect 21010 8730 21016 8732
rect 21072 8730 21096 8732
rect 21152 8730 21176 8732
rect 21232 8730 21256 8732
rect 21312 8730 21318 8732
rect 21072 8678 21074 8730
rect 21254 8678 21256 8730
rect 21010 8676 21016 8678
rect 21072 8676 21096 8678
rect 21152 8676 21176 8678
rect 21232 8676 21256 8678
rect 21312 8676 21318 8678
rect 21010 8667 21318 8676
rect 21560 8634 21588 11194
rect 22928 8832 22980 8838
rect 22928 8774 22980 8780
rect 19984 8628 20036 8634
rect 19984 8570 20036 8576
rect 21548 8628 21600 8634
rect 21548 8570 21600 8576
rect 20352 8492 20404 8498
rect 20352 8434 20404 8440
rect 22192 8492 22244 8498
rect 22192 8434 22244 8440
rect 19950 8188 20258 8197
rect 19950 8186 19956 8188
rect 20012 8186 20036 8188
rect 20092 8186 20116 8188
rect 20172 8186 20196 8188
rect 20252 8186 20258 8188
rect 20012 8134 20014 8186
rect 20194 8134 20196 8186
rect 19950 8132 19956 8134
rect 20012 8132 20036 8134
rect 20092 8132 20116 8134
rect 20172 8132 20196 8134
rect 20252 8132 20258 8134
rect 19950 8123 20258 8132
rect 20260 8016 20312 8022
rect 20260 7958 20312 7964
rect 20272 7546 20300 7958
rect 20260 7540 20312 7546
rect 20260 7482 20312 7488
rect 19524 7472 19576 7478
rect 19524 7414 19576 7420
rect 19616 7404 19668 7410
rect 19616 7346 19668 7352
rect 19260 6718 19472 6746
rect 19260 6662 19288 6718
rect 19248 6656 19300 6662
rect 19248 6598 19300 6604
rect 19340 6656 19392 6662
rect 19340 6598 19392 6604
rect 18788 6180 18840 6186
rect 18788 6122 18840 6128
rect 17776 6112 17828 6118
rect 17776 6054 17828 6060
rect 16946 5128 17002 5137
rect 16946 5063 17002 5072
rect 17132 4140 17184 4146
rect 17132 4082 17184 4088
rect 16856 3936 16908 3942
rect 16856 3878 16908 3884
rect 16868 2922 16896 3878
rect 16856 2916 16908 2922
rect 16856 2858 16908 2864
rect 16764 2440 16816 2446
rect 16764 2382 16816 2388
rect 16948 2440 17000 2446
rect 17144 2417 17172 4082
rect 17316 3936 17368 3942
rect 17316 3878 17368 3884
rect 17408 3936 17460 3942
rect 17408 3878 17460 3884
rect 17328 3738 17356 3878
rect 17224 3732 17276 3738
rect 17224 3674 17276 3680
rect 17316 3732 17368 3738
rect 17316 3674 17368 3680
rect 17236 3398 17264 3674
rect 17224 3392 17276 3398
rect 17224 3334 17276 3340
rect 17420 3210 17448 3878
rect 17500 3596 17552 3602
rect 17500 3538 17552 3544
rect 17328 3182 17448 3210
rect 16948 2382 17000 2388
rect 17130 2408 17186 2417
rect 16856 2304 16908 2310
rect 16856 2246 16908 2252
rect 16672 1284 16724 1290
rect 16672 1226 16724 1232
rect 16868 56 16896 2246
rect 16960 1698 16988 2382
rect 17130 2343 17186 2352
rect 17132 2304 17184 2310
rect 17132 2246 17184 2252
rect 16948 1692 17000 1698
rect 16948 1634 17000 1640
rect 17144 56 17172 2246
rect 17328 1465 17356 3182
rect 17512 2446 17540 3538
rect 17788 2854 17816 6054
rect 17960 5568 18012 5574
rect 17960 5510 18012 5516
rect 18052 5568 18104 5574
rect 18052 5510 18104 5516
rect 17868 3460 17920 3466
rect 17868 3402 17920 3408
rect 17776 2848 17828 2854
rect 17776 2790 17828 2796
rect 17684 2644 17736 2650
rect 17684 2586 17736 2592
rect 17500 2440 17552 2446
rect 17500 2382 17552 2388
rect 17408 2304 17460 2310
rect 17408 2246 17460 2252
rect 17314 1456 17370 1465
rect 17314 1391 17370 1400
rect 17420 56 17448 2246
rect 17696 56 17724 2586
rect 17880 2106 17908 3402
rect 17972 2446 18000 5510
rect 18064 5370 18092 5510
rect 18052 5364 18104 5370
rect 18052 5306 18104 5312
rect 19352 4729 19380 6598
rect 19444 5302 19472 6718
rect 19432 5296 19484 5302
rect 19432 5238 19484 5244
rect 19432 5024 19484 5030
rect 19432 4966 19484 4972
rect 19338 4720 19394 4729
rect 19338 4655 19394 4664
rect 18052 4140 18104 4146
rect 18052 4082 18104 4088
rect 17960 2440 18012 2446
rect 17960 2382 18012 2388
rect 17960 2304 18012 2310
rect 17960 2246 18012 2252
rect 17868 2100 17920 2106
rect 17868 2042 17920 2048
rect 17972 56 18000 2246
rect 18064 1329 18092 4082
rect 18972 4072 19024 4078
rect 18972 4014 19024 4020
rect 18512 4004 18564 4010
rect 18512 3946 18564 3952
rect 18880 4004 18932 4010
rect 18880 3946 18932 3952
rect 18524 3126 18552 3946
rect 18696 3936 18748 3942
rect 18696 3878 18748 3884
rect 18512 3120 18564 3126
rect 18512 3062 18564 3068
rect 18512 2848 18564 2854
rect 18512 2790 18564 2796
rect 18236 2576 18288 2582
rect 18236 2518 18288 2524
rect 18050 1320 18106 1329
rect 18050 1255 18106 1264
rect 18248 56 18276 2518
rect 18524 2446 18552 2790
rect 18512 2440 18564 2446
rect 18512 2382 18564 2388
rect 18512 2304 18564 2310
rect 18512 2246 18564 2252
rect 18524 56 18552 2246
rect 18708 1698 18736 3878
rect 18892 2774 18920 3946
rect 18800 2746 18920 2774
rect 18696 1692 18748 1698
rect 18696 1634 18748 1640
rect 18800 1306 18828 2746
rect 18880 2644 18932 2650
rect 18880 2586 18932 2592
rect 18892 2038 18920 2586
rect 18984 2553 19012 4014
rect 19340 3528 19392 3534
rect 19340 3470 19392 3476
rect 19156 3392 19208 3398
rect 19156 3334 19208 3340
rect 19064 2576 19116 2582
rect 18970 2544 19026 2553
rect 19064 2518 19116 2524
rect 18970 2479 19026 2488
rect 18880 2032 18932 2038
rect 18880 1974 18932 1980
rect 18972 2032 19024 2038
rect 18972 1974 19024 1980
rect 18708 1278 18828 1306
rect 18708 1193 18736 1278
rect 18694 1184 18750 1193
rect 18694 1119 18750 1128
rect 18800 56 18920 82
rect 15304 14 15424 42
rect 15474 0 15530 56
rect 15750 0 15806 56
rect 16026 0 16082 56
rect 16302 0 16358 56
rect 16578 0 16634 56
rect 16854 0 16910 56
rect 17130 0 17186 56
rect 17406 0 17462 56
rect 17682 0 17738 56
rect 17958 0 18014 56
rect 18234 0 18290 56
rect 18510 0 18566 56
rect 18786 54 18920 56
rect 18786 0 18842 54
rect 18892 42 18920 54
rect 18984 42 19012 1974
rect 19076 1766 19104 2518
rect 19168 1766 19196 3334
rect 19352 2938 19380 3470
rect 19444 3058 19472 4966
rect 19524 3460 19576 3466
rect 19524 3402 19576 3408
rect 19432 3052 19484 3058
rect 19432 2994 19484 3000
rect 19352 2910 19472 2938
rect 19340 2848 19392 2854
rect 19340 2790 19392 2796
rect 19064 1760 19116 1766
rect 19064 1702 19116 1708
rect 19156 1760 19208 1766
rect 19156 1702 19208 1708
rect 19064 1420 19116 1426
rect 19064 1362 19116 1368
rect 19076 56 19104 1362
rect 19352 56 19380 2790
rect 19444 2582 19472 2910
rect 19536 2650 19564 3402
rect 19524 2644 19576 2650
rect 19524 2586 19576 2592
rect 19432 2576 19484 2582
rect 19628 2530 19656 7346
rect 19950 7100 20258 7109
rect 19950 7098 19956 7100
rect 20012 7098 20036 7100
rect 20092 7098 20116 7100
rect 20172 7098 20196 7100
rect 20252 7098 20258 7100
rect 20012 7046 20014 7098
rect 20194 7046 20196 7098
rect 19950 7044 19956 7046
rect 20012 7044 20036 7046
rect 20092 7044 20116 7046
rect 20172 7044 20196 7046
rect 20252 7044 20258 7046
rect 19950 7035 20258 7044
rect 19708 6656 19760 6662
rect 19708 6598 19760 6604
rect 19720 6458 19748 6598
rect 19708 6452 19760 6458
rect 19708 6394 19760 6400
rect 19950 6012 20258 6021
rect 19950 6010 19956 6012
rect 20012 6010 20036 6012
rect 20092 6010 20116 6012
rect 20172 6010 20196 6012
rect 20252 6010 20258 6012
rect 20012 5958 20014 6010
rect 20194 5958 20196 6010
rect 19950 5956 19956 5958
rect 20012 5956 20036 5958
rect 20092 5956 20116 5958
rect 20172 5956 20196 5958
rect 20252 5956 20258 5958
rect 19950 5947 20258 5956
rect 20364 5574 20392 8434
rect 20536 8424 20588 8430
rect 20536 8366 20588 8372
rect 20548 5642 20576 8366
rect 21640 8084 21692 8090
rect 21640 8026 21692 8032
rect 21652 7886 21680 8026
rect 21640 7880 21692 7886
rect 21640 7822 21692 7828
rect 21010 7644 21318 7653
rect 21010 7642 21016 7644
rect 21072 7642 21096 7644
rect 21152 7642 21176 7644
rect 21232 7642 21256 7644
rect 21312 7642 21318 7644
rect 21072 7590 21074 7642
rect 21254 7590 21256 7642
rect 21010 7588 21016 7590
rect 21072 7588 21096 7590
rect 21152 7588 21176 7590
rect 21232 7588 21256 7590
rect 21312 7588 21318 7590
rect 21010 7579 21318 7588
rect 21640 7540 21692 7546
rect 21640 7482 21692 7488
rect 20904 7404 20956 7410
rect 20904 7346 20956 7352
rect 20916 6934 20944 7346
rect 20904 6928 20956 6934
rect 20904 6870 20956 6876
rect 21010 6556 21318 6565
rect 21010 6554 21016 6556
rect 21072 6554 21096 6556
rect 21152 6554 21176 6556
rect 21232 6554 21256 6556
rect 21312 6554 21318 6556
rect 21072 6502 21074 6554
rect 21254 6502 21256 6554
rect 21010 6500 21016 6502
rect 21072 6500 21096 6502
rect 21152 6500 21176 6502
rect 21232 6500 21256 6502
rect 21312 6500 21318 6502
rect 21010 6491 21318 6500
rect 20904 6112 20956 6118
rect 20904 6054 20956 6060
rect 20536 5636 20588 5642
rect 20536 5578 20588 5584
rect 19800 5568 19852 5574
rect 19800 5510 19852 5516
rect 20352 5568 20404 5574
rect 20352 5510 20404 5516
rect 19812 4049 19840 5510
rect 19950 4924 20258 4933
rect 19950 4922 19956 4924
rect 20012 4922 20036 4924
rect 20092 4922 20116 4924
rect 20172 4922 20196 4924
rect 20252 4922 20258 4924
rect 20012 4870 20014 4922
rect 20194 4870 20196 4922
rect 19950 4868 19956 4870
rect 20012 4868 20036 4870
rect 20092 4868 20116 4870
rect 20172 4868 20196 4870
rect 20252 4868 20258 4870
rect 19950 4859 20258 4868
rect 20916 4593 20944 6054
rect 21010 5468 21318 5477
rect 21010 5466 21016 5468
rect 21072 5466 21096 5468
rect 21152 5466 21176 5468
rect 21232 5466 21256 5468
rect 21312 5466 21318 5468
rect 21072 5414 21074 5466
rect 21254 5414 21256 5466
rect 21010 5412 21016 5414
rect 21072 5412 21096 5414
rect 21152 5412 21176 5414
rect 21232 5412 21256 5414
rect 21312 5412 21318 5414
rect 21010 5403 21318 5412
rect 20902 4584 20958 4593
rect 20902 4519 20958 4528
rect 20352 4480 20404 4486
rect 20352 4422 20404 4428
rect 19798 4040 19854 4049
rect 19798 3975 19854 3984
rect 19800 3936 19852 3942
rect 19800 3878 19852 3884
rect 19812 2990 19840 3878
rect 19950 3836 20258 3845
rect 19950 3834 19956 3836
rect 20012 3834 20036 3836
rect 20092 3834 20116 3836
rect 20172 3834 20196 3836
rect 20252 3834 20258 3836
rect 20012 3782 20014 3834
rect 20194 3782 20196 3834
rect 19950 3780 19956 3782
rect 20012 3780 20036 3782
rect 20092 3780 20116 3782
rect 20172 3780 20196 3782
rect 20252 3780 20258 3782
rect 19950 3771 20258 3780
rect 19892 3664 19944 3670
rect 19892 3606 19944 3612
rect 19708 2984 19760 2990
rect 19708 2926 19760 2932
rect 19800 2984 19852 2990
rect 19800 2926 19852 2932
rect 19432 2518 19484 2524
rect 19536 2502 19656 2530
rect 19432 2440 19484 2446
rect 19432 2382 19484 2388
rect 19444 1834 19472 2382
rect 19432 1828 19484 1834
rect 19432 1770 19484 1776
rect 19536 1358 19564 2502
rect 19720 2417 19748 2926
rect 19904 2922 19932 3606
rect 20364 3466 20392 4422
rect 21010 4380 21318 4389
rect 21010 4378 21016 4380
rect 21072 4378 21096 4380
rect 21152 4378 21176 4380
rect 21232 4378 21256 4380
rect 21312 4378 21318 4380
rect 21072 4326 21074 4378
rect 21254 4326 21256 4378
rect 21010 4324 21016 4326
rect 21072 4324 21096 4326
rect 21152 4324 21176 4326
rect 21232 4324 21256 4326
rect 21312 4324 21318 4326
rect 21010 4315 21318 4324
rect 20904 4004 20956 4010
rect 20904 3946 20956 3952
rect 20720 3528 20772 3534
rect 20720 3470 20772 3476
rect 20352 3460 20404 3466
rect 20352 3402 20404 3408
rect 20260 3392 20312 3398
rect 20260 3334 20312 3340
rect 20444 3392 20496 3398
rect 20444 3334 20496 3340
rect 20272 3126 20300 3334
rect 20260 3120 20312 3126
rect 20260 3062 20312 3068
rect 20456 3040 20484 3334
rect 20628 3188 20680 3194
rect 20628 3130 20680 3136
rect 20364 3012 20484 3040
rect 19892 2916 19944 2922
rect 19892 2858 19944 2864
rect 19800 2848 19852 2854
rect 19800 2790 19852 2796
rect 19706 2408 19762 2417
rect 19706 2343 19762 2352
rect 19616 2304 19668 2310
rect 19616 2246 19668 2252
rect 19708 2304 19760 2310
rect 19708 2246 19760 2252
rect 19524 1352 19576 1358
rect 19524 1294 19576 1300
rect 19628 56 19656 2246
rect 19720 2038 19748 2246
rect 19812 2038 19840 2790
rect 19950 2748 20258 2757
rect 19950 2746 19956 2748
rect 20012 2746 20036 2748
rect 20092 2746 20116 2748
rect 20172 2746 20196 2748
rect 20252 2746 20258 2748
rect 20012 2694 20014 2746
rect 20194 2694 20196 2746
rect 19950 2692 19956 2694
rect 20012 2692 20036 2694
rect 20092 2692 20116 2694
rect 20172 2692 20196 2694
rect 20252 2692 20258 2694
rect 19950 2683 20258 2692
rect 19892 2576 19944 2582
rect 20364 2530 20392 3012
rect 20536 2916 20588 2922
rect 20536 2858 20588 2864
rect 20444 2848 20496 2854
rect 20444 2790 20496 2796
rect 19892 2518 19944 2524
rect 19708 2032 19760 2038
rect 19708 1974 19760 1980
rect 19800 2032 19852 2038
rect 19800 1974 19852 1980
rect 19904 56 19932 2518
rect 20088 2502 20392 2530
rect 19984 2440 20036 2446
rect 19984 2382 20036 2388
rect 19996 1902 20024 2382
rect 19984 1896 20036 1902
rect 19984 1838 20036 1844
rect 20088 1737 20116 2502
rect 20352 2440 20404 2446
rect 20352 2382 20404 2388
rect 20168 2304 20220 2310
rect 20168 2246 20220 2252
rect 20260 2304 20312 2310
rect 20260 2246 20312 2252
rect 20074 1728 20130 1737
rect 20074 1663 20130 1672
rect 20180 1426 20208 2246
rect 20168 1420 20220 1426
rect 20168 1362 20220 1368
rect 20272 1170 20300 2246
rect 20364 1970 20392 2382
rect 20352 1964 20404 1970
rect 20352 1906 20404 1912
rect 20180 1142 20300 1170
rect 20180 56 20208 1142
rect 20456 56 20484 2790
rect 20548 2514 20576 2858
rect 20536 2508 20588 2514
rect 20536 2450 20588 2456
rect 20534 2408 20590 2417
rect 20640 2378 20668 3130
rect 20534 2343 20536 2352
rect 20588 2343 20590 2352
rect 20628 2372 20680 2378
rect 20536 2314 20588 2320
rect 20628 2314 20680 2320
rect 20732 1873 20760 3470
rect 20812 3392 20864 3398
rect 20812 3334 20864 3340
rect 20824 3194 20852 3334
rect 20812 3188 20864 3194
rect 20812 3130 20864 3136
rect 20916 3058 20944 3946
rect 21456 3664 21508 3670
rect 21456 3606 21508 3612
rect 21364 3460 21416 3466
rect 21364 3402 21416 3408
rect 21010 3292 21318 3301
rect 21010 3290 21016 3292
rect 21072 3290 21096 3292
rect 21152 3290 21176 3292
rect 21232 3290 21256 3292
rect 21312 3290 21318 3292
rect 21072 3238 21074 3290
rect 21254 3238 21256 3290
rect 21010 3236 21016 3238
rect 21072 3236 21096 3238
rect 21152 3236 21176 3238
rect 21232 3236 21256 3238
rect 21312 3236 21318 3238
rect 21010 3227 21318 3236
rect 21376 3058 21404 3402
rect 20904 3052 20956 3058
rect 20904 2994 20956 3000
rect 21364 3052 21416 3058
rect 21364 2994 21416 3000
rect 21468 2922 21496 3606
rect 21456 2916 21508 2922
rect 21456 2858 21508 2864
rect 20812 2848 20864 2854
rect 20812 2790 20864 2796
rect 21548 2848 21600 2854
rect 21548 2790 21600 2796
rect 20718 1864 20774 1873
rect 20718 1799 20774 1808
rect 20824 1442 20852 2790
rect 21456 2644 21508 2650
rect 21456 2586 21508 2592
rect 21364 2304 21416 2310
rect 21364 2246 21416 2252
rect 21010 2204 21318 2213
rect 21010 2202 21016 2204
rect 21072 2202 21096 2204
rect 21152 2202 21176 2204
rect 21232 2202 21256 2204
rect 21312 2202 21318 2204
rect 21072 2150 21074 2202
rect 21254 2150 21256 2202
rect 21010 2148 21016 2150
rect 21072 2148 21096 2150
rect 21152 2148 21176 2150
rect 21232 2148 21256 2150
rect 21312 2148 21318 2150
rect 21010 2139 21318 2148
rect 20732 1414 20852 1442
rect 20732 56 20760 1414
rect 21376 218 21404 2246
rect 21192 190 21404 218
rect 21008 56 21128 82
rect 18892 14 19012 42
rect 19062 0 19118 56
rect 19338 0 19394 56
rect 19614 0 19670 56
rect 19890 0 19946 56
rect 20166 0 20222 56
rect 20442 0 20498 56
rect 20718 0 20774 56
rect 20994 54 21128 56
rect 20994 0 21050 54
rect 21100 42 21128 54
rect 21192 42 21220 190
rect 21284 56 21404 82
rect 21100 14 21220 42
rect 21270 54 21404 56
rect 21270 0 21326 54
rect 21376 42 21404 54
rect 21468 42 21496 2586
rect 21560 56 21588 2790
rect 21652 2689 21680 7482
rect 22008 4140 22060 4146
rect 22008 4082 22060 4088
rect 21732 3528 21784 3534
rect 21732 3470 21784 3476
rect 21638 2680 21694 2689
rect 21638 2615 21694 2624
rect 21640 2440 21692 2446
rect 21640 2382 21692 2388
rect 21652 2106 21680 2382
rect 21640 2100 21692 2106
rect 21640 2042 21692 2048
rect 21744 2009 21772 3470
rect 21824 2576 21876 2582
rect 21824 2518 21876 2524
rect 21730 2000 21786 2009
rect 21730 1935 21786 1944
rect 21836 56 21864 2518
rect 22020 2106 22048 4082
rect 22204 4010 22232 8434
rect 22940 7546 22968 8774
rect 23124 8634 23152 11194
rect 24216 9172 24268 9178
rect 24216 9114 24268 9120
rect 23388 8900 23440 8906
rect 23388 8842 23440 8848
rect 23112 8628 23164 8634
rect 23112 8570 23164 8576
rect 23112 8492 23164 8498
rect 23112 8434 23164 8440
rect 22928 7540 22980 7546
rect 22928 7482 22980 7488
rect 22836 6248 22888 6254
rect 22836 6190 22888 6196
rect 22376 4140 22428 4146
rect 22376 4082 22428 4088
rect 22192 4004 22244 4010
rect 22192 3946 22244 3952
rect 22388 3602 22416 4082
rect 22744 3732 22796 3738
rect 22744 3674 22796 3680
rect 22284 3596 22336 3602
rect 22284 3538 22336 3544
rect 22376 3596 22428 3602
rect 22376 3538 22428 3544
rect 22296 2514 22324 3538
rect 22756 3058 22784 3674
rect 22744 3052 22796 3058
rect 22744 2994 22796 3000
rect 22376 2916 22428 2922
rect 22376 2858 22428 2864
rect 22284 2508 22336 2514
rect 22284 2450 22336 2456
rect 22388 2446 22416 2858
rect 22652 2848 22704 2854
rect 22652 2790 22704 2796
rect 22468 2644 22520 2650
rect 22468 2586 22520 2592
rect 22376 2440 22428 2446
rect 22376 2382 22428 2388
rect 22100 2304 22152 2310
rect 22100 2246 22152 2252
rect 22008 2100 22060 2106
rect 22008 2042 22060 2048
rect 22112 56 22140 2246
rect 22480 1170 22508 2586
rect 22388 1142 22508 1170
rect 22388 56 22416 1142
rect 22664 56 22692 2790
rect 22744 2440 22796 2446
rect 22744 2382 22796 2388
rect 22756 1902 22784 2382
rect 22744 1896 22796 1902
rect 22744 1838 22796 1844
rect 22848 1154 22876 6190
rect 23020 5024 23072 5030
rect 23020 4966 23072 4972
rect 23032 4185 23060 4966
rect 23018 4176 23074 4185
rect 23018 4111 23074 4120
rect 23124 4010 23152 8434
rect 23400 5370 23428 8842
rect 23664 8492 23716 8498
rect 23664 8434 23716 8440
rect 23388 5364 23440 5370
rect 23388 5306 23440 5312
rect 23480 5024 23532 5030
rect 23480 4966 23532 4972
rect 23492 4690 23520 4966
rect 23480 4684 23532 4690
rect 23480 4626 23532 4632
rect 23296 4140 23348 4146
rect 23296 4082 23348 4088
rect 23112 4004 23164 4010
rect 23112 3946 23164 3952
rect 23308 3738 23336 4082
rect 23676 4010 23704 8434
rect 23940 7880 23992 7886
rect 23940 7822 23992 7828
rect 23952 7342 23980 7822
rect 24228 7546 24256 9114
rect 24688 8634 24716 11194
rect 24952 9444 25004 9450
rect 24952 9386 25004 9392
rect 24676 8628 24728 8634
rect 24676 8570 24728 8576
rect 24216 7540 24268 7546
rect 24216 7482 24268 7488
rect 24308 7404 24360 7410
rect 24308 7346 24360 7352
rect 23940 7336 23992 7342
rect 23940 7278 23992 7284
rect 24032 7336 24084 7342
rect 24032 7278 24084 7284
rect 23664 4004 23716 4010
rect 23664 3946 23716 3952
rect 23296 3732 23348 3738
rect 23296 3674 23348 3680
rect 23940 3460 23992 3466
rect 23940 3402 23992 3408
rect 23204 2848 23256 2854
rect 23204 2790 23256 2796
rect 23756 2848 23808 2854
rect 23756 2790 23808 2796
rect 22928 2576 22980 2582
rect 22928 2518 22980 2524
rect 22836 1148 22888 1154
rect 22836 1090 22888 1096
rect 22940 56 22968 2518
rect 23216 56 23244 2790
rect 23296 2440 23348 2446
rect 23296 2382 23348 2388
rect 23664 2440 23716 2446
rect 23664 2382 23716 2388
rect 23308 2038 23336 2382
rect 23572 2304 23624 2310
rect 23492 2264 23572 2292
rect 23296 2032 23348 2038
rect 23296 1974 23348 1980
rect 23492 56 23520 2264
rect 23572 2246 23624 2252
rect 23676 2106 23704 2382
rect 23664 2100 23716 2106
rect 23664 2042 23716 2048
rect 23768 56 23796 2790
rect 23952 2514 23980 3402
rect 23940 2508 23992 2514
rect 23940 2450 23992 2456
rect 24044 56 24072 7278
rect 24124 3664 24176 3670
rect 24124 3606 24176 3612
rect 24136 2582 24164 3606
rect 24124 2576 24176 2582
rect 24124 2518 24176 2524
rect 24320 56 24348 7346
rect 24584 6928 24636 6934
rect 24584 6870 24636 6876
rect 24596 56 24624 6870
rect 24964 6662 24992 9386
rect 25320 9376 25372 9382
rect 25320 9318 25372 9324
rect 25134 8528 25190 8537
rect 25134 8463 25190 8472
rect 25044 8424 25096 8430
rect 25044 8366 25096 8372
rect 24952 6656 25004 6662
rect 24952 6598 25004 6604
rect 25056 4826 25084 8366
rect 25148 7546 25176 8463
rect 25332 7546 25360 9318
rect 26252 8634 26280 11194
rect 27010 8732 27318 8741
rect 27010 8730 27016 8732
rect 27072 8730 27096 8732
rect 27152 8730 27176 8732
rect 27232 8730 27256 8732
rect 27312 8730 27318 8732
rect 27072 8678 27074 8730
rect 27254 8678 27256 8730
rect 27010 8676 27016 8678
rect 27072 8676 27096 8678
rect 27152 8676 27176 8678
rect 27232 8676 27256 8678
rect 27312 8676 27318 8678
rect 27010 8667 27318 8676
rect 27816 8634 27844 11194
rect 29380 8634 29408 11194
rect 30102 9888 30158 9897
rect 30102 9823 30158 9832
rect 29920 8968 29972 8974
rect 29920 8910 29972 8916
rect 26240 8628 26292 8634
rect 26240 8570 26292 8576
rect 27804 8628 27856 8634
rect 27804 8570 27856 8576
rect 29368 8628 29420 8634
rect 29368 8570 29420 8576
rect 29932 8498 29960 8910
rect 30116 8634 30144 9823
rect 30838 9616 30894 9625
rect 30838 9551 30894 9560
rect 30656 9308 30708 9314
rect 30656 9250 30708 9256
rect 30288 9104 30340 9110
rect 30288 9046 30340 9052
rect 30470 9072 30526 9081
rect 30104 8628 30156 8634
rect 30104 8570 30156 8576
rect 30300 8498 30328 9046
rect 30470 9007 30526 9016
rect 30484 8634 30512 9007
rect 30472 8628 30524 8634
rect 30472 8570 30524 8576
rect 30668 8498 30696 9250
rect 26424 8492 26476 8498
rect 26424 8434 26476 8440
rect 29000 8492 29052 8498
rect 29000 8434 29052 8440
rect 29920 8492 29972 8498
rect 29920 8434 29972 8440
rect 30288 8492 30340 8498
rect 30288 8434 30340 8440
rect 30656 8492 30708 8498
rect 30656 8434 30708 8440
rect 25950 8188 26258 8197
rect 25950 8186 25956 8188
rect 26012 8186 26036 8188
rect 26092 8186 26116 8188
rect 26172 8186 26196 8188
rect 26252 8186 26258 8188
rect 26012 8134 26014 8186
rect 26194 8134 26196 8186
rect 25950 8132 25956 8134
rect 26012 8132 26036 8134
rect 26092 8132 26116 8134
rect 26172 8132 26196 8134
rect 26252 8132 26258 8134
rect 25950 8123 26258 8132
rect 25136 7540 25188 7546
rect 25136 7482 25188 7488
rect 25320 7540 25372 7546
rect 25320 7482 25372 7488
rect 25688 7472 25740 7478
rect 25688 7414 25740 7420
rect 25136 6180 25188 6186
rect 25136 6122 25188 6128
rect 25044 4820 25096 4826
rect 25044 4762 25096 4768
rect 24858 2680 24914 2689
rect 24858 2615 24914 2624
rect 24872 56 24900 2615
rect 25148 56 25176 6122
rect 25226 3496 25282 3505
rect 25226 3431 25228 3440
rect 25280 3431 25282 3440
rect 25228 3402 25280 3408
rect 25412 1352 25464 1358
rect 25412 1294 25464 1300
rect 25424 56 25452 1294
rect 25700 56 25728 7414
rect 25872 7404 25924 7410
rect 25872 7346 25924 7352
rect 25780 3392 25832 3398
rect 25780 3334 25832 3340
rect 25792 3097 25820 3334
rect 25778 3088 25834 3097
rect 25778 3023 25834 3032
rect 25884 1442 25912 7346
rect 25950 7100 26258 7109
rect 25950 7098 25956 7100
rect 26012 7098 26036 7100
rect 26092 7098 26116 7100
rect 26172 7098 26196 7100
rect 26252 7098 26258 7100
rect 26012 7046 26014 7098
rect 26194 7046 26196 7098
rect 25950 7044 25956 7046
rect 26012 7044 26036 7046
rect 26092 7044 26116 7046
rect 26172 7044 26196 7046
rect 26252 7044 26258 7046
rect 25950 7035 26258 7044
rect 26332 6792 26384 6798
rect 26332 6734 26384 6740
rect 25950 6012 26258 6021
rect 25950 6010 25956 6012
rect 26012 6010 26036 6012
rect 26092 6010 26116 6012
rect 26172 6010 26196 6012
rect 26252 6010 26258 6012
rect 26012 5958 26014 6010
rect 26194 5958 26196 6010
rect 25950 5956 25956 5958
rect 26012 5956 26036 5958
rect 26092 5956 26116 5958
rect 26172 5956 26196 5958
rect 26252 5956 26258 5958
rect 25950 5947 26258 5956
rect 26056 5568 26108 5574
rect 26108 5528 26280 5556
rect 26056 5510 26108 5516
rect 26252 5166 26280 5528
rect 26240 5160 26292 5166
rect 26240 5102 26292 5108
rect 25950 4924 26258 4933
rect 25950 4922 25956 4924
rect 26012 4922 26036 4924
rect 26092 4922 26116 4924
rect 26172 4922 26196 4924
rect 26252 4922 26258 4924
rect 26012 4870 26014 4922
rect 26194 4870 26196 4922
rect 25950 4868 25956 4870
rect 26012 4868 26036 4870
rect 26092 4868 26116 4870
rect 26172 4868 26196 4870
rect 26252 4868 26258 4870
rect 25950 4859 26258 4868
rect 25950 3836 26258 3845
rect 25950 3834 25956 3836
rect 26012 3834 26036 3836
rect 26092 3834 26116 3836
rect 26172 3834 26196 3836
rect 26252 3834 26258 3836
rect 26012 3782 26014 3834
rect 26194 3782 26196 3834
rect 25950 3780 25956 3782
rect 26012 3780 26036 3782
rect 26092 3780 26116 3782
rect 26172 3780 26196 3782
rect 26252 3780 26258 3782
rect 25950 3771 26258 3780
rect 26240 3392 26292 3398
rect 26240 3334 26292 3340
rect 26252 2961 26280 3334
rect 26238 2952 26294 2961
rect 26238 2887 26294 2896
rect 25950 2748 26258 2757
rect 25950 2746 25956 2748
rect 26012 2746 26036 2748
rect 26092 2746 26116 2748
rect 26172 2746 26196 2748
rect 26252 2746 26258 2748
rect 26012 2694 26014 2746
rect 26194 2694 26196 2746
rect 25950 2692 25956 2694
rect 26012 2692 26036 2694
rect 26092 2692 26116 2694
rect 26172 2692 26196 2694
rect 26252 2692 26258 2694
rect 25950 2683 26258 2692
rect 26344 1578 26372 6734
rect 26436 4010 26464 8434
rect 26792 8016 26844 8022
rect 26792 7958 26844 7964
rect 26804 7750 26832 7958
rect 26792 7744 26844 7750
rect 26792 7686 26844 7692
rect 27010 7644 27318 7653
rect 27010 7642 27016 7644
rect 27072 7642 27096 7644
rect 27152 7642 27176 7644
rect 27232 7642 27256 7644
rect 27312 7642 27318 7644
rect 27072 7590 27074 7642
rect 27254 7590 27256 7642
rect 27010 7588 27016 7590
rect 27072 7588 27096 7590
rect 27152 7588 27176 7590
rect 27232 7588 27256 7590
rect 27312 7588 27318 7590
rect 27010 7579 27318 7588
rect 27010 6556 27318 6565
rect 27010 6554 27016 6556
rect 27072 6554 27096 6556
rect 27152 6554 27176 6556
rect 27232 6554 27256 6556
rect 27312 6554 27318 6556
rect 27072 6502 27074 6554
rect 27254 6502 27256 6554
rect 27010 6500 27016 6502
rect 27072 6500 27096 6502
rect 27152 6500 27176 6502
rect 27232 6500 27256 6502
rect 27312 6500 27318 6502
rect 27010 6491 27318 6500
rect 27620 6452 27672 6458
rect 27620 6394 27672 6400
rect 26792 5568 26844 5574
rect 26792 5510 26844 5516
rect 26516 5228 26568 5234
rect 26516 5170 26568 5176
rect 26424 4004 26476 4010
rect 26424 3946 26476 3952
rect 26252 1550 26372 1578
rect 25884 1414 26004 1442
rect 25976 56 26004 1414
rect 26252 56 26280 1550
rect 26528 56 26556 5170
rect 26804 56 26832 5510
rect 27010 5468 27318 5477
rect 27010 5466 27016 5468
rect 27072 5466 27096 5468
rect 27152 5466 27176 5468
rect 27232 5466 27256 5468
rect 27312 5466 27318 5468
rect 27072 5414 27074 5466
rect 27254 5414 27256 5466
rect 27010 5412 27016 5414
rect 27072 5412 27096 5414
rect 27152 5412 27176 5414
rect 27232 5412 27256 5414
rect 27312 5412 27318 5414
rect 27010 5403 27318 5412
rect 27632 5166 27660 6394
rect 29012 5370 29040 8434
rect 30472 8424 30524 8430
rect 30472 8366 30524 8372
rect 30380 8084 30432 8090
rect 30380 8026 30432 8032
rect 30392 6322 30420 8026
rect 30380 6316 30432 6322
rect 30380 6258 30432 6264
rect 30484 5846 30512 8366
rect 30852 8090 30880 9551
rect 30944 8634 30972 11194
rect 31482 9344 31538 9353
rect 31482 9279 31538 9288
rect 31022 8800 31078 8809
rect 31022 8735 31078 8744
rect 30932 8628 30984 8634
rect 30932 8570 30984 8576
rect 31036 8090 31064 8735
rect 31390 8528 31446 8537
rect 31390 8463 31446 8472
rect 31404 8090 31432 8463
rect 30840 8084 30892 8090
rect 30840 8026 30892 8032
rect 31024 8084 31076 8090
rect 31024 8026 31076 8032
rect 31392 8084 31444 8090
rect 31392 8026 31444 8032
rect 30840 7880 30892 7886
rect 30840 7822 30892 7828
rect 30852 7002 30880 7822
rect 31496 7546 31524 9279
rect 32404 8424 32456 8430
rect 32404 8366 32456 8372
rect 31852 8356 31904 8362
rect 31852 8298 31904 8304
rect 31864 7993 31892 8298
rect 32416 8265 32444 8366
rect 32402 8256 32458 8265
rect 31950 8188 32258 8197
rect 32402 8191 32458 8200
rect 31950 8186 31956 8188
rect 32012 8186 32036 8188
rect 32092 8186 32116 8188
rect 32172 8186 32196 8188
rect 32252 8186 32258 8188
rect 32012 8134 32014 8186
rect 32194 8134 32196 8186
rect 31950 8132 31956 8134
rect 32012 8132 32036 8134
rect 32092 8132 32116 8134
rect 32172 8132 32196 8134
rect 32252 8132 32258 8134
rect 31950 8123 32258 8132
rect 31850 7984 31906 7993
rect 31850 7919 31906 7928
rect 31760 7744 31812 7750
rect 32128 7744 32180 7750
rect 31760 7686 31812 7692
rect 32126 7712 32128 7721
rect 32180 7712 32182 7721
rect 31484 7540 31536 7546
rect 31484 7482 31536 7488
rect 31772 7449 31800 7686
rect 32126 7647 32182 7656
rect 31758 7440 31814 7449
rect 31300 7404 31352 7410
rect 31758 7375 31814 7384
rect 31300 7346 31352 7352
rect 31312 7313 31340 7346
rect 31298 7304 31354 7313
rect 31298 7239 31354 7248
rect 31950 7100 32258 7109
rect 31950 7098 31956 7100
rect 32012 7098 32036 7100
rect 32092 7098 32116 7100
rect 32172 7098 32196 7100
rect 32252 7098 32258 7100
rect 32012 7046 32014 7098
rect 32194 7046 32196 7098
rect 31950 7044 31956 7046
rect 32012 7044 32036 7046
rect 32092 7044 32116 7046
rect 32172 7044 32196 7046
rect 32252 7044 32258 7046
rect 31950 7035 32258 7044
rect 30840 6996 30892 7002
rect 30840 6938 30892 6944
rect 32508 6914 32536 11194
rect 32772 7200 32824 7206
rect 32770 7168 32772 7177
rect 32824 7168 32826 7177
rect 32770 7103 32826 7112
rect 31758 6896 31814 6905
rect 31758 6831 31814 6840
rect 32324 6886 32536 6914
rect 31576 6792 31628 6798
rect 31576 6734 31628 6740
rect 31668 6792 31720 6798
rect 31668 6734 31720 6740
rect 31484 6724 31536 6730
rect 31484 6666 31536 6672
rect 31392 6656 31444 6662
rect 31390 6624 31392 6633
rect 31444 6624 31446 6633
rect 31390 6559 31446 6568
rect 31496 6322 31524 6666
rect 31588 6390 31616 6734
rect 31576 6384 31628 6390
rect 31576 6326 31628 6332
rect 31484 6316 31536 6322
rect 31484 6258 31536 6264
rect 31482 6216 31538 6225
rect 31482 6151 31538 6160
rect 31496 6118 31524 6151
rect 31484 6112 31536 6118
rect 31484 6054 31536 6060
rect 31208 5908 31260 5914
rect 31208 5850 31260 5856
rect 30472 5840 30524 5846
rect 30472 5782 30524 5788
rect 31220 5710 31248 5850
rect 29276 5704 29328 5710
rect 29276 5646 29328 5652
rect 29552 5704 29604 5710
rect 29552 5646 29604 5652
rect 31208 5704 31260 5710
rect 31208 5646 31260 5652
rect 29000 5364 29052 5370
rect 29000 5306 29052 5312
rect 29092 5228 29144 5234
rect 29092 5170 29144 5176
rect 27344 5160 27396 5166
rect 27344 5102 27396 5108
rect 27620 5160 27672 5166
rect 27620 5102 27672 5108
rect 27010 4380 27318 4389
rect 27010 4378 27016 4380
rect 27072 4378 27096 4380
rect 27152 4378 27176 4380
rect 27232 4378 27256 4380
rect 27312 4378 27318 4380
rect 27072 4326 27074 4378
rect 27254 4326 27256 4378
rect 27010 4324 27016 4326
rect 27072 4324 27096 4326
rect 27152 4324 27176 4326
rect 27232 4324 27256 4326
rect 27312 4324 27318 4326
rect 27010 4315 27318 4324
rect 27010 3292 27318 3301
rect 27010 3290 27016 3292
rect 27072 3290 27096 3292
rect 27152 3290 27176 3292
rect 27232 3290 27256 3292
rect 27312 3290 27318 3292
rect 27072 3238 27074 3290
rect 27254 3238 27256 3290
rect 27010 3236 27016 3238
rect 27072 3236 27096 3238
rect 27152 3236 27176 3238
rect 27232 3236 27256 3238
rect 27312 3236 27318 3238
rect 27010 3227 27318 3236
rect 27010 2204 27318 2213
rect 27010 2202 27016 2204
rect 27072 2202 27096 2204
rect 27152 2202 27176 2204
rect 27232 2202 27256 2204
rect 27312 2202 27318 2204
rect 27072 2150 27074 2202
rect 27254 2150 27256 2202
rect 27010 2148 27016 2150
rect 27072 2148 27096 2150
rect 27152 2148 27176 2150
rect 27232 2148 27256 2150
rect 27312 2148 27318 2150
rect 27010 2139 27318 2148
rect 27068 1148 27120 1154
rect 27068 1090 27120 1096
rect 27080 56 27108 1090
rect 27356 56 27384 5102
rect 28724 4548 28776 4554
rect 28724 4490 28776 4496
rect 28448 4140 28500 4146
rect 28448 4082 28500 4088
rect 28172 4072 28224 4078
rect 28172 4014 28224 4020
rect 27896 3732 27948 3738
rect 27896 3674 27948 3680
rect 27620 3596 27672 3602
rect 27620 3538 27672 3544
rect 27632 56 27660 3538
rect 27908 56 27936 3674
rect 28184 56 28212 4014
rect 28460 56 28488 4082
rect 28736 56 28764 4490
rect 29000 4072 29052 4078
rect 28998 4040 29000 4049
rect 29052 4040 29054 4049
rect 28998 3975 29054 3984
rect 29104 2666 29132 5170
rect 29012 2638 29132 2666
rect 29012 56 29040 2638
rect 29288 56 29316 5646
rect 29564 56 29592 5646
rect 31680 5574 31708 6734
rect 31772 6662 31800 6831
rect 32324 6662 32352 6886
rect 31760 6656 31812 6662
rect 31760 6598 31812 6604
rect 32312 6656 32364 6662
rect 32312 6598 32364 6604
rect 31852 6452 31904 6458
rect 31852 6394 31904 6400
rect 31864 6361 31892 6394
rect 31850 6352 31906 6361
rect 31850 6287 31906 6296
rect 31852 6112 31904 6118
rect 31852 6054 31904 6060
rect 31668 5568 31720 5574
rect 31760 5568 31812 5574
rect 31668 5510 31720 5516
rect 31758 5536 31760 5545
rect 31812 5536 31814 5545
rect 31758 5471 31814 5480
rect 31484 5024 31536 5030
rect 31484 4966 31536 4972
rect 31496 4729 31524 4966
rect 31482 4720 31538 4729
rect 31482 4655 31538 4664
rect 31864 4622 31892 6054
rect 31950 6012 32258 6021
rect 31950 6010 31956 6012
rect 32012 6010 32036 6012
rect 32092 6010 32116 6012
rect 32172 6010 32196 6012
rect 32252 6010 32258 6012
rect 32012 5958 32014 6010
rect 32194 5958 32196 6010
rect 31950 5956 31956 5958
rect 32012 5956 32036 5958
rect 32092 5956 32116 5958
rect 32172 5956 32196 5958
rect 32252 5956 32258 5958
rect 31950 5947 32258 5956
rect 32036 5840 32088 5846
rect 32128 5840 32180 5846
rect 32036 5782 32088 5788
rect 32126 5808 32128 5817
rect 32180 5808 32182 5817
rect 32048 5273 32076 5782
rect 32126 5743 32182 5752
rect 32034 5264 32090 5273
rect 32034 5199 32090 5208
rect 32864 5024 32916 5030
rect 32862 4992 32864 5001
rect 32916 4992 32918 5001
rect 31950 4924 32258 4933
rect 32862 4927 32918 4936
rect 31950 4922 31956 4924
rect 32012 4922 32036 4924
rect 32092 4922 32116 4924
rect 32172 4922 32196 4924
rect 32252 4922 32258 4924
rect 32012 4870 32014 4922
rect 32194 4870 32196 4922
rect 31950 4868 31956 4870
rect 32012 4868 32036 4870
rect 32092 4868 32116 4870
rect 32172 4868 32196 4870
rect 32252 4868 32258 4870
rect 31950 4859 32258 4868
rect 31852 4616 31904 4622
rect 31852 4558 31904 4564
rect 31300 4480 31352 4486
rect 31300 4422 31352 4428
rect 31760 4480 31812 4486
rect 32128 4480 32180 4486
rect 31760 4422 31812 4428
rect 32126 4448 32128 4457
rect 32180 4448 32182 4457
rect 31312 4146 31340 4422
rect 31772 4185 31800 4422
rect 32126 4383 32182 4392
rect 31758 4176 31814 4185
rect 31300 4140 31352 4146
rect 31758 4111 31814 4120
rect 31300 4082 31352 4088
rect 31300 3936 31352 3942
rect 31300 3878 31352 3884
rect 31484 3936 31536 3942
rect 32864 3936 32916 3942
rect 31484 3878 31536 3884
rect 32862 3904 32864 3913
rect 32916 3904 32918 3913
rect 30932 3188 30984 3194
rect 30932 3130 30984 3136
rect 30944 2446 30972 3130
rect 31312 3058 31340 3878
rect 31496 3641 31524 3878
rect 31950 3836 32258 3845
rect 32862 3839 32918 3848
rect 31950 3834 31956 3836
rect 32012 3834 32036 3836
rect 32092 3834 32116 3836
rect 32172 3834 32196 3836
rect 32252 3834 32258 3836
rect 32012 3782 32014 3834
rect 32194 3782 32196 3834
rect 31950 3780 31956 3782
rect 32012 3780 32036 3782
rect 32092 3780 32116 3782
rect 32172 3780 32196 3782
rect 32252 3780 32258 3782
rect 31950 3771 32258 3780
rect 31482 3632 31538 3641
rect 31482 3567 31538 3576
rect 31668 3392 31720 3398
rect 31668 3334 31720 3340
rect 31760 3392 31812 3398
rect 32128 3392 32180 3398
rect 31760 3334 31812 3340
rect 32126 3360 32128 3369
rect 32180 3360 32182 3369
rect 31680 3058 31708 3334
rect 31772 3097 31800 3334
rect 32126 3295 32182 3304
rect 31758 3088 31814 3097
rect 31300 3052 31352 3058
rect 31300 2994 31352 3000
rect 31668 3052 31720 3058
rect 31758 3023 31814 3032
rect 31668 2994 31720 3000
rect 31760 2848 31812 2854
rect 32864 2848 32916 2854
rect 31760 2790 31812 2796
rect 32862 2816 32864 2825
rect 32916 2816 32918 2825
rect 31772 2553 31800 2790
rect 31950 2748 32258 2757
rect 32862 2751 32918 2760
rect 31950 2746 31956 2748
rect 32012 2746 32036 2748
rect 32092 2746 32116 2748
rect 32172 2746 32196 2748
rect 32252 2746 32258 2748
rect 32012 2694 32014 2746
rect 32194 2694 32196 2746
rect 31950 2692 31956 2694
rect 32012 2692 32036 2694
rect 32092 2692 32116 2694
rect 32172 2692 32196 2694
rect 32252 2692 32258 2694
rect 31950 2683 32258 2692
rect 31758 2544 31814 2553
rect 31758 2479 31814 2488
rect 30932 2440 30984 2446
rect 30932 2382 30984 2388
rect 31300 2440 31352 2446
rect 31300 2382 31352 2388
rect 30748 2304 30800 2310
rect 30748 2246 30800 2252
rect 31116 2304 31168 2310
rect 31116 2246 31168 2252
rect 30760 2009 30788 2246
rect 30746 2000 30802 2009
rect 30746 1935 30802 1944
rect 31128 1737 31156 2246
rect 31114 1728 31170 1737
rect 31312 1698 31340 2382
rect 31484 2304 31536 2310
rect 31852 2304 31904 2310
rect 31484 2246 31536 2252
rect 31850 2272 31852 2281
rect 31904 2272 31906 2281
rect 31114 1663 31170 1672
rect 31300 1692 31352 1698
rect 31300 1634 31352 1640
rect 31496 1465 31524 2246
rect 31850 2207 31906 2216
rect 31482 1456 31538 1465
rect 31482 1391 31538 1400
rect 21376 14 21496 42
rect 21546 0 21602 56
rect 21822 0 21878 56
rect 22098 0 22154 56
rect 22374 0 22430 56
rect 22650 0 22706 56
rect 22926 0 22982 56
rect 23202 0 23258 56
rect 23478 0 23534 56
rect 23754 0 23810 56
rect 24030 0 24086 56
rect 24306 0 24362 56
rect 24582 0 24638 56
rect 24858 0 24914 56
rect 25134 0 25190 56
rect 25410 0 25466 56
rect 25686 0 25742 56
rect 25962 0 26018 56
rect 26238 0 26294 56
rect 26514 0 26570 56
rect 26790 0 26846 56
rect 27066 0 27122 56
rect 27342 0 27398 56
rect 27618 0 27674 56
rect 27894 0 27950 56
rect 28170 0 28226 56
rect 28446 0 28502 56
rect 28722 0 28778 56
rect 28998 0 29054 56
rect 29274 0 29330 56
rect 29550 0 29606 56
<< via2 >>
rect 3016 8730 3072 8732
rect 3096 8730 3152 8732
rect 3176 8730 3232 8732
rect 3256 8730 3312 8732
rect 3016 8678 3062 8730
rect 3062 8678 3072 8730
rect 3096 8678 3126 8730
rect 3126 8678 3138 8730
rect 3138 8678 3152 8730
rect 3176 8678 3190 8730
rect 3190 8678 3202 8730
rect 3202 8678 3232 8730
rect 3256 8678 3266 8730
rect 3266 8678 3312 8730
rect 3016 8676 3072 8678
rect 3096 8676 3152 8678
rect 3176 8676 3232 8678
rect 3256 8676 3312 8678
rect 2870 8608 2926 8664
rect 4802 9288 4858 9344
rect 1582 8492 1638 8528
rect 1582 8472 1584 8492
rect 1584 8472 1636 8492
rect 1636 8472 1638 8492
rect 2870 8336 2926 8392
rect 1956 8186 2012 8188
rect 2036 8186 2092 8188
rect 2116 8186 2172 8188
rect 2196 8186 2252 8188
rect 1956 8134 2002 8186
rect 2002 8134 2012 8186
rect 2036 8134 2066 8186
rect 2066 8134 2078 8186
rect 2078 8134 2092 8186
rect 2116 8134 2130 8186
rect 2130 8134 2142 8186
rect 2142 8134 2172 8186
rect 2196 8134 2206 8186
rect 2206 8134 2252 8186
rect 1956 8132 2012 8134
rect 2036 8132 2092 8134
rect 2116 8132 2172 8134
rect 2196 8132 2252 8134
rect 3016 7642 3072 7644
rect 3096 7642 3152 7644
rect 3176 7642 3232 7644
rect 3256 7642 3312 7644
rect 3016 7590 3062 7642
rect 3062 7590 3072 7642
rect 3096 7590 3126 7642
rect 3126 7590 3138 7642
rect 3138 7590 3152 7642
rect 3176 7590 3190 7642
rect 3190 7590 3202 7642
rect 3202 7590 3232 7642
rect 3256 7590 3266 7642
rect 3266 7590 3312 7642
rect 3016 7588 3072 7590
rect 3096 7588 3152 7590
rect 3176 7588 3232 7590
rect 3256 7588 3312 7590
rect 7378 8880 7434 8936
rect 6826 7792 6882 7848
rect 1956 7098 2012 7100
rect 2036 7098 2092 7100
rect 2116 7098 2172 7100
rect 2196 7098 2252 7100
rect 1956 7046 2002 7098
rect 2002 7046 2012 7098
rect 2036 7046 2066 7098
rect 2066 7046 2078 7098
rect 2078 7046 2092 7098
rect 2116 7046 2130 7098
rect 2130 7046 2142 7098
rect 2142 7046 2172 7098
rect 2196 7046 2206 7098
rect 2206 7046 2252 7098
rect 1956 7044 2012 7046
rect 2036 7044 2092 7046
rect 2116 7044 2172 7046
rect 2196 7044 2252 7046
rect 5538 7248 5594 7304
rect 5906 7268 5962 7304
rect 5906 7248 5908 7268
rect 5908 7248 5960 7268
rect 5960 7248 5962 7268
rect 3016 6554 3072 6556
rect 3096 6554 3152 6556
rect 3176 6554 3232 6556
rect 3256 6554 3312 6556
rect 3016 6502 3062 6554
rect 3062 6502 3072 6554
rect 3096 6502 3126 6554
rect 3126 6502 3138 6554
rect 3138 6502 3152 6554
rect 3176 6502 3190 6554
rect 3190 6502 3202 6554
rect 3202 6502 3232 6554
rect 3256 6502 3266 6554
rect 3266 6502 3312 6554
rect 3016 6500 3072 6502
rect 3096 6500 3152 6502
rect 3176 6500 3232 6502
rect 3256 6500 3312 6502
rect 1956 6010 2012 6012
rect 2036 6010 2092 6012
rect 2116 6010 2172 6012
rect 2196 6010 2252 6012
rect 1956 5958 2002 6010
rect 2002 5958 2012 6010
rect 2036 5958 2066 6010
rect 2066 5958 2078 6010
rect 2078 5958 2092 6010
rect 2116 5958 2130 6010
rect 2130 5958 2142 6010
rect 2142 5958 2172 6010
rect 2196 5958 2206 6010
rect 2206 5958 2252 6010
rect 1956 5956 2012 5958
rect 2036 5956 2092 5958
rect 2116 5956 2172 5958
rect 2196 5956 2252 5958
rect 3016 5466 3072 5468
rect 3096 5466 3152 5468
rect 3176 5466 3232 5468
rect 3256 5466 3312 5468
rect 3016 5414 3062 5466
rect 3062 5414 3072 5466
rect 3096 5414 3126 5466
rect 3126 5414 3138 5466
rect 3138 5414 3152 5466
rect 3176 5414 3190 5466
rect 3190 5414 3202 5466
rect 3202 5414 3232 5466
rect 3256 5414 3266 5466
rect 3266 5414 3312 5466
rect 3016 5412 3072 5414
rect 3096 5412 3152 5414
rect 3176 5412 3232 5414
rect 3256 5412 3312 5414
rect 1956 4922 2012 4924
rect 2036 4922 2092 4924
rect 2116 4922 2172 4924
rect 2196 4922 2252 4924
rect 1956 4870 2002 4922
rect 2002 4870 2012 4922
rect 2036 4870 2066 4922
rect 2066 4870 2078 4922
rect 2078 4870 2092 4922
rect 2116 4870 2130 4922
rect 2130 4870 2142 4922
rect 2142 4870 2172 4922
rect 2196 4870 2206 4922
rect 2206 4870 2252 4922
rect 1956 4868 2012 4870
rect 2036 4868 2092 4870
rect 2116 4868 2172 4870
rect 2196 4868 2252 4870
rect 3016 4378 3072 4380
rect 3096 4378 3152 4380
rect 3176 4378 3232 4380
rect 3256 4378 3312 4380
rect 3016 4326 3062 4378
rect 3062 4326 3072 4378
rect 3096 4326 3126 4378
rect 3126 4326 3138 4378
rect 3138 4326 3152 4378
rect 3176 4326 3190 4378
rect 3190 4326 3202 4378
rect 3202 4326 3232 4378
rect 3256 4326 3266 4378
rect 3266 4326 3312 4378
rect 3016 4324 3072 4326
rect 3096 4324 3152 4326
rect 3176 4324 3232 4326
rect 3256 4324 3312 4326
rect 1956 3834 2012 3836
rect 2036 3834 2092 3836
rect 2116 3834 2172 3836
rect 2196 3834 2252 3836
rect 1956 3782 2002 3834
rect 2002 3782 2012 3834
rect 2036 3782 2066 3834
rect 2066 3782 2078 3834
rect 2078 3782 2092 3834
rect 2116 3782 2130 3834
rect 2130 3782 2142 3834
rect 2142 3782 2172 3834
rect 2196 3782 2206 3834
rect 2206 3782 2252 3834
rect 1956 3780 2012 3782
rect 2036 3780 2092 3782
rect 2116 3780 2172 3782
rect 2196 3780 2252 3782
rect 3016 3290 3072 3292
rect 3096 3290 3152 3292
rect 3176 3290 3232 3292
rect 3256 3290 3312 3292
rect 3016 3238 3062 3290
rect 3062 3238 3072 3290
rect 3096 3238 3126 3290
rect 3126 3238 3138 3290
rect 3138 3238 3152 3290
rect 3176 3238 3190 3290
rect 3190 3238 3202 3290
rect 3202 3238 3232 3290
rect 3256 3238 3266 3290
rect 3266 3238 3312 3290
rect 3016 3236 3072 3238
rect 3096 3236 3152 3238
rect 3176 3236 3232 3238
rect 3256 3236 3312 3238
rect 1956 2746 2012 2748
rect 2036 2746 2092 2748
rect 2116 2746 2172 2748
rect 2196 2746 2252 2748
rect 1956 2694 2002 2746
rect 2002 2694 2012 2746
rect 2036 2694 2066 2746
rect 2066 2694 2078 2746
rect 2078 2694 2092 2746
rect 2116 2694 2130 2746
rect 2130 2694 2142 2746
rect 2142 2694 2172 2746
rect 2196 2694 2206 2746
rect 2206 2694 2252 2746
rect 1956 2692 2012 2694
rect 2036 2692 2092 2694
rect 2116 2692 2172 2694
rect 2196 2692 2252 2694
rect 2870 2216 2926 2272
rect 3016 2202 3072 2204
rect 3096 2202 3152 2204
rect 3176 2202 3232 2204
rect 3256 2202 3312 2204
rect 3016 2150 3062 2202
rect 3062 2150 3072 2202
rect 3096 2150 3126 2202
rect 3126 2150 3138 2202
rect 3138 2150 3152 2202
rect 3176 2150 3190 2202
rect 3190 2150 3202 2202
rect 3202 2150 3232 2202
rect 3256 2150 3266 2202
rect 3266 2150 3312 2202
rect 3016 2148 3072 2150
rect 3096 2148 3152 2150
rect 3176 2148 3232 2150
rect 3256 2148 3312 2150
rect 2870 1808 2926 1864
rect 5538 6296 5594 6352
rect 7746 9560 7802 9616
rect 7654 8200 7710 8256
rect 9016 8730 9072 8732
rect 9096 8730 9152 8732
rect 9176 8730 9232 8732
rect 9256 8730 9312 8732
rect 9016 8678 9062 8730
rect 9062 8678 9072 8730
rect 9096 8678 9126 8730
rect 9126 8678 9138 8730
rect 9138 8678 9152 8730
rect 9176 8678 9190 8730
rect 9190 8678 9202 8730
rect 9202 8678 9232 8730
rect 9256 8678 9266 8730
rect 9266 8678 9312 8730
rect 9016 8676 9072 8678
rect 9096 8676 9152 8678
rect 9176 8676 9232 8678
rect 9256 8676 9312 8678
rect 12438 9016 12494 9072
rect 7956 8186 8012 8188
rect 8036 8186 8092 8188
rect 8116 8186 8172 8188
rect 8196 8186 8252 8188
rect 7956 8134 8002 8186
rect 8002 8134 8012 8186
rect 8036 8134 8066 8186
rect 8066 8134 8078 8186
rect 8078 8134 8092 8186
rect 8116 8134 8130 8186
rect 8130 8134 8142 8186
rect 8142 8134 8172 8186
rect 8196 8134 8206 8186
rect 8206 8134 8252 8186
rect 7956 8132 8012 8134
rect 8036 8132 8092 8134
rect 8116 8132 8172 8134
rect 8196 8132 8252 8134
rect 9016 7642 9072 7644
rect 9096 7642 9152 7644
rect 9176 7642 9232 7644
rect 9256 7642 9312 7644
rect 9016 7590 9062 7642
rect 9062 7590 9072 7642
rect 9096 7590 9126 7642
rect 9126 7590 9138 7642
rect 9138 7590 9152 7642
rect 9176 7590 9190 7642
rect 9190 7590 9202 7642
rect 9202 7590 9232 7642
rect 9256 7590 9266 7642
rect 9266 7590 9312 7642
rect 9016 7588 9072 7590
rect 9096 7588 9152 7590
rect 9176 7588 9232 7590
rect 9256 7588 9312 7590
rect 13956 8186 14012 8188
rect 14036 8186 14092 8188
rect 14116 8186 14172 8188
rect 14196 8186 14252 8188
rect 13956 8134 14002 8186
rect 14002 8134 14012 8186
rect 14036 8134 14066 8186
rect 14066 8134 14078 8186
rect 14078 8134 14092 8186
rect 14116 8134 14130 8186
rect 14130 8134 14142 8186
rect 14142 8134 14172 8186
rect 14196 8134 14206 8186
rect 14206 8134 14252 8186
rect 13956 8132 14012 8134
rect 14036 8132 14092 8134
rect 14116 8132 14172 8134
rect 14196 8132 14252 8134
rect 15016 8730 15072 8732
rect 15096 8730 15152 8732
rect 15176 8730 15232 8732
rect 15256 8730 15312 8732
rect 15016 8678 15062 8730
rect 15062 8678 15072 8730
rect 15096 8678 15126 8730
rect 15126 8678 15138 8730
rect 15138 8678 15152 8730
rect 15176 8678 15190 8730
rect 15190 8678 15202 8730
rect 15202 8678 15232 8730
rect 15256 8678 15266 8730
rect 15266 8678 15312 8730
rect 15016 8676 15072 8678
rect 15096 8676 15152 8678
rect 15176 8676 15232 8678
rect 15256 8676 15312 8678
rect 17130 9832 17186 9888
rect 15106 8336 15162 8392
rect 6274 6840 6330 6896
rect 7956 7098 8012 7100
rect 8036 7098 8092 7100
rect 8116 7098 8172 7100
rect 8196 7098 8252 7100
rect 7956 7046 8002 7098
rect 8002 7046 8012 7098
rect 8036 7046 8066 7098
rect 8066 7046 8078 7098
rect 8078 7046 8092 7098
rect 8116 7046 8130 7098
rect 8130 7046 8142 7098
rect 8142 7046 8172 7098
rect 8196 7046 8206 7098
rect 8206 7046 8252 7098
rect 7956 7044 8012 7046
rect 8036 7044 8092 7046
rect 8116 7044 8172 7046
rect 8196 7044 8252 7046
rect 7956 6010 8012 6012
rect 8036 6010 8092 6012
rect 8116 6010 8172 6012
rect 8196 6010 8252 6012
rect 7956 5958 8002 6010
rect 8002 5958 8012 6010
rect 8036 5958 8066 6010
rect 8066 5958 8078 6010
rect 8078 5958 8092 6010
rect 8116 5958 8130 6010
rect 8130 5958 8142 6010
rect 8142 5958 8172 6010
rect 8196 5958 8206 6010
rect 8206 5958 8252 6010
rect 7956 5956 8012 5958
rect 8036 5956 8092 5958
rect 8116 5956 8172 5958
rect 8196 5956 8252 5958
rect 7956 4922 8012 4924
rect 8036 4922 8092 4924
rect 8116 4922 8172 4924
rect 8196 4922 8252 4924
rect 7956 4870 8002 4922
rect 8002 4870 8012 4922
rect 8036 4870 8066 4922
rect 8066 4870 8078 4922
rect 8078 4870 8092 4922
rect 8116 4870 8130 4922
rect 8130 4870 8142 4922
rect 8142 4870 8172 4922
rect 8196 4870 8206 4922
rect 8206 4870 8252 4922
rect 7956 4868 8012 4870
rect 8036 4868 8092 4870
rect 8116 4868 8172 4870
rect 8196 4868 8252 4870
rect 7956 3834 8012 3836
rect 8036 3834 8092 3836
rect 8116 3834 8172 3836
rect 8196 3834 8252 3836
rect 7956 3782 8002 3834
rect 8002 3782 8012 3834
rect 8036 3782 8066 3834
rect 8066 3782 8078 3834
rect 8078 3782 8092 3834
rect 8116 3782 8130 3834
rect 8130 3782 8142 3834
rect 8142 3782 8172 3834
rect 8196 3782 8206 3834
rect 8206 3782 8252 3834
rect 7956 3780 8012 3782
rect 8036 3780 8092 3782
rect 8116 3780 8172 3782
rect 8196 3780 8252 3782
rect 7956 2746 8012 2748
rect 8036 2746 8092 2748
rect 8116 2746 8172 2748
rect 8196 2746 8252 2748
rect 7956 2694 8002 2746
rect 8002 2694 8012 2746
rect 8036 2694 8066 2746
rect 8066 2694 8078 2746
rect 8078 2694 8092 2746
rect 8116 2694 8130 2746
rect 8130 2694 8142 2746
rect 8142 2694 8172 2746
rect 8196 2694 8206 2746
rect 8206 2694 8252 2746
rect 7956 2692 8012 2694
rect 8036 2692 8092 2694
rect 8116 2692 8172 2694
rect 8196 2692 8252 2694
rect 10966 6704 11022 6760
rect 9016 6554 9072 6556
rect 9096 6554 9152 6556
rect 9176 6554 9232 6556
rect 9256 6554 9312 6556
rect 9016 6502 9062 6554
rect 9062 6502 9072 6554
rect 9096 6502 9126 6554
rect 9126 6502 9138 6554
rect 9138 6502 9152 6554
rect 9176 6502 9190 6554
rect 9190 6502 9202 6554
rect 9202 6502 9232 6554
rect 9256 6502 9266 6554
rect 9266 6502 9312 6554
rect 9016 6500 9072 6502
rect 9096 6500 9152 6502
rect 9176 6500 9232 6502
rect 9256 6500 9312 6502
rect 9016 5466 9072 5468
rect 9096 5466 9152 5468
rect 9176 5466 9232 5468
rect 9256 5466 9312 5468
rect 9016 5414 9062 5466
rect 9062 5414 9072 5466
rect 9096 5414 9126 5466
rect 9126 5414 9138 5466
rect 9138 5414 9152 5466
rect 9176 5414 9190 5466
rect 9190 5414 9202 5466
rect 9202 5414 9232 5466
rect 9256 5414 9266 5466
rect 9266 5414 9312 5466
rect 9016 5412 9072 5414
rect 9096 5412 9152 5414
rect 9176 5412 9232 5414
rect 9256 5412 9312 5414
rect 9016 4378 9072 4380
rect 9096 4378 9152 4380
rect 9176 4378 9232 4380
rect 9256 4378 9312 4380
rect 9016 4326 9062 4378
rect 9062 4326 9072 4378
rect 9096 4326 9126 4378
rect 9126 4326 9138 4378
rect 9138 4326 9152 4378
rect 9176 4326 9190 4378
rect 9190 4326 9202 4378
rect 9202 4326 9232 4378
rect 9256 4326 9266 4378
rect 9266 4326 9312 4378
rect 9016 4324 9072 4326
rect 9096 4324 9152 4326
rect 9176 4324 9232 4326
rect 9256 4324 9312 4326
rect 9016 3290 9072 3292
rect 9096 3290 9152 3292
rect 9176 3290 9232 3292
rect 9256 3290 9312 3292
rect 9016 3238 9062 3290
rect 9062 3238 9072 3290
rect 9096 3238 9126 3290
rect 9126 3238 9138 3290
rect 9138 3238 9152 3290
rect 9176 3238 9190 3290
rect 9190 3238 9202 3290
rect 9202 3238 9232 3290
rect 9256 3238 9266 3290
rect 9266 3238 9312 3290
rect 9016 3236 9072 3238
rect 9096 3236 9152 3238
rect 9176 3236 9232 3238
rect 9256 3236 9312 3238
rect 9016 2202 9072 2204
rect 9096 2202 9152 2204
rect 9176 2202 9232 2204
rect 9256 2202 9312 2204
rect 9016 2150 9062 2202
rect 9062 2150 9072 2202
rect 9096 2150 9126 2202
rect 9126 2150 9138 2202
rect 9138 2150 9152 2202
rect 9176 2150 9190 2202
rect 9190 2150 9202 2202
rect 9202 2150 9232 2202
rect 9256 2150 9266 2202
rect 9266 2150 9312 2202
rect 9016 2148 9072 2150
rect 9096 2148 9152 2150
rect 9176 2148 9232 2150
rect 9256 2148 9312 2150
rect 12714 5480 12770 5536
rect 11886 5208 11942 5264
rect 10782 2352 10838 2408
rect 10506 1264 10562 1320
rect 10230 1128 10286 1184
rect 12530 3984 12586 4040
rect 13082 3576 13138 3632
rect 13910 7420 13912 7440
rect 13912 7420 13964 7440
rect 13964 7420 13966 7440
rect 13910 7384 13966 7420
rect 14554 7928 14610 7984
rect 13956 7098 14012 7100
rect 14036 7098 14092 7100
rect 14116 7098 14172 7100
rect 14196 7098 14252 7100
rect 13956 7046 14002 7098
rect 14002 7046 14012 7098
rect 14036 7046 14066 7098
rect 14066 7046 14078 7098
rect 14078 7046 14092 7098
rect 14116 7046 14130 7098
rect 14130 7046 14142 7098
rect 14142 7046 14172 7098
rect 14196 7046 14206 7098
rect 14206 7046 14252 7098
rect 13956 7044 14012 7046
rect 14036 7044 14092 7046
rect 14116 7044 14172 7046
rect 14196 7044 14252 7046
rect 15016 7642 15072 7644
rect 15096 7642 15152 7644
rect 15176 7642 15232 7644
rect 15256 7642 15312 7644
rect 15016 7590 15062 7642
rect 15062 7590 15072 7642
rect 15096 7590 15126 7642
rect 15126 7590 15138 7642
rect 15138 7590 15152 7642
rect 15176 7590 15190 7642
rect 15190 7590 15202 7642
rect 15202 7590 15232 7642
rect 15256 7590 15266 7642
rect 15266 7590 15312 7642
rect 15016 7588 15072 7590
rect 15096 7588 15152 7590
rect 15176 7588 15232 7590
rect 15256 7588 15312 7590
rect 15016 6554 15072 6556
rect 15096 6554 15152 6556
rect 15176 6554 15232 6556
rect 15256 6554 15312 6556
rect 15016 6502 15062 6554
rect 15062 6502 15072 6554
rect 15096 6502 15126 6554
rect 15126 6502 15138 6554
rect 15138 6502 15152 6554
rect 15176 6502 15190 6554
rect 15190 6502 15202 6554
rect 15202 6502 15232 6554
rect 15256 6502 15266 6554
rect 15266 6502 15312 6554
rect 15016 6500 15072 6502
rect 15096 6500 15152 6502
rect 15176 6500 15232 6502
rect 15256 6500 15312 6502
rect 13956 6010 14012 6012
rect 14036 6010 14092 6012
rect 14116 6010 14172 6012
rect 14196 6010 14252 6012
rect 13956 5958 14002 6010
rect 14002 5958 14012 6010
rect 14036 5958 14066 6010
rect 14066 5958 14078 6010
rect 14078 5958 14092 6010
rect 14116 5958 14130 6010
rect 14130 5958 14142 6010
rect 14142 5958 14172 6010
rect 14196 5958 14206 6010
rect 14206 5958 14252 6010
rect 13956 5956 14012 5958
rect 14036 5956 14092 5958
rect 14116 5956 14172 5958
rect 14196 5956 14252 5958
rect 13726 5752 13782 5808
rect 13956 4922 14012 4924
rect 14036 4922 14092 4924
rect 14116 4922 14172 4924
rect 14196 4922 14252 4924
rect 13956 4870 14002 4922
rect 14002 4870 14012 4922
rect 14036 4870 14066 4922
rect 14066 4870 14078 4922
rect 14078 4870 14092 4922
rect 14116 4870 14130 4922
rect 14130 4870 14142 4922
rect 14142 4870 14172 4922
rect 14196 4870 14206 4922
rect 14206 4870 14252 4922
rect 13956 4868 14012 4870
rect 14036 4868 14092 4870
rect 14116 4868 14172 4870
rect 14196 4868 14252 4870
rect 13956 3834 14012 3836
rect 14036 3834 14092 3836
rect 14116 3834 14172 3836
rect 14196 3834 14252 3836
rect 13956 3782 14002 3834
rect 14002 3782 14012 3834
rect 14036 3782 14066 3834
rect 14066 3782 14078 3834
rect 14078 3782 14092 3834
rect 14116 3782 14130 3834
rect 14130 3782 14142 3834
rect 14142 3782 14172 3834
rect 14196 3782 14206 3834
rect 14206 3782 14252 3834
rect 13956 3780 14012 3782
rect 14036 3780 14092 3782
rect 14116 3780 14172 3782
rect 14196 3780 14252 3782
rect 13956 2746 14012 2748
rect 14036 2746 14092 2748
rect 14116 2746 14172 2748
rect 14196 2746 14252 2748
rect 13956 2694 14002 2746
rect 14002 2694 14012 2746
rect 14036 2694 14066 2746
rect 14066 2694 14078 2746
rect 14078 2694 14092 2746
rect 14116 2694 14130 2746
rect 14130 2694 14142 2746
rect 14142 2694 14172 2746
rect 14196 2694 14206 2746
rect 14206 2694 14252 2746
rect 13956 2692 14012 2694
rect 14036 2692 14092 2694
rect 14116 2692 14172 2694
rect 14196 2692 14252 2694
rect 15016 5466 15072 5468
rect 15096 5466 15152 5468
rect 15176 5466 15232 5468
rect 15256 5466 15312 5468
rect 15016 5414 15062 5466
rect 15062 5414 15072 5466
rect 15096 5414 15126 5466
rect 15126 5414 15138 5466
rect 15138 5414 15152 5466
rect 15176 5414 15190 5466
rect 15190 5414 15202 5466
rect 15202 5414 15232 5466
rect 15256 5414 15266 5466
rect 15266 5414 15312 5466
rect 15016 5412 15072 5414
rect 15096 5412 15152 5414
rect 15176 5412 15232 5414
rect 15256 5412 15312 5414
rect 15016 4378 15072 4380
rect 15096 4378 15152 4380
rect 15176 4378 15232 4380
rect 15256 4378 15312 4380
rect 15016 4326 15062 4378
rect 15062 4326 15072 4378
rect 15096 4326 15126 4378
rect 15126 4326 15138 4378
rect 15138 4326 15152 4378
rect 15176 4326 15190 4378
rect 15190 4326 15202 4378
rect 15202 4326 15232 4378
rect 15256 4326 15266 4378
rect 15266 4326 15312 4378
rect 15016 4324 15072 4326
rect 15096 4324 15152 4326
rect 15176 4324 15232 4326
rect 15256 4324 15312 4326
rect 15016 3290 15072 3292
rect 15096 3290 15152 3292
rect 15176 3290 15232 3292
rect 15256 3290 15312 3292
rect 15016 3238 15062 3290
rect 15062 3238 15072 3290
rect 15096 3238 15126 3290
rect 15126 3238 15138 3290
rect 15138 3238 15152 3290
rect 15176 3238 15190 3290
rect 15190 3238 15202 3290
rect 15202 3238 15232 3290
rect 15256 3238 15266 3290
rect 15266 3238 15312 3290
rect 15016 3236 15072 3238
rect 15096 3236 15152 3238
rect 15176 3236 15232 3238
rect 15256 3236 15312 3238
rect 15016 2202 15072 2204
rect 15096 2202 15152 2204
rect 15176 2202 15232 2204
rect 15256 2202 15312 2204
rect 15016 2150 15062 2202
rect 15062 2150 15072 2202
rect 15096 2150 15126 2202
rect 15126 2150 15138 2202
rect 15138 2150 15152 2202
rect 15176 2150 15190 2202
rect 15190 2150 15202 2202
rect 15202 2150 15232 2202
rect 15256 2150 15266 2202
rect 15266 2150 15312 2202
rect 15016 2148 15072 2150
rect 15096 2148 15152 2150
rect 15176 2148 15232 2150
rect 15256 2148 15312 2150
rect 16486 6160 16542 6216
rect 21016 8730 21072 8732
rect 21096 8730 21152 8732
rect 21176 8730 21232 8732
rect 21256 8730 21312 8732
rect 21016 8678 21062 8730
rect 21062 8678 21072 8730
rect 21096 8678 21126 8730
rect 21126 8678 21138 8730
rect 21138 8678 21152 8730
rect 21176 8678 21190 8730
rect 21190 8678 21202 8730
rect 21202 8678 21232 8730
rect 21256 8678 21266 8730
rect 21266 8678 21312 8730
rect 21016 8676 21072 8678
rect 21096 8676 21152 8678
rect 21176 8676 21232 8678
rect 21256 8676 21312 8678
rect 19956 8186 20012 8188
rect 20036 8186 20092 8188
rect 20116 8186 20172 8188
rect 20196 8186 20252 8188
rect 19956 8134 20002 8186
rect 20002 8134 20012 8186
rect 20036 8134 20066 8186
rect 20066 8134 20078 8186
rect 20078 8134 20092 8186
rect 20116 8134 20130 8186
rect 20130 8134 20142 8186
rect 20142 8134 20172 8186
rect 20196 8134 20206 8186
rect 20206 8134 20252 8186
rect 19956 8132 20012 8134
rect 20036 8132 20092 8134
rect 20116 8132 20172 8134
rect 20196 8132 20252 8134
rect 16946 5072 17002 5128
rect 17130 2352 17186 2408
rect 17314 1400 17370 1456
rect 19338 4664 19394 4720
rect 18050 1264 18106 1320
rect 18970 2488 19026 2544
rect 18694 1128 18750 1184
rect 19956 7098 20012 7100
rect 20036 7098 20092 7100
rect 20116 7098 20172 7100
rect 20196 7098 20252 7100
rect 19956 7046 20002 7098
rect 20002 7046 20012 7098
rect 20036 7046 20066 7098
rect 20066 7046 20078 7098
rect 20078 7046 20092 7098
rect 20116 7046 20130 7098
rect 20130 7046 20142 7098
rect 20142 7046 20172 7098
rect 20196 7046 20206 7098
rect 20206 7046 20252 7098
rect 19956 7044 20012 7046
rect 20036 7044 20092 7046
rect 20116 7044 20172 7046
rect 20196 7044 20252 7046
rect 19956 6010 20012 6012
rect 20036 6010 20092 6012
rect 20116 6010 20172 6012
rect 20196 6010 20252 6012
rect 19956 5958 20002 6010
rect 20002 5958 20012 6010
rect 20036 5958 20066 6010
rect 20066 5958 20078 6010
rect 20078 5958 20092 6010
rect 20116 5958 20130 6010
rect 20130 5958 20142 6010
rect 20142 5958 20172 6010
rect 20196 5958 20206 6010
rect 20206 5958 20252 6010
rect 19956 5956 20012 5958
rect 20036 5956 20092 5958
rect 20116 5956 20172 5958
rect 20196 5956 20252 5958
rect 21016 7642 21072 7644
rect 21096 7642 21152 7644
rect 21176 7642 21232 7644
rect 21256 7642 21312 7644
rect 21016 7590 21062 7642
rect 21062 7590 21072 7642
rect 21096 7590 21126 7642
rect 21126 7590 21138 7642
rect 21138 7590 21152 7642
rect 21176 7590 21190 7642
rect 21190 7590 21202 7642
rect 21202 7590 21232 7642
rect 21256 7590 21266 7642
rect 21266 7590 21312 7642
rect 21016 7588 21072 7590
rect 21096 7588 21152 7590
rect 21176 7588 21232 7590
rect 21256 7588 21312 7590
rect 21016 6554 21072 6556
rect 21096 6554 21152 6556
rect 21176 6554 21232 6556
rect 21256 6554 21312 6556
rect 21016 6502 21062 6554
rect 21062 6502 21072 6554
rect 21096 6502 21126 6554
rect 21126 6502 21138 6554
rect 21138 6502 21152 6554
rect 21176 6502 21190 6554
rect 21190 6502 21202 6554
rect 21202 6502 21232 6554
rect 21256 6502 21266 6554
rect 21266 6502 21312 6554
rect 21016 6500 21072 6502
rect 21096 6500 21152 6502
rect 21176 6500 21232 6502
rect 21256 6500 21312 6502
rect 19956 4922 20012 4924
rect 20036 4922 20092 4924
rect 20116 4922 20172 4924
rect 20196 4922 20252 4924
rect 19956 4870 20002 4922
rect 20002 4870 20012 4922
rect 20036 4870 20066 4922
rect 20066 4870 20078 4922
rect 20078 4870 20092 4922
rect 20116 4870 20130 4922
rect 20130 4870 20142 4922
rect 20142 4870 20172 4922
rect 20196 4870 20206 4922
rect 20206 4870 20252 4922
rect 19956 4868 20012 4870
rect 20036 4868 20092 4870
rect 20116 4868 20172 4870
rect 20196 4868 20252 4870
rect 21016 5466 21072 5468
rect 21096 5466 21152 5468
rect 21176 5466 21232 5468
rect 21256 5466 21312 5468
rect 21016 5414 21062 5466
rect 21062 5414 21072 5466
rect 21096 5414 21126 5466
rect 21126 5414 21138 5466
rect 21138 5414 21152 5466
rect 21176 5414 21190 5466
rect 21190 5414 21202 5466
rect 21202 5414 21232 5466
rect 21256 5414 21266 5466
rect 21266 5414 21312 5466
rect 21016 5412 21072 5414
rect 21096 5412 21152 5414
rect 21176 5412 21232 5414
rect 21256 5412 21312 5414
rect 20902 4528 20958 4584
rect 19798 3984 19854 4040
rect 19956 3834 20012 3836
rect 20036 3834 20092 3836
rect 20116 3834 20172 3836
rect 20196 3834 20252 3836
rect 19956 3782 20002 3834
rect 20002 3782 20012 3834
rect 20036 3782 20066 3834
rect 20066 3782 20078 3834
rect 20078 3782 20092 3834
rect 20116 3782 20130 3834
rect 20130 3782 20142 3834
rect 20142 3782 20172 3834
rect 20196 3782 20206 3834
rect 20206 3782 20252 3834
rect 19956 3780 20012 3782
rect 20036 3780 20092 3782
rect 20116 3780 20172 3782
rect 20196 3780 20252 3782
rect 21016 4378 21072 4380
rect 21096 4378 21152 4380
rect 21176 4378 21232 4380
rect 21256 4378 21312 4380
rect 21016 4326 21062 4378
rect 21062 4326 21072 4378
rect 21096 4326 21126 4378
rect 21126 4326 21138 4378
rect 21138 4326 21152 4378
rect 21176 4326 21190 4378
rect 21190 4326 21202 4378
rect 21202 4326 21232 4378
rect 21256 4326 21266 4378
rect 21266 4326 21312 4378
rect 21016 4324 21072 4326
rect 21096 4324 21152 4326
rect 21176 4324 21232 4326
rect 21256 4324 21312 4326
rect 19706 2352 19762 2408
rect 19956 2746 20012 2748
rect 20036 2746 20092 2748
rect 20116 2746 20172 2748
rect 20196 2746 20252 2748
rect 19956 2694 20002 2746
rect 20002 2694 20012 2746
rect 20036 2694 20066 2746
rect 20066 2694 20078 2746
rect 20078 2694 20092 2746
rect 20116 2694 20130 2746
rect 20130 2694 20142 2746
rect 20142 2694 20172 2746
rect 20196 2694 20206 2746
rect 20206 2694 20252 2746
rect 19956 2692 20012 2694
rect 20036 2692 20092 2694
rect 20116 2692 20172 2694
rect 20196 2692 20252 2694
rect 20074 1672 20130 1728
rect 20534 2372 20590 2408
rect 20534 2352 20536 2372
rect 20536 2352 20588 2372
rect 20588 2352 20590 2372
rect 21016 3290 21072 3292
rect 21096 3290 21152 3292
rect 21176 3290 21232 3292
rect 21256 3290 21312 3292
rect 21016 3238 21062 3290
rect 21062 3238 21072 3290
rect 21096 3238 21126 3290
rect 21126 3238 21138 3290
rect 21138 3238 21152 3290
rect 21176 3238 21190 3290
rect 21190 3238 21202 3290
rect 21202 3238 21232 3290
rect 21256 3238 21266 3290
rect 21266 3238 21312 3290
rect 21016 3236 21072 3238
rect 21096 3236 21152 3238
rect 21176 3236 21232 3238
rect 21256 3236 21312 3238
rect 20718 1808 20774 1864
rect 21016 2202 21072 2204
rect 21096 2202 21152 2204
rect 21176 2202 21232 2204
rect 21256 2202 21312 2204
rect 21016 2150 21062 2202
rect 21062 2150 21072 2202
rect 21096 2150 21126 2202
rect 21126 2150 21138 2202
rect 21138 2150 21152 2202
rect 21176 2150 21190 2202
rect 21190 2150 21202 2202
rect 21202 2150 21232 2202
rect 21256 2150 21266 2202
rect 21266 2150 21312 2202
rect 21016 2148 21072 2150
rect 21096 2148 21152 2150
rect 21176 2148 21232 2150
rect 21256 2148 21312 2150
rect 21638 2624 21694 2680
rect 21730 1944 21786 2000
rect 23018 4120 23074 4176
rect 25134 8472 25190 8528
rect 27016 8730 27072 8732
rect 27096 8730 27152 8732
rect 27176 8730 27232 8732
rect 27256 8730 27312 8732
rect 27016 8678 27062 8730
rect 27062 8678 27072 8730
rect 27096 8678 27126 8730
rect 27126 8678 27138 8730
rect 27138 8678 27152 8730
rect 27176 8678 27190 8730
rect 27190 8678 27202 8730
rect 27202 8678 27232 8730
rect 27256 8678 27266 8730
rect 27266 8678 27312 8730
rect 27016 8676 27072 8678
rect 27096 8676 27152 8678
rect 27176 8676 27232 8678
rect 27256 8676 27312 8678
rect 30102 9832 30158 9888
rect 30838 9560 30894 9616
rect 30470 9016 30526 9072
rect 25956 8186 26012 8188
rect 26036 8186 26092 8188
rect 26116 8186 26172 8188
rect 26196 8186 26252 8188
rect 25956 8134 26002 8186
rect 26002 8134 26012 8186
rect 26036 8134 26066 8186
rect 26066 8134 26078 8186
rect 26078 8134 26092 8186
rect 26116 8134 26130 8186
rect 26130 8134 26142 8186
rect 26142 8134 26172 8186
rect 26196 8134 26206 8186
rect 26206 8134 26252 8186
rect 25956 8132 26012 8134
rect 26036 8132 26092 8134
rect 26116 8132 26172 8134
rect 26196 8132 26252 8134
rect 24858 2624 24914 2680
rect 25226 3460 25282 3496
rect 25226 3440 25228 3460
rect 25228 3440 25280 3460
rect 25280 3440 25282 3460
rect 25778 3032 25834 3088
rect 25956 7098 26012 7100
rect 26036 7098 26092 7100
rect 26116 7098 26172 7100
rect 26196 7098 26252 7100
rect 25956 7046 26002 7098
rect 26002 7046 26012 7098
rect 26036 7046 26066 7098
rect 26066 7046 26078 7098
rect 26078 7046 26092 7098
rect 26116 7046 26130 7098
rect 26130 7046 26142 7098
rect 26142 7046 26172 7098
rect 26196 7046 26206 7098
rect 26206 7046 26252 7098
rect 25956 7044 26012 7046
rect 26036 7044 26092 7046
rect 26116 7044 26172 7046
rect 26196 7044 26252 7046
rect 25956 6010 26012 6012
rect 26036 6010 26092 6012
rect 26116 6010 26172 6012
rect 26196 6010 26252 6012
rect 25956 5958 26002 6010
rect 26002 5958 26012 6010
rect 26036 5958 26066 6010
rect 26066 5958 26078 6010
rect 26078 5958 26092 6010
rect 26116 5958 26130 6010
rect 26130 5958 26142 6010
rect 26142 5958 26172 6010
rect 26196 5958 26206 6010
rect 26206 5958 26252 6010
rect 25956 5956 26012 5958
rect 26036 5956 26092 5958
rect 26116 5956 26172 5958
rect 26196 5956 26252 5958
rect 25956 4922 26012 4924
rect 26036 4922 26092 4924
rect 26116 4922 26172 4924
rect 26196 4922 26252 4924
rect 25956 4870 26002 4922
rect 26002 4870 26012 4922
rect 26036 4870 26066 4922
rect 26066 4870 26078 4922
rect 26078 4870 26092 4922
rect 26116 4870 26130 4922
rect 26130 4870 26142 4922
rect 26142 4870 26172 4922
rect 26196 4870 26206 4922
rect 26206 4870 26252 4922
rect 25956 4868 26012 4870
rect 26036 4868 26092 4870
rect 26116 4868 26172 4870
rect 26196 4868 26252 4870
rect 25956 3834 26012 3836
rect 26036 3834 26092 3836
rect 26116 3834 26172 3836
rect 26196 3834 26252 3836
rect 25956 3782 26002 3834
rect 26002 3782 26012 3834
rect 26036 3782 26066 3834
rect 26066 3782 26078 3834
rect 26078 3782 26092 3834
rect 26116 3782 26130 3834
rect 26130 3782 26142 3834
rect 26142 3782 26172 3834
rect 26196 3782 26206 3834
rect 26206 3782 26252 3834
rect 25956 3780 26012 3782
rect 26036 3780 26092 3782
rect 26116 3780 26172 3782
rect 26196 3780 26252 3782
rect 26238 2896 26294 2952
rect 25956 2746 26012 2748
rect 26036 2746 26092 2748
rect 26116 2746 26172 2748
rect 26196 2746 26252 2748
rect 25956 2694 26002 2746
rect 26002 2694 26012 2746
rect 26036 2694 26066 2746
rect 26066 2694 26078 2746
rect 26078 2694 26092 2746
rect 26116 2694 26130 2746
rect 26130 2694 26142 2746
rect 26142 2694 26172 2746
rect 26196 2694 26206 2746
rect 26206 2694 26252 2746
rect 25956 2692 26012 2694
rect 26036 2692 26092 2694
rect 26116 2692 26172 2694
rect 26196 2692 26252 2694
rect 27016 7642 27072 7644
rect 27096 7642 27152 7644
rect 27176 7642 27232 7644
rect 27256 7642 27312 7644
rect 27016 7590 27062 7642
rect 27062 7590 27072 7642
rect 27096 7590 27126 7642
rect 27126 7590 27138 7642
rect 27138 7590 27152 7642
rect 27176 7590 27190 7642
rect 27190 7590 27202 7642
rect 27202 7590 27232 7642
rect 27256 7590 27266 7642
rect 27266 7590 27312 7642
rect 27016 7588 27072 7590
rect 27096 7588 27152 7590
rect 27176 7588 27232 7590
rect 27256 7588 27312 7590
rect 27016 6554 27072 6556
rect 27096 6554 27152 6556
rect 27176 6554 27232 6556
rect 27256 6554 27312 6556
rect 27016 6502 27062 6554
rect 27062 6502 27072 6554
rect 27096 6502 27126 6554
rect 27126 6502 27138 6554
rect 27138 6502 27152 6554
rect 27176 6502 27190 6554
rect 27190 6502 27202 6554
rect 27202 6502 27232 6554
rect 27256 6502 27266 6554
rect 27266 6502 27312 6554
rect 27016 6500 27072 6502
rect 27096 6500 27152 6502
rect 27176 6500 27232 6502
rect 27256 6500 27312 6502
rect 27016 5466 27072 5468
rect 27096 5466 27152 5468
rect 27176 5466 27232 5468
rect 27256 5466 27312 5468
rect 27016 5414 27062 5466
rect 27062 5414 27072 5466
rect 27096 5414 27126 5466
rect 27126 5414 27138 5466
rect 27138 5414 27152 5466
rect 27176 5414 27190 5466
rect 27190 5414 27202 5466
rect 27202 5414 27232 5466
rect 27256 5414 27266 5466
rect 27266 5414 27312 5466
rect 27016 5412 27072 5414
rect 27096 5412 27152 5414
rect 27176 5412 27232 5414
rect 27256 5412 27312 5414
rect 31482 9288 31538 9344
rect 31022 8744 31078 8800
rect 31390 8472 31446 8528
rect 32402 8200 32458 8256
rect 31956 8186 32012 8188
rect 32036 8186 32092 8188
rect 32116 8186 32172 8188
rect 32196 8186 32252 8188
rect 31956 8134 32002 8186
rect 32002 8134 32012 8186
rect 32036 8134 32066 8186
rect 32066 8134 32078 8186
rect 32078 8134 32092 8186
rect 32116 8134 32130 8186
rect 32130 8134 32142 8186
rect 32142 8134 32172 8186
rect 32196 8134 32206 8186
rect 32206 8134 32252 8186
rect 31956 8132 32012 8134
rect 32036 8132 32092 8134
rect 32116 8132 32172 8134
rect 32196 8132 32252 8134
rect 31850 7928 31906 7984
rect 32126 7692 32128 7712
rect 32128 7692 32180 7712
rect 32180 7692 32182 7712
rect 32126 7656 32182 7692
rect 31758 7384 31814 7440
rect 31298 7248 31354 7304
rect 31956 7098 32012 7100
rect 32036 7098 32092 7100
rect 32116 7098 32172 7100
rect 32196 7098 32252 7100
rect 31956 7046 32002 7098
rect 32002 7046 32012 7098
rect 32036 7046 32066 7098
rect 32066 7046 32078 7098
rect 32078 7046 32092 7098
rect 32116 7046 32130 7098
rect 32130 7046 32142 7098
rect 32142 7046 32172 7098
rect 32196 7046 32206 7098
rect 32206 7046 32252 7098
rect 31956 7044 32012 7046
rect 32036 7044 32092 7046
rect 32116 7044 32172 7046
rect 32196 7044 32252 7046
rect 32770 7148 32772 7168
rect 32772 7148 32824 7168
rect 32824 7148 32826 7168
rect 32770 7112 32826 7148
rect 31758 6840 31814 6896
rect 31390 6604 31392 6624
rect 31392 6604 31444 6624
rect 31444 6604 31446 6624
rect 31390 6568 31446 6604
rect 31482 6160 31538 6216
rect 27016 4378 27072 4380
rect 27096 4378 27152 4380
rect 27176 4378 27232 4380
rect 27256 4378 27312 4380
rect 27016 4326 27062 4378
rect 27062 4326 27072 4378
rect 27096 4326 27126 4378
rect 27126 4326 27138 4378
rect 27138 4326 27152 4378
rect 27176 4326 27190 4378
rect 27190 4326 27202 4378
rect 27202 4326 27232 4378
rect 27256 4326 27266 4378
rect 27266 4326 27312 4378
rect 27016 4324 27072 4326
rect 27096 4324 27152 4326
rect 27176 4324 27232 4326
rect 27256 4324 27312 4326
rect 27016 3290 27072 3292
rect 27096 3290 27152 3292
rect 27176 3290 27232 3292
rect 27256 3290 27312 3292
rect 27016 3238 27062 3290
rect 27062 3238 27072 3290
rect 27096 3238 27126 3290
rect 27126 3238 27138 3290
rect 27138 3238 27152 3290
rect 27176 3238 27190 3290
rect 27190 3238 27202 3290
rect 27202 3238 27232 3290
rect 27256 3238 27266 3290
rect 27266 3238 27312 3290
rect 27016 3236 27072 3238
rect 27096 3236 27152 3238
rect 27176 3236 27232 3238
rect 27256 3236 27312 3238
rect 27016 2202 27072 2204
rect 27096 2202 27152 2204
rect 27176 2202 27232 2204
rect 27256 2202 27312 2204
rect 27016 2150 27062 2202
rect 27062 2150 27072 2202
rect 27096 2150 27126 2202
rect 27126 2150 27138 2202
rect 27138 2150 27152 2202
rect 27176 2150 27190 2202
rect 27190 2150 27202 2202
rect 27202 2150 27232 2202
rect 27256 2150 27266 2202
rect 27266 2150 27312 2202
rect 27016 2148 27072 2150
rect 27096 2148 27152 2150
rect 27176 2148 27232 2150
rect 27256 2148 27312 2150
rect 28998 4020 29000 4040
rect 29000 4020 29052 4040
rect 29052 4020 29054 4040
rect 28998 3984 29054 4020
rect 31850 6296 31906 6352
rect 31758 5516 31760 5536
rect 31760 5516 31812 5536
rect 31812 5516 31814 5536
rect 31758 5480 31814 5516
rect 31482 4664 31538 4720
rect 31956 6010 32012 6012
rect 32036 6010 32092 6012
rect 32116 6010 32172 6012
rect 32196 6010 32252 6012
rect 31956 5958 32002 6010
rect 32002 5958 32012 6010
rect 32036 5958 32066 6010
rect 32066 5958 32078 6010
rect 32078 5958 32092 6010
rect 32116 5958 32130 6010
rect 32130 5958 32142 6010
rect 32142 5958 32172 6010
rect 32196 5958 32206 6010
rect 32206 5958 32252 6010
rect 31956 5956 32012 5958
rect 32036 5956 32092 5958
rect 32116 5956 32172 5958
rect 32196 5956 32252 5958
rect 32126 5788 32128 5808
rect 32128 5788 32180 5808
rect 32180 5788 32182 5808
rect 32126 5752 32182 5788
rect 32034 5208 32090 5264
rect 32862 4972 32864 4992
rect 32864 4972 32916 4992
rect 32916 4972 32918 4992
rect 32862 4936 32918 4972
rect 31956 4922 32012 4924
rect 32036 4922 32092 4924
rect 32116 4922 32172 4924
rect 32196 4922 32252 4924
rect 31956 4870 32002 4922
rect 32002 4870 32012 4922
rect 32036 4870 32066 4922
rect 32066 4870 32078 4922
rect 32078 4870 32092 4922
rect 32116 4870 32130 4922
rect 32130 4870 32142 4922
rect 32142 4870 32172 4922
rect 32196 4870 32206 4922
rect 32206 4870 32252 4922
rect 31956 4868 32012 4870
rect 32036 4868 32092 4870
rect 32116 4868 32172 4870
rect 32196 4868 32252 4870
rect 32126 4428 32128 4448
rect 32128 4428 32180 4448
rect 32180 4428 32182 4448
rect 32126 4392 32182 4428
rect 31758 4120 31814 4176
rect 32862 3884 32864 3904
rect 32864 3884 32916 3904
rect 32916 3884 32918 3904
rect 32862 3848 32918 3884
rect 31956 3834 32012 3836
rect 32036 3834 32092 3836
rect 32116 3834 32172 3836
rect 32196 3834 32252 3836
rect 31956 3782 32002 3834
rect 32002 3782 32012 3834
rect 32036 3782 32066 3834
rect 32066 3782 32078 3834
rect 32078 3782 32092 3834
rect 32116 3782 32130 3834
rect 32130 3782 32142 3834
rect 32142 3782 32172 3834
rect 32196 3782 32206 3834
rect 32206 3782 32252 3834
rect 31956 3780 32012 3782
rect 32036 3780 32092 3782
rect 32116 3780 32172 3782
rect 32196 3780 32252 3782
rect 31482 3576 31538 3632
rect 32126 3340 32128 3360
rect 32128 3340 32180 3360
rect 32180 3340 32182 3360
rect 32126 3304 32182 3340
rect 31758 3032 31814 3088
rect 32862 2796 32864 2816
rect 32864 2796 32916 2816
rect 32916 2796 32918 2816
rect 32862 2760 32918 2796
rect 31956 2746 32012 2748
rect 32036 2746 32092 2748
rect 32116 2746 32172 2748
rect 32196 2746 32252 2748
rect 31956 2694 32002 2746
rect 32002 2694 32012 2746
rect 32036 2694 32066 2746
rect 32066 2694 32078 2746
rect 32078 2694 32092 2746
rect 32116 2694 32130 2746
rect 32130 2694 32142 2746
rect 32142 2694 32172 2746
rect 32196 2694 32206 2746
rect 32206 2694 32252 2746
rect 31956 2692 32012 2694
rect 32036 2692 32092 2694
rect 32116 2692 32172 2694
rect 32196 2692 32252 2694
rect 31758 2488 31814 2544
rect 30746 1944 30802 2000
rect 31114 1672 31170 1728
rect 31850 2252 31852 2272
rect 31852 2252 31904 2272
rect 31904 2252 31906 2272
rect 31850 2216 31906 2252
rect 31482 1400 31538 1456
<< metal3 >>
rect 0 9890 120 9920
rect 17125 9890 17191 9893
rect 0 9888 17191 9890
rect 0 9832 17130 9888
rect 17186 9832 17191 9888
rect 0 9830 17191 9832
rect 0 9800 120 9830
rect 17125 9827 17191 9830
rect 30097 9890 30163 9893
rect 33630 9890 33750 9920
rect 30097 9888 33750 9890
rect 30097 9832 30102 9888
rect 30158 9832 33750 9888
rect 30097 9830 33750 9832
rect 30097 9827 30163 9830
rect 33630 9800 33750 9830
rect 0 9618 120 9648
rect 7741 9618 7807 9621
rect 0 9616 7807 9618
rect 0 9560 7746 9616
rect 7802 9560 7807 9616
rect 0 9558 7807 9560
rect 0 9528 120 9558
rect 7741 9555 7807 9558
rect 30833 9618 30899 9621
rect 33630 9618 33750 9648
rect 30833 9616 33750 9618
rect 30833 9560 30838 9616
rect 30894 9560 33750 9616
rect 30833 9558 33750 9560
rect 30833 9555 30899 9558
rect 33630 9528 33750 9558
rect 0 9346 120 9376
rect 4797 9346 4863 9349
rect 0 9344 4863 9346
rect 0 9288 4802 9344
rect 4858 9288 4863 9344
rect 0 9286 4863 9288
rect 0 9256 120 9286
rect 4797 9283 4863 9286
rect 31477 9346 31543 9349
rect 33630 9346 33750 9376
rect 31477 9344 33750 9346
rect 31477 9288 31482 9344
rect 31538 9288 33750 9344
rect 31477 9286 33750 9288
rect 31477 9283 31543 9286
rect 33630 9256 33750 9286
rect 0 9074 120 9104
rect 12433 9074 12499 9077
rect 0 9072 12499 9074
rect 0 9016 12438 9072
rect 12494 9016 12499 9072
rect 0 9014 12499 9016
rect 0 8984 120 9014
rect 12433 9011 12499 9014
rect 30465 9074 30531 9077
rect 33630 9074 33750 9104
rect 30465 9072 33750 9074
rect 30465 9016 30470 9072
rect 30526 9016 33750 9072
rect 30465 9014 33750 9016
rect 30465 9011 30531 9014
rect 33630 8984 33750 9014
rect 7373 8938 7439 8941
rect 2822 8936 7439 8938
rect 2822 8880 7378 8936
rect 7434 8880 7439 8936
rect 2822 8878 7439 8880
rect 0 8802 120 8832
rect 2822 8802 2882 8878
rect 7373 8875 7439 8878
rect 0 8742 2882 8802
rect 31017 8802 31083 8805
rect 33630 8802 33750 8832
rect 31017 8800 33750 8802
rect 31017 8744 31022 8800
rect 31078 8744 33750 8800
rect 31017 8742 33750 8744
rect 0 8712 120 8742
rect 31017 8739 31083 8742
rect 3006 8736 3322 8737
rect 3006 8672 3012 8736
rect 3076 8672 3092 8736
rect 3156 8672 3172 8736
rect 3236 8672 3252 8736
rect 3316 8672 3322 8736
rect 3006 8671 3322 8672
rect 9006 8736 9322 8737
rect 9006 8672 9012 8736
rect 9076 8672 9092 8736
rect 9156 8672 9172 8736
rect 9236 8672 9252 8736
rect 9316 8672 9322 8736
rect 9006 8671 9322 8672
rect 15006 8736 15322 8737
rect 15006 8672 15012 8736
rect 15076 8672 15092 8736
rect 15156 8672 15172 8736
rect 15236 8672 15252 8736
rect 15316 8672 15322 8736
rect 15006 8671 15322 8672
rect 21006 8736 21322 8737
rect 21006 8672 21012 8736
rect 21076 8672 21092 8736
rect 21156 8672 21172 8736
rect 21236 8672 21252 8736
rect 21316 8672 21322 8736
rect 21006 8671 21322 8672
rect 27006 8736 27322 8737
rect 27006 8672 27012 8736
rect 27076 8672 27092 8736
rect 27156 8672 27172 8736
rect 27236 8672 27252 8736
rect 27316 8672 27322 8736
rect 33630 8712 33750 8742
rect 27006 8671 27322 8672
rect 2865 8666 2931 8669
rect 1350 8664 2931 8666
rect 1350 8608 2870 8664
rect 2926 8608 2931 8664
rect 1350 8606 2931 8608
rect 0 8530 120 8560
rect 1350 8530 1410 8606
rect 2865 8603 2931 8606
rect 0 8470 1410 8530
rect 1577 8530 1643 8533
rect 25129 8530 25195 8533
rect 1577 8528 25195 8530
rect 1577 8472 1582 8528
rect 1638 8472 25134 8528
rect 25190 8472 25195 8528
rect 1577 8470 25195 8472
rect 0 8440 120 8470
rect 1577 8467 1643 8470
rect 25129 8467 25195 8470
rect 31385 8530 31451 8533
rect 33630 8530 33750 8560
rect 31385 8528 33750 8530
rect 31385 8472 31390 8528
rect 31446 8472 33750 8528
rect 31385 8470 33750 8472
rect 31385 8467 31451 8470
rect 33630 8440 33750 8470
rect 2865 8394 2931 8397
rect 15101 8394 15167 8397
rect 1718 8334 2514 8394
rect 0 8258 120 8288
rect 1718 8258 1778 8334
rect 0 8198 1778 8258
rect 2454 8258 2514 8334
rect 2865 8392 15167 8394
rect 2865 8336 2870 8392
rect 2926 8336 15106 8392
rect 15162 8336 15167 8392
rect 2865 8334 15167 8336
rect 2865 8331 2931 8334
rect 15101 8331 15167 8334
rect 7649 8258 7715 8261
rect 2454 8256 7715 8258
rect 2454 8200 7654 8256
rect 7710 8200 7715 8256
rect 2454 8198 7715 8200
rect 0 8168 120 8198
rect 7649 8195 7715 8198
rect 32397 8258 32463 8261
rect 33630 8258 33750 8288
rect 32397 8256 33750 8258
rect 32397 8200 32402 8256
rect 32458 8200 33750 8256
rect 32397 8198 33750 8200
rect 32397 8195 32463 8198
rect 1946 8192 2262 8193
rect 1946 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2262 8192
rect 1946 8127 2262 8128
rect 7946 8192 8262 8193
rect 7946 8128 7952 8192
rect 8016 8128 8032 8192
rect 8096 8128 8112 8192
rect 8176 8128 8192 8192
rect 8256 8128 8262 8192
rect 7946 8127 8262 8128
rect 13946 8192 14262 8193
rect 13946 8128 13952 8192
rect 14016 8128 14032 8192
rect 14096 8128 14112 8192
rect 14176 8128 14192 8192
rect 14256 8128 14262 8192
rect 13946 8127 14262 8128
rect 19946 8192 20262 8193
rect 19946 8128 19952 8192
rect 20016 8128 20032 8192
rect 20096 8128 20112 8192
rect 20176 8128 20192 8192
rect 20256 8128 20262 8192
rect 19946 8127 20262 8128
rect 25946 8192 26262 8193
rect 25946 8128 25952 8192
rect 26016 8128 26032 8192
rect 26096 8128 26112 8192
rect 26176 8128 26192 8192
rect 26256 8128 26262 8192
rect 25946 8127 26262 8128
rect 31946 8192 32262 8193
rect 31946 8128 31952 8192
rect 32016 8128 32032 8192
rect 32096 8128 32112 8192
rect 32176 8128 32192 8192
rect 32256 8128 32262 8192
rect 33630 8168 33750 8198
rect 31946 8127 32262 8128
rect 0 7986 120 8016
rect 14549 7986 14615 7989
rect 0 7984 14615 7986
rect 0 7928 14554 7984
rect 14610 7928 14615 7984
rect 0 7926 14615 7928
rect 0 7896 120 7926
rect 14549 7923 14615 7926
rect 31845 7986 31911 7989
rect 33630 7986 33750 8016
rect 31845 7984 33750 7986
rect 31845 7928 31850 7984
rect 31906 7928 33750 7984
rect 31845 7926 33750 7928
rect 31845 7923 31911 7926
rect 33630 7896 33750 7926
rect 6821 7850 6887 7853
rect 2822 7848 6887 7850
rect 2822 7792 6826 7848
rect 6882 7792 6887 7848
rect 2822 7790 6887 7792
rect 0 7714 120 7744
rect 2822 7714 2882 7790
rect 6821 7787 6887 7790
rect 0 7654 2882 7714
rect 32121 7714 32187 7717
rect 33630 7714 33750 7744
rect 32121 7712 33750 7714
rect 32121 7656 32126 7712
rect 32182 7656 33750 7712
rect 32121 7654 33750 7656
rect 0 7624 120 7654
rect 32121 7651 32187 7654
rect 3006 7648 3322 7649
rect 3006 7584 3012 7648
rect 3076 7584 3092 7648
rect 3156 7584 3172 7648
rect 3236 7584 3252 7648
rect 3316 7584 3322 7648
rect 3006 7583 3322 7584
rect 9006 7648 9322 7649
rect 9006 7584 9012 7648
rect 9076 7584 9092 7648
rect 9156 7584 9172 7648
rect 9236 7584 9252 7648
rect 9316 7584 9322 7648
rect 9006 7583 9322 7584
rect 15006 7648 15322 7649
rect 15006 7584 15012 7648
rect 15076 7584 15092 7648
rect 15156 7584 15172 7648
rect 15236 7584 15252 7648
rect 15316 7584 15322 7648
rect 15006 7583 15322 7584
rect 21006 7648 21322 7649
rect 21006 7584 21012 7648
rect 21076 7584 21092 7648
rect 21156 7584 21172 7648
rect 21236 7584 21252 7648
rect 21316 7584 21322 7648
rect 21006 7583 21322 7584
rect 27006 7648 27322 7649
rect 27006 7584 27012 7648
rect 27076 7584 27092 7648
rect 27156 7584 27172 7648
rect 27236 7584 27252 7648
rect 27316 7584 27322 7648
rect 33630 7624 33750 7654
rect 27006 7583 27322 7584
rect 0 7442 120 7472
rect 13905 7442 13971 7445
rect 0 7440 13971 7442
rect 0 7384 13910 7440
rect 13966 7384 13971 7440
rect 0 7382 13971 7384
rect 0 7352 120 7382
rect 13905 7379 13971 7382
rect 31753 7442 31819 7445
rect 33630 7442 33750 7472
rect 31753 7440 33750 7442
rect 31753 7384 31758 7440
rect 31814 7384 33750 7440
rect 31753 7382 33750 7384
rect 31753 7379 31819 7382
rect 33630 7352 33750 7382
rect 5533 7306 5599 7309
rect 1718 7304 5599 7306
rect 1718 7248 5538 7304
rect 5594 7248 5599 7304
rect 1718 7246 5599 7248
rect 0 7170 120 7200
rect 1718 7170 1778 7246
rect 5533 7243 5599 7246
rect 5901 7306 5967 7309
rect 31293 7306 31359 7309
rect 5901 7304 31359 7306
rect 5901 7248 5906 7304
rect 5962 7248 31298 7304
rect 31354 7248 31359 7304
rect 5901 7246 31359 7248
rect 5901 7243 5967 7246
rect 31293 7243 31359 7246
rect 0 7110 1778 7170
rect 32765 7170 32831 7173
rect 33630 7170 33750 7200
rect 32765 7168 33750 7170
rect 32765 7112 32770 7168
rect 32826 7112 33750 7168
rect 32765 7110 33750 7112
rect 0 7080 120 7110
rect 32765 7107 32831 7110
rect 1946 7104 2262 7105
rect 1946 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2262 7104
rect 1946 7039 2262 7040
rect 7946 7104 8262 7105
rect 7946 7040 7952 7104
rect 8016 7040 8032 7104
rect 8096 7040 8112 7104
rect 8176 7040 8192 7104
rect 8256 7040 8262 7104
rect 7946 7039 8262 7040
rect 13946 7104 14262 7105
rect 13946 7040 13952 7104
rect 14016 7040 14032 7104
rect 14096 7040 14112 7104
rect 14176 7040 14192 7104
rect 14256 7040 14262 7104
rect 13946 7039 14262 7040
rect 19946 7104 20262 7105
rect 19946 7040 19952 7104
rect 20016 7040 20032 7104
rect 20096 7040 20112 7104
rect 20176 7040 20192 7104
rect 20256 7040 20262 7104
rect 19946 7039 20262 7040
rect 25946 7104 26262 7105
rect 25946 7040 25952 7104
rect 26016 7040 26032 7104
rect 26096 7040 26112 7104
rect 26176 7040 26192 7104
rect 26256 7040 26262 7104
rect 25946 7039 26262 7040
rect 31946 7104 32262 7105
rect 31946 7040 31952 7104
rect 32016 7040 32032 7104
rect 32096 7040 32112 7104
rect 32176 7040 32192 7104
rect 32256 7040 32262 7104
rect 33630 7080 33750 7110
rect 31946 7039 32262 7040
rect 0 6898 120 6928
rect 6269 6898 6335 6901
rect 0 6896 6335 6898
rect 0 6840 6274 6896
rect 6330 6840 6335 6896
rect 0 6838 6335 6840
rect 0 6808 120 6838
rect 6269 6835 6335 6838
rect 31753 6898 31819 6901
rect 33630 6898 33750 6928
rect 31753 6896 33750 6898
rect 31753 6840 31758 6896
rect 31814 6840 33750 6896
rect 31753 6838 33750 6840
rect 31753 6835 31819 6838
rect 33630 6808 33750 6838
rect 10961 6762 11027 6765
rect 2822 6760 11027 6762
rect 2822 6704 10966 6760
rect 11022 6704 11027 6760
rect 2822 6702 11027 6704
rect 0 6626 120 6656
rect 2822 6626 2882 6702
rect 10961 6699 11027 6702
rect 0 6566 2882 6626
rect 31385 6626 31451 6629
rect 33630 6626 33750 6656
rect 31385 6624 33750 6626
rect 31385 6568 31390 6624
rect 31446 6568 33750 6624
rect 31385 6566 33750 6568
rect 0 6536 120 6566
rect 31385 6563 31451 6566
rect 3006 6560 3322 6561
rect 3006 6496 3012 6560
rect 3076 6496 3092 6560
rect 3156 6496 3172 6560
rect 3236 6496 3252 6560
rect 3316 6496 3322 6560
rect 3006 6495 3322 6496
rect 9006 6560 9322 6561
rect 9006 6496 9012 6560
rect 9076 6496 9092 6560
rect 9156 6496 9172 6560
rect 9236 6496 9252 6560
rect 9316 6496 9322 6560
rect 9006 6495 9322 6496
rect 15006 6560 15322 6561
rect 15006 6496 15012 6560
rect 15076 6496 15092 6560
rect 15156 6496 15172 6560
rect 15236 6496 15252 6560
rect 15316 6496 15322 6560
rect 15006 6495 15322 6496
rect 21006 6560 21322 6561
rect 21006 6496 21012 6560
rect 21076 6496 21092 6560
rect 21156 6496 21172 6560
rect 21236 6496 21252 6560
rect 21316 6496 21322 6560
rect 21006 6495 21322 6496
rect 27006 6560 27322 6561
rect 27006 6496 27012 6560
rect 27076 6496 27092 6560
rect 27156 6496 27172 6560
rect 27236 6496 27252 6560
rect 27316 6496 27322 6560
rect 33630 6536 33750 6566
rect 27006 6495 27322 6496
rect 0 6354 120 6384
rect 5533 6354 5599 6357
rect 0 6352 5599 6354
rect 0 6296 5538 6352
rect 5594 6296 5599 6352
rect 0 6294 5599 6296
rect 0 6264 120 6294
rect 5533 6291 5599 6294
rect 31845 6354 31911 6357
rect 33630 6354 33750 6384
rect 31845 6352 33750 6354
rect 31845 6296 31850 6352
rect 31906 6296 33750 6352
rect 31845 6294 33750 6296
rect 31845 6291 31911 6294
rect 33630 6264 33750 6294
rect 16481 6218 16547 6221
rect 1718 6216 16547 6218
rect 1718 6160 16486 6216
rect 16542 6160 16547 6216
rect 1718 6158 16547 6160
rect 0 6082 120 6112
rect 1718 6082 1778 6158
rect 16481 6155 16547 6158
rect 31477 6218 31543 6221
rect 31477 6216 32690 6218
rect 31477 6160 31482 6216
rect 31538 6160 32690 6216
rect 31477 6158 32690 6160
rect 31477 6155 31543 6158
rect 0 6022 1778 6082
rect 32630 6082 32690 6158
rect 33630 6082 33750 6112
rect 32630 6022 33750 6082
rect 0 5992 120 6022
rect 1946 6016 2262 6017
rect 1946 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2262 6016
rect 1946 5951 2262 5952
rect 7946 6016 8262 6017
rect 7946 5952 7952 6016
rect 8016 5952 8032 6016
rect 8096 5952 8112 6016
rect 8176 5952 8192 6016
rect 8256 5952 8262 6016
rect 7946 5951 8262 5952
rect 13946 6016 14262 6017
rect 13946 5952 13952 6016
rect 14016 5952 14032 6016
rect 14096 5952 14112 6016
rect 14176 5952 14192 6016
rect 14256 5952 14262 6016
rect 13946 5951 14262 5952
rect 19946 6016 20262 6017
rect 19946 5952 19952 6016
rect 20016 5952 20032 6016
rect 20096 5952 20112 6016
rect 20176 5952 20192 6016
rect 20256 5952 20262 6016
rect 19946 5951 20262 5952
rect 25946 6016 26262 6017
rect 25946 5952 25952 6016
rect 26016 5952 26032 6016
rect 26096 5952 26112 6016
rect 26176 5952 26192 6016
rect 26256 5952 26262 6016
rect 25946 5951 26262 5952
rect 31946 6016 32262 6017
rect 31946 5952 31952 6016
rect 32016 5952 32032 6016
rect 32096 5952 32112 6016
rect 32176 5952 32192 6016
rect 32256 5952 32262 6016
rect 33630 5992 33750 6022
rect 31946 5951 32262 5952
rect 0 5810 120 5840
rect 13721 5810 13787 5813
rect 0 5808 13787 5810
rect 0 5752 13726 5808
rect 13782 5752 13787 5808
rect 0 5750 13787 5752
rect 0 5720 120 5750
rect 13721 5747 13787 5750
rect 32121 5810 32187 5813
rect 33630 5810 33750 5840
rect 32121 5808 33750 5810
rect 32121 5752 32126 5808
rect 32182 5752 33750 5808
rect 32121 5750 33750 5752
rect 32121 5747 32187 5750
rect 33630 5720 33750 5750
rect 2822 5614 3618 5674
rect 0 5538 120 5568
rect 2822 5538 2882 5614
rect 0 5478 2882 5538
rect 3558 5538 3618 5614
rect 8710 5614 9506 5674
rect 8710 5538 8770 5614
rect 3558 5478 8770 5538
rect 9446 5538 9506 5614
rect 12709 5538 12775 5541
rect 9446 5536 12775 5538
rect 9446 5480 12714 5536
rect 12770 5480 12775 5536
rect 9446 5478 12775 5480
rect 0 5448 120 5478
rect 12709 5475 12775 5478
rect 31753 5538 31819 5541
rect 33630 5538 33750 5568
rect 31753 5536 33750 5538
rect 31753 5480 31758 5536
rect 31814 5480 33750 5536
rect 31753 5478 33750 5480
rect 31753 5475 31819 5478
rect 3006 5472 3322 5473
rect 3006 5408 3012 5472
rect 3076 5408 3092 5472
rect 3156 5408 3172 5472
rect 3236 5408 3252 5472
rect 3316 5408 3322 5472
rect 3006 5407 3322 5408
rect 9006 5472 9322 5473
rect 9006 5408 9012 5472
rect 9076 5408 9092 5472
rect 9156 5408 9172 5472
rect 9236 5408 9252 5472
rect 9316 5408 9322 5472
rect 9006 5407 9322 5408
rect 15006 5472 15322 5473
rect 15006 5408 15012 5472
rect 15076 5408 15092 5472
rect 15156 5408 15172 5472
rect 15236 5408 15252 5472
rect 15316 5408 15322 5472
rect 15006 5407 15322 5408
rect 21006 5472 21322 5473
rect 21006 5408 21012 5472
rect 21076 5408 21092 5472
rect 21156 5408 21172 5472
rect 21236 5408 21252 5472
rect 21316 5408 21322 5472
rect 21006 5407 21322 5408
rect 27006 5472 27322 5473
rect 27006 5408 27012 5472
rect 27076 5408 27092 5472
rect 27156 5408 27172 5472
rect 27236 5408 27252 5472
rect 27316 5408 27322 5472
rect 33630 5448 33750 5478
rect 27006 5407 27322 5408
rect 0 5266 120 5296
rect 11881 5266 11947 5269
rect 0 5264 11947 5266
rect 0 5208 11886 5264
rect 11942 5208 11947 5264
rect 0 5206 11947 5208
rect 0 5176 120 5206
rect 11881 5203 11947 5206
rect 32029 5266 32095 5269
rect 33630 5266 33750 5296
rect 32029 5264 33750 5266
rect 32029 5208 32034 5264
rect 32090 5208 33750 5264
rect 32029 5206 33750 5208
rect 32029 5203 32095 5206
rect 33630 5176 33750 5206
rect 16941 5130 17007 5133
rect 1718 5128 17007 5130
rect 1718 5072 16946 5128
rect 17002 5072 17007 5128
rect 1718 5070 17007 5072
rect 0 4994 120 5024
rect 1718 4994 1778 5070
rect 16941 5067 17007 5070
rect 0 4934 1778 4994
rect 32857 4994 32923 4997
rect 33630 4994 33750 5024
rect 32857 4992 33750 4994
rect 32857 4936 32862 4992
rect 32918 4936 33750 4992
rect 32857 4934 33750 4936
rect 0 4904 120 4934
rect 32857 4931 32923 4934
rect 1946 4928 2262 4929
rect 1946 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2262 4928
rect 1946 4863 2262 4864
rect 7946 4928 8262 4929
rect 7946 4864 7952 4928
rect 8016 4864 8032 4928
rect 8096 4864 8112 4928
rect 8176 4864 8192 4928
rect 8256 4864 8262 4928
rect 7946 4863 8262 4864
rect 13946 4928 14262 4929
rect 13946 4864 13952 4928
rect 14016 4864 14032 4928
rect 14096 4864 14112 4928
rect 14176 4864 14192 4928
rect 14256 4864 14262 4928
rect 13946 4863 14262 4864
rect 19946 4928 20262 4929
rect 19946 4864 19952 4928
rect 20016 4864 20032 4928
rect 20096 4864 20112 4928
rect 20176 4864 20192 4928
rect 20256 4864 20262 4928
rect 19946 4863 20262 4864
rect 25946 4928 26262 4929
rect 25946 4864 25952 4928
rect 26016 4864 26032 4928
rect 26096 4864 26112 4928
rect 26176 4864 26192 4928
rect 26256 4864 26262 4928
rect 25946 4863 26262 4864
rect 31946 4928 32262 4929
rect 31946 4864 31952 4928
rect 32016 4864 32032 4928
rect 32096 4864 32112 4928
rect 32176 4864 32192 4928
rect 32256 4864 32262 4928
rect 33630 4904 33750 4934
rect 31946 4863 32262 4864
rect 0 4722 120 4752
rect 19333 4722 19399 4725
rect 0 4720 19399 4722
rect 0 4664 19338 4720
rect 19394 4664 19399 4720
rect 0 4662 19399 4664
rect 0 4632 120 4662
rect 19333 4659 19399 4662
rect 31477 4722 31543 4725
rect 33630 4722 33750 4752
rect 31477 4720 33750 4722
rect 31477 4664 31482 4720
rect 31538 4664 33750 4720
rect 31477 4662 33750 4664
rect 31477 4659 31543 4662
rect 33630 4632 33750 4662
rect 20897 4586 20963 4589
rect 2822 4584 20963 4586
rect 2822 4528 20902 4584
rect 20958 4528 20963 4584
rect 2822 4526 20963 4528
rect 0 4450 120 4480
rect 2822 4450 2882 4526
rect 20897 4523 20963 4526
rect 0 4390 2882 4450
rect 32121 4450 32187 4453
rect 33630 4450 33750 4480
rect 32121 4448 33750 4450
rect 32121 4392 32126 4448
rect 32182 4392 33750 4448
rect 32121 4390 33750 4392
rect 0 4360 120 4390
rect 32121 4387 32187 4390
rect 3006 4384 3322 4385
rect 3006 4320 3012 4384
rect 3076 4320 3092 4384
rect 3156 4320 3172 4384
rect 3236 4320 3252 4384
rect 3316 4320 3322 4384
rect 3006 4319 3322 4320
rect 9006 4384 9322 4385
rect 9006 4320 9012 4384
rect 9076 4320 9092 4384
rect 9156 4320 9172 4384
rect 9236 4320 9252 4384
rect 9316 4320 9322 4384
rect 9006 4319 9322 4320
rect 15006 4384 15322 4385
rect 15006 4320 15012 4384
rect 15076 4320 15092 4384
rect 15156 4320 15172 4384
rect 15236 4320 15252 4384
rect 15316 4320 15322 4384
rect 15006 4319 15322 4320
rect 21006 4384 21322 4385
rect 21006 4320 21012 4384
rect 21076 4320 21092 4384
rect 21156 4320 21172 4384
rect 21236 4320 21252 4384
rect 21316 4320 21322 4384
rect 21006 4319 21322 4320
rect 27006 4384 27322 4385
rect 27006 4320 27012 4384
rect 27076 4320 27092 4384
rect 27156 4320 27172 4384
rect 27236 4320 27252 4384
rect 27316 4320 27322 4384
rect 33630 4360 33750 4390
rect 27006 4319 27322 4320
rect 0 4178 120 4208
rect 23013 4178 23079 4181
rect 0 4176 23079 4178
rect 0 4120 23018 4176
rect 23074 4120 23079 4176
rect 0 4118 23079 4120
rect 0 4088 120 4118
rect 23013 4115 23079 4118
rect 31753 4178 31819 4181
rect 33630 4178 33750 4208
rect 31753 4176 33750 4178
rect 31753 4120 31758 4176
rect 31814 4120 33750 4176
rect 31753 4118 33750 4120
rect 31753 4115 31819 4118
rect 33630 4088 33750 4118
rect 12525 4042 12591 4045
rect 1718 4040 12591 4042
rect 1718 3984 12530 4040
rect 12586 3984 12591 4040
rect 1718 3982 12591 3984
rect 0 3906 120 3936
rect 1718 3906 1778 3982
rect 12525 3979 12591 3982
rect 19793 4042 19859 4045
rect 28993 4042 29059 4045
rect 19793 4040 29059 4042
rect 19793 3984 19798 4040
rect 19854 3984 28998 4040
rect 29054 3984 29059 4040
rect 19793 3982 29059 3984
rect 19793 3979 19859 3982
rect 28993 3979 29059 3982
rect 0 3846 1778 3906
rect 32857 3906 32923 3909
rect 33630 3906 33750 3936
rect 32857 3904 33750 3906
rect 32857 3848 32862 3904
rect 32918 3848 33750 3904
rect 32857 3846 33750 3848
rect 0 3816 120 3846
rect 32857 3843 32923 3846
rect 1946 3840 2262 3841
rect 1946 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2262 3840
rect 1946 3775 2262 3776
rect 7946 3840 8262 3841
rect 7946 3776 7952 3840
rect 8016 3776 8032 3840
rect 8096 3776 8112 3840
rect 8176 3776 8192 3840
rect 8256 3776 8262 3840
rect 7946 3775 8262 3776
rect 13946 3840 14262 3841
rect 13946 3776 13952 3840
rect 14016 3776 14032 3840
rect 14096 3776 14112 3840
rect 14176 3776 14192 3840
rect 14256 3776 14262 3840
rect 13946 3775 14262 3776
rect 19946 3840 20262 3841
rect 19946 3776 19952 3840
rect 20016 3776 20032 3840
rect 20096 3776 20112 3840
rect 20176 3776 20192 3840
rect 20256 3776 20262 3840
rect 19946 3775 20262 3776
rect 25946 3840 26262 3841
rect 25946 3776 25952 3840
rect 26016 3776 26032 3840
rect 26096 3776 26112 3840
rect 26176 3776 26192 3840
rect 26256 3776 26262 3840
rect 25946 3775 26262 3776
rect 31946 3840 32262 3841
rect 31946 3776 31952 3840
rect 32016 3776 32032 3840
rect 32096 3776 32112 3840
rect 32176 3776 32192 3840
rect 32256 3776 32262 3840
rect 33630 3816 33750 3846
rect 31946 3775 32262 3776
rect 0 3634 120 3664
rect 13077 3634 13143 3637
rect 0 3632 13143 3634
rect 0 3576 13082 3632
rect 13138 3576 13143 3632
rect 0 3574 13143 3576
rect 0 3544 120 3574
rect 13077 3571 13143 3574
rect 31477 3634 31543 3637
rect 33630 3634 33750 3664
rect 31477 3632 33750 3634
rect 31477 3576 31482 3632
rect 31538 3576 33750 3632
rect 31477 3574 33750 3576
rect 31477 3571 31543 3574
rect 33630 3544 33750 3574
rect 25221 3498 25287 3501
rect 2822 3496 25287 3498
rect 2822 3440 25226 3496
rect 25282 3440 25287 3496
rect 2822 3438 25287 3440
rect 0 3362 120 3392
rect 2822 3362 2882 3438
rect 25221 3435 25287 3438
rect 0 3302 2882 3362
rect 32121 3362 32187 3365
rect 33630 3362 33750 3392
rect 32121 3360 33750 3362
rect 32121 3304 32126 3360
rect 32182 3304 33750 3360
rect 32121 3302 33750 3304
rect 0 3272 120 3302
rect 32121 3299 32187 3302
rect 3006 3296 3322 3297
rect 3006 3232 3012 3296
rect 3076 3232 3092 3296
rect 3156 3232 3172 3296
rect 3236 3232 3252 3296
rect 3316 3232 3322 3296
rect 3006 3231 3322 3232
rect 9006 3296 9322 3297
rect 9006 3232 9012 3296
rect 9076 3232 9092 3296
rect 9156 3232 9172 3296
rect 9236 3232 9252 3296
rect 9316 3232 9322 3296
rect 9006 3231 9322 3232
rect 15006 3296 15322 3297
rect 15006 3232 15012 3296
rect 15076 3232 15092 3296
rect 15156 3232 15172 3296
rect 15236 3232 15252 3296
rect 15316 3232 15322 3296
rect 15006 3231 15322 3232
rect 21006 3296 21322 3297
rect 21006 3232 21012 3296
rect 21076 3232 21092 3296
rect 21156 3232 21172 3296
rect 21236 3232 21252 3296
rect 21316 3232 21322 3296
rect 21006 3231 21322 3232
rect 27006 3296 27322 3297
rect 27006 3232 27012 3296
rect 27076 3232 27092 3296
rect 27156 3232 27172 3296
rect 27236 3232 27252 3296
rect 27316 3232 27322 3296
rect 33630 3272 33750 3302
rect 27006 3231 27322 3232
rect 0 3090 120 3120
rect 25773 3090 25839 3093
rect 0 3088 25839 3090
rect 0 3032 25778 3088
rect 25834 3032 25839 3088
rect 0 3030 25839 3032
rect 0 3000 120 3030
rect 25773 3027 25839 3030
rect 31753 3090 31819 3093
rect 33630 3090 33750 3120
rect 31753 3088 33750 3090
rect 31753 3032 31758 3088
rect 31814 3032 33750 3088
rect 31753 3030 33750 3032
rect 31753 3027 31819 3030
rect 33630 3000 33750 3030
rect 26233 2954 26299 2957
rect 1718 2952 26299 2954
rect 1718 2896 26238 2952
rect 26294 2896 26299 2952
rect 1718 2894 26299 2896
rect 0 2818 120 2848
rect 1718 2818 1778 2894
rect 26233 2891 26299 2894
rect 0 2758 1778 2818
rect 32857 2818 32923 2821
rect 33630 2818 33750 2848
rect 32857 2816 33750 2818
rect 32857 2760 32862 2816
rect 32918 2760 33750 2816
rect 32857 2758 33750 2760
rect 0 2728 120 2758
rect 32857 2755 32923 2758
rect 1946 2752 2262 2753
rect 1946 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2262 2752
rect 1946 2687 2262 2688
rect 7946 2752 8262 2753
rect 7946 2688 7952 2752
rect 8016 2688 8032 2752
rect 8096 2688 8112 2752
rect 8176 2688 8192 2752
rect 8256 2688 8262 2752
rect 7946 2687 8262 2688
rect 13946 2752 14262 2753
rect 13946 2688 13952 2752
rect 14016 2688 14032 2752
rect 14096 2688 14112 2752
rect 14176 2688 14192 2752
rect 14256 2688 14262 2752
rect 13946 2687 14262 2688
rect 19946 2752 20262 2753
rect 19946 2688 19952 2752
rect 20016 2688 20032 2752
rect 20096 2688 20112 2752
rect 20176 2688 20192 2752
rect 20256 2688 20262 2752
rect 19946 2687 20262 2688
rect 25946 2752 26262 2753
rect 25946 2688 25952 2752
rect 26016 2688 26032 2752
rect 26096 2688 26112 2752
rect 26176 2688 26192 2752
rect 26256 2688 26262 2752
rect 25946 2687 26262 2688
rect 31946 2752 32262 2753
rect 31946 2688 31952 2752
rect 32016 2688 32032 2752
rect 32096 2688 32112 2752
rect 32176 2688 32192 2752
rect 32256 2688 32262 2752
rect 33630 2728 33750 2758
rect 31946 2687 32262 2688
rect 21633 2682 21699 2685
rect 24853 2682 24919 2685
rect 21633 2680 24919 2682
rect 21633 2624 21638 2680
rect 21694 2624 24858 2680
rect 24914 2624 24919 2680
rect 21633 2622 24919 2624
rect 21633 2619 21699 2622
rect 24853 2619 24919 2622
rect 0 2546 120 2576
rect 18965 2546 19031 2549
rect 0 2544 19031 2546
rect 0 2488 18970 2544
rect 19026 2488 19031 2544
rect 0 2486 19031 2488
rect 0 2456 120 2486
rect 18965 2483 19031 2486
rect 31753 2546 31819 2549
rect 33630 2546 33750 2576
rect 31753 2544 33750 2546
rect 31753 2488 31758 2544
rect 31814 2488 33750 2544
rect 31753 2486 33750 2488
rect 31753 2483 31819 2486
rect 33630 2456 33750 2486
rect 10777 2410 10843 2413
rect 17125 2410 17191 2413
rect 10777 2408 17191 2410
rect 10777 2352 10782 2408
rect 10838 2352 17130 2408
rect 17186 2352 17191 2408
rect 10777 2350 17191 2352
rect 10777 2347 10843 2350
rect 17125 2347 17191 2350
rect 19701 2410 19767 2413
rect 20529 2410 20595 2413
rect 19701 2408 20595 2410
rect 19701 2352 19706 2408
rect 19762 2352 20534 2408
rect 20590 2352 20595 2408
rect 19701 2350 20595 2352
rect 19701 2347 19767 2350
rect 20529 2347 20595 2350
rect 0 2274 120 2304
rect 2865 2274 2931 2277
rect 0 2272 2931 2274
rect 0 2216 2870 2272
rect 2926 2216 2931 2272
rect 0 2214 2931 2216
rect 0 2184 120 2214
rect 2865 2211 2931 2214
rect 31845 2274 31911 2277
rect 33630 2274 33750 2304
rect 31845 2272 33750 2274
rect 31845 2216 31850 2272
rect 31906 2216 33750 2272
rect 31845 2214 33750 2216
rect 31845 2211 31911 2214
rect 3006 2208 3322 2209
rect 3006 2144 3012 2208
rect 3076 2144 3092 2208
rect 3156 2144 3172 2208
rect 3236 2144 3252 2208
rect 3316 2144 3322 2208
rect 3006 2143 3322 2144
rect 9006 2208 9322 2209
rect 9006 2144 9012 2208
rect 9076 2144 9092 2208
rect 9156 2144 9172 2208
rect 9236 2144 9252 2208
rect 9316 2144 9322 2208
rect 9006 2143 9322 2144
rect 15006 2208 15322 2209
rect 15006 2144 15012 2208
rect 15076 2144 15092 2208
rect 15156 2144 15172 2208
rect 15236 2144 15252 2208
rect 15316 2144 15322 2208
rect 15006 2143 15322 2144
rect 21006 2208 21322 2209
rect 21006 2144 21012 2208
rect 21076 2144 21092 2208
rect 21156 2144 21172 2208
rect 21236 2144 21252 2208
rect 21316 2144 21322 2208
rect 21006 2143 21322 2144
rect 27006 2208 27322 2209
rect 27006 2144 27012 2208
rect 27076 2144 27092 2208
rect 27156 2144 27172 2208
rect 27236 2144 27252 2208
rect 27316 2144 27322 2208
rect 33630 2184 33750 2214
rect 27006 2143 27322 2144
rect 0 2002 120 2032
rect 21725 2002 21791 2005
rect 0 2000 21791 2002
rect 0 1944 21730 2000
rect 21786 1944 21791 2000
rect 0 1942 21791 1944
rect 0 1912 120 1942
rect 21725 1939 21791 1942
rect 30741 2002 30807 2005
rect 33630 2002 33750 2032
rect 30741 2000 33750 2002
rect 30741 1944 30746 2000
rect 30802 1944 33750 2000
rect 30741 1942 33750 1944
rect 30741 1939 30807 1942
rect 33630 1912 33750 1942
rect 2865 1866 2931 1869
rect 20713 1866 20779 1869
rect 2865 1864 20779 1866
rect 2865 1808 2870 1864
rect 2926 1808 20718 1864
rect 20774 1808 20779 1864
rect 2865 1806 20779 1808
rect 2865 1803 2931 1806
rect 20713 1803 20779 1806
rect 0 1730 120 1760
rect 20069 1730 20135 1733
rect 0 1728 20135 1730
rect 0 1672 20074 1728
rect 20130 1672 20135 1728
rect 0 1670 20135 1672
rect 0 1640 120 1670
rect 20069 1667 20135 1670
rect 31109 1730 31175 1733
rect 33630 1730 33750 1760
rect 31109 1728 33750 1730
rect 31109 1672 31114 1728
rect 31170 1672 33750 1728
rect 31109 1670 33750 1672
rect 31109 1667 31175 1670
rect 33630 1640 33750 1670
rect 0 1458 120 1488
rect 17309 1458 17375 1461
rect 0 1456 17375 1458
rect 0 1400 17314 1456
rect 17370 1400 17375 1456
rect 0 1398 17375 1400
rect 0 1368 120 1398
rect 17309 1395 17375 1398
rect 31477 1458 31543 1461
rect 33630 1458 33750 1488
rect 31477 1456 33750 1458
rect 31477 1400 31482 1456
rect 31538 1400 33750 1456
rect 31477 1398 33750 1400
rect 31477 1395 31543 1398
rect 33630 1368 33750 1398
rect 10501 1322 10567 1325
rect 18045 1322 18111 1325
rect 10501 1320 18111 1322
rect 10501 1264 10506 1320
rect 10562 1264 18050 1320
rect 18106 1264 18111 1320
rect 10501 1262 18111 1264
rect 10501 1259 10567 1262
rect 18045 1259 18111 1262
rect 10225 1186 10291 1189
rect 18689 1186 18755 1189
rect 10225 1184 18755 1186
rect 10225 1128 10230 1184
rect 10286 1128 18694 1184
rect 18750 1128 18755 1184
rect 10225 1126 18755 1128
rect 10225 1123 10291 1126
rect 18689 1123 18755 1126
<< via3 >>
rect 3012 8732 3076 8736
rect 3012 8676 3016 8732
rect 3016 8676 3072 8732
rect 3072 8676 3076 8732
rect 3012 8672 3076 8676
rect 3092 8732 3156 8736
rect 3092 8676 3096 8732
rect 3096 8676 3152 8732
rect 3152 8676 3156 8732
rect 3092 8672 3156 8676
rect 3172 8732 3236 8736
rect 3172 8676 3176 8732
rect 3176 8676 3232 8732
rect 3232 8676 3236 8732
rect 3172 8672 3236 8676
rect 3252 8732 3316 8736
rect 3252 8676 3256 8732
rect 3256 8676 3312 8732
rect 3312 8676 3316 8732
rect 3252 8672 3316 8676
rect 9012 8732 9076 8736
rect 9012 8676 9016 8732
rect 9016 8676 9072 8732
rect 9072 8676 9076 8732
rect 9012 8672 9076 8676
rect 9092 8732 9156 8736
rect 9092 8676 9096 8732
rect 9096 8676 9152 8732
rect 9152 8676 9156 8732
rect 9092 8672 9156 8676
rect 9172 8732 9236 8736
rect 9172 8676 9176 8732
rect 9176 8676 9232 8732
rect 9232 8676 9236 8732
rect 9172 8672 9236 8676
rect 9252 8732 9316 8736
rect 9252 8676 9256 8732
rect 9256 8676 9312 8732
rect 9312 8676 9316 8732
rect 9252 8672 9316 8676
rect 15012 8732 15076 8736
rect 15012 8676 15016 8732
rect 15016 8676 15072 8732
rect 15072 8676 15076 8732
rect 15012 8672 15076 8676
rect 15092 8732 15156 8736
rect 15092 8676 15096 8732
rect 15096 8676 15152 8732
rect 15152 8676 15156 8732
rect 15092 8672 15156 8676
rect 15172 8732 15236 8736
rect 15172 8676 15176 8732
rect 15176 8676 15232 8732
rect 15232 8676 15236 8732
rect 15172 8672 15236 8676
rect 15252 8732 15316 8736
rect 15252 8676 15256 8732
rect 15256 8676 15312 8732
rect 15312 8676 15316 8732
rect 15252 8672 15316 8676
rect 21012 8732 21076 8736
rect 21012 8676 21016 8732
rect 21016 8676 21072 8732
rect 21072 8676 21076 8732
rect 21012 8672 21076 8676
rect 21092 8732 21156 8736
rect 21092 8676 21096 8732
rect 21096 8676 21152 8732
rect 21152 8676 21156 8732
rect 21092 8672 21156 8676
rect 21172 8732 21236 8736
rect 21172 8676 21176 8732
rect 21176 8676 21232 8732
rect 21232 8676 21236 8732
rect 21172 8672 21236 8676
rect 21252 8732 21316 8736
rect 21252 8676 21256 8732
rect 21256 8676 21312 8732
rect 21312 8676 21316 8732
rect 21252 8672 21316 8676
rect 27012 8732 27076 8736
rect 27012 8676 27016 8732
rect 27016 8676 27072 8732
rect 27072 8676 27076 8732
rect 27012 8672 27076 8676
rect 27092 8732 27156 8736
rect 27092 8676 27096 8732
rect 27096 8676 27152 8732
rect 27152 8676 27156 8732
rect 27092 8672 27156 8676
rect 27172 8732 27236 8736
rect 27172 8676 27176 8732
rect 27176 8676 27232 8732
rect 27232 8676 27236 8732
rect 27172 8672 27236 8676
rect 27252 8732 27316 8736
rect 27252 8676 27256 8732
rect 27256 8676 27312 8732
rect 27312 8676 27316 8732
rect 27252 8672 27316 8676
rect 1952 8188 2016 8192
rect 1952 8132 1956 8188
rect 1956 8132 2012 8188
rect 2012 8132 2016 8188
rect 1952 8128 2016 8132
rect 2032 8188 2096 8192
rect 2032 8132 2036 8188
rect 2036 8132 2092 8188
rect 2092 8132 2096 8188
rect 2032 8128 2096 8132
rect 2112 8188 2176 8192
rect 2112 8132 2116 8188
rect 2116 8132 2172 8188
rect 2172 8132 2176 8188
rect 2112 8128 2176 8132
rect 2192 8188 2256 8192
rect 2192 8132 2196 8188
rect 2196 8132 2252 8188
rect 2252 8132 2256 8188
rect 2192 8128 2256 8132
rect 7952 8188 8016 8192
rect 7952 8132 7956 8188
rect 7956 8132 8012 8188
rect 8012 8132 8016 8188
rect 7952 8128 8016 8132
rect 8032 8188 8096 8192
rect 8032 8132 8036 8188
rect 8036 8132 8092 8188
rect 8092 8132 8096 8188
rect 8032 8128 8096 8132
rect 8112 8188 8176 8192
rect 8112 8132 8116 8188
rect 8116 8132 8172 8188
rect 8172 8132 8176 8188
rect 8112 8128 8176 8132
rect 8192 8188 8256 8192
rect 8192 8132 8196 8188
rect 8196 8132 8252 8188
rect 8252 8132 8256 8188
rect 8192 8128 8256 8132
rect 13952 8188 14016 8192
rect 13952 8132 13956 8188
rect 13956 8132 14012 8188
rect 14012 8132 14016 8188
rect 13952 8128 14016 8132
rect 14032 8188 14096 8192
rect 14032 8132 14036 8188
rect 14036 8132 14092 8188
rect 14092 8132 14096 8188
rect 14032 8128 14096 8132
rect 14112 8188 14176 8192
rect 14112 8132 14116 8188
rect 14116 8132 14172 8188
rect 14172 8132 14176 8188
rect 14112 8128 14176 8132
rect 14192 8188 14256 8192
rect 14192 8132 14196 8188
rect 14196 8132 14252 8188
rect 14252 8132 14256 8188
rect 14192 8128 14256 8132
rect 19952 8188 20016 8192
rect 19952 8132 19956 8188
rect 19956 8132 20012 8188
rect 20012 8132 20016 8188
rect 19952 8128 20016 8132
rect 20032 8188 20096 8192
rect 20032 8132 20036 8188
rect 20036 8132 20092 8188
rect 20092 8132 20096 8188
rect 20032 8128 20096 8132
rect 20112 8188 20176 8192
rect 20112 8132 20116 8188
rect 20116 8132 20172 8188
rect 20172 8132 20176 8188
rect 20112 8128 20176 8132
rect 20192 8188 20256 8192
rect 20192 8132 20196 8188
rect 20196 8132 20252 8188
rect 20252 8132 20256 8188
rect 20192 8128 20256 8132
rect 25952 8188 26016 8192
rect 25952 8132 25956 8188
rect 25956 8132 26012 8188
rect 26012 8132 26016 8188
rect 25952 8128 26016 8132
rect 26032 8188 26096 8192
rect 26032 8132 26036 8188
rect 26036 8132 26092 8188
rect 26092 8132 26096 8188
rect 26032 8128 26096 8132
rect 26112 8188 26176 8192
rect 26112 8132 26116 8188
rect 26116 8132 26172 8188
rect 26172 8132 26176 8188
rect 26112 8128 26176 8132
rect 26192 8188 26256 8192
rect 26192 8132 26196 8188
rect 26196 8132 26252 8188
rect 26252 8132 26256 8188
rect 26192 8128 26256 8132
rect 31952 8188 32016 8192
rect 31952 8132 31956 8188
rect 31956 8132 32012 8188
rect 32012 8132 32016 8188
rect 31952 8128 32016 8132
rect 32032 8188 32096 8192
rect 32032 8132 32036 8188
rect 32036 8132 32092 8188
rect 32092 8132 32096 8188
rect 32032 8128 32096 8132
rect 32112 8188 32176 8192
rect 32112 8132 32116 8188
rect 32116 8132 32172 8188
rect 32172 8132 32176 8188
rect 32112 8128 32176 8132
rect 32192 8188 32256 8192
rect 32192 8132 32196 8188
rect 32196 8132 32252 8188
rect 32252 8132 32256 8188
rect 32192 8128 32256 8132
rect 3012 7644 3076 7648
rect 3012 7588 3016 7644
rect 3016 7588 3072 7644
rect 3072 7588 3076 7644
rect 3012 7584 3076 7588
rect 3092 7644 3156 7648
rect 3092 7588 3096 7644
rect 3096 7588 3152 7644
rect 3152 7588 3156 7644
rect 3092 7584 3156 7588
rect 3172 7644 3236 7648
rect 3172 7588 3176 7644
rect 3176 7588 3232 7644
rect 3232 7588 3236 7644
rect 3172 7584 3236 7588
rect 3252 7644 3316 7648
rect 3252 7588 3256 7644
rect 3256 7588 3312 7644
rect 3312 7588 3316 7644
rect 3252 7584 3316 7588
rect 9012 7644 9076 7648
rect 9012 7588 9016 7644
rect 9016 7588 9072 7644
rect 9072 7588 9076 7644
rect 9012 7584 9076 7588
rect 9092 7644 9156 7648
rect 9092 7588 9096 7644
rect 9096 7588 9152 7644
rect 9152 7588 9156 7644
rect 9092 7584 9156 7588
rect 9172 7644 9236 7648
rect 9172 7588 9176 7644
rect 9176 7588 9232 7644
rect 9232 7588 9236 7644
rect 9172 7584 9236 7588
rect 9252 7644 9316 7648
rect 9252 7588 9256 7644
rect 9256 7588 9312 7644
rect 9312 7588 9316 7644
rect 9252 7584 9316 7588
rect 15012 7644 15076 7648
rect 15012 7588 15016 7644
rect 15016 7588 15072 7644
rect 15072 7588 15076 7644
rect 15012 7584 15076 7588
rect 15092 7644 15156 7648
rect 15092 7588 15096 7644
rect 15096 7588 15152 7644
rect 15152 7588 15156 7644
rect 15092 7584 15156 7588
rect 15172 7644 15236 7648
rect 15172 7588 15176 7644
rect 15176 7588 15232 7644
rect 15232 7588 15236 7644
rect 15172 7584 15236 7588
rect 15252 7644 15316 7648
rect 15252 7588 15256 7644
rect 15256 7588 15312 7644
rect 15312 7588 15316 7644
rect 15252 7584 15316 7588
rect 21012 7644 21076 7648
rect 21012 7588 21016 7644
rect 21016 7588 21072 7644
rect 21072 7588 21076 7644
rect 21012 7584 21076 7588
rect 21092 7644 21156 7648
rect 21092 7588 21096 7644
rect 21096 7588 21152 7644
rect 21152 7588 21156 7644
rect 21092 7584 21156 7588
rect 21172 7644 21236 7648
rect 21172 7588 21176 7644
rect 21176 7588 21232 7644
rect 21232 7588 21236 7644
rect 21172 7584 21236 7588
rect 21252 7644 21316 7648
rect 21252 7588 21256 7644
rect 21256 7588 21312 7644
rect 21312 7588 21316 7644
rect 21252 7584 21316 7588
rect 27012 7644 27076 7648
rect 27012 7588 27016 7644
rect 27016 7588 27072 7644
rect 27072 7588 27076 7644
rect 27012 7584 27076 7588
rect 27092 7644 27156 7648
rect 27092 7588 27096 7644
rect 27096 7588 27152 7644
rect 27152 7588 27156 7644
rect 27092 7584 27156 7588
rect 27172 7644 27236 7648
rect 27172 7588 27176 7644
rect 27176 7588 27232 7644
rect 27232 7588 27236 7644
rect 27172 7584 27236 7588
rect 27252 7644 27316 7648
rect 27252 7588 27256 7644
rect 27256 7588 27312 7644
rect 27312 7588 27316 7644
rect 27252 7584 27316 7588
rect 1952 7100 2016 7104
rect 1952 7044 1956 7100
rect 1956 7044 2012 7100
rect 2012 7044 2016 7100
rect 1952 7040 2016 7044
rect 2032 7100 2096 7104
rect 2032 7044 2036 7100
rect 2036 7044 2092 7100
rect 2092 7044 2096 7100
rect 2032 7040 2096 7044
rect 2112 7100 2176 7104
rect 2112 7044 2116 7100
rect 2116 7044 2172 7100
rect 2172 7044 2176 7100
rect 2112 7040 2176 7044
rect 2192 7100 2256 7104
rect 2192 7044 2196 7100
rect 2196 7044 2252 7100
rect 2252 7044 2256 7100
rect 2192 7040 2256 7044
rect 7952 7100 8016 7104
rect 7952 7044 7956 7100
rect 7956 7044 8012 7100
rect 8012 7044 8016 7100
rect 7952 7040 8016 7044
rect 8032 7100 8096 7104
rect 8032 7044 8036 7100
rect 8036 7044 8092 7100
rect 8092 7044 8096 7100
rect 8032 7040 8096 7044
rect 8112 7100 8176 7104
rect 8112 7044 8116 7100
rect 8116 7044 8172 7100
rect 8172 7044 8176 7100
rect 8112 7040 8176 7044
rect 8192 7100 8256 7104
rect 8192 7044 8196 7100
rect 8196 7044 8252 7100
rect 8252 7044 8256 7100
rect 8192 7040 8256 7044
rect 13952 7100 14016 7104
rect 13952 7044 13956 7100
rect 13956 7044 14012 7100
rect 14012 7044 14016 7100
rect 13952 7040 14016 7044
rect 14032 7100 14096 7104
rect 14032 7044 14036 7100
rect 14036 7044 14092 7100
rect 14092 7044 14096 7100
rect 14032 7040 14096 7044
rect 14112 7100 14176 7104
rect 14112 7044 14116 7100
rect 14116 7044 14172 7100
rect 14172 7044 14176 7100
rect 14112 7040 14176 7044
rect 14192 7100 14256 7104
rect 14192 7044 14196 7100
rect 14196 7044 14252 7100
rect 14252 7044 14256 7100
rect 14192 7040 14256 7044
rect 19952 7100 20016 7104
rect 19952 7044 19956 7100
rect 19956 7044 20012 7100
rect 20012 7044 20016 7100
rect 19952 7040 20016 7044
rect 20032 7100 20096 7104
rect 20032 7044 20036 7100
rect 20036 7044 20092 7100
rect 20092 7044 20096 7100
rect 20032 7040 20096 7044
rect 20112 7100 20176 7104
rect 20112 7044 20116 7100
rect 20116 7044 20172 7100
rect 20172 7044 20176 7100
rect 20112 7040 20176 7044
rect 20192 7100 20256 7104
rect 20192 7044 20196 7100
rect 20196 7044 20252 7100
rect 20252 7044 20256 7100
rect 20192 7040 20256 7044
rect 25952 7100 26016 7104
rect 25952 7044 25956 7100
rect 25956 7044 26012 7100
rect 26012 7044 26016 7100
rect 25952 7040 26016 7044
rect 26032 7100 26096 7104
rect 26032 7044 26036 7100
rect 26036 7044 26092 7100
rect 26092 7044 26096 7100
rect 26032 7040 26096 7044
rect 26112 7100 26176 7104
rect 26112 7044 26116 7100
rect 26116 7044 26172 7100
rect 26172 7044 26176 7100
rect 26112 7040 26176 7044
rect 26192 7100 26256 7104
rect 26192 7044 26196 7100
rect 26196 7044 26252 7100
rect 26252 7044 26256 7100
rect 26192 7040 26256 7044
rect 31952 7100 32016 7104
rect 31952 7044 31956 7100
rect 31956 7044 32012 7100
rect 32012 7044 32016 7100
rect 31952 7040 32016 7044
rect 32032 7100 32096 7104
rect 32032 7044 32036 7100
rect 32036 7044 32092 7100
rect 32092 7044 32096 7100
rect 32032 7040 32096 7044
rect 32112 7100 32176 7104
rect 32112 7044 32116 7100
rect 32116 7044 32172 7100
rect 32172 7044 32176 7100
rect 32112 7040 32176 7044
rect 32192 7100 32256 7104
rect 32192 7044 32196 7100
rect 32196 7044 32252 7100
rect 32252 7044 32256 7100
rect 32192 7040 32256 7044
rect 3012 6556 3076 6560
rect 3012 6500 3016 6556
rect 3016 6500 3072 6556
rect 3072 6500 3076 6556
rect 3012 6496 3076 6500
rect 3092 6556 3156 6560
rect 3092 6500 3096 6556
rect 3096 6500 3152 6556
rect 3152 6500 3156 6556
rect 3092 6496 3156 6500
rect 3172 6556 3236 6560
rect 3172 6500 3176 6556
rect 3176 6500 3232 6556
rect 3232 6500 3236 6556
rect 3172 6496 3236 6500
rect 3252 6556 3316 6560
rect 3252 6500 3256 6556
rect 3256 6500 3312 6556
rect 3312 6500 3316 6556
rect 3252 6496 3316 6500
rect 9012 6556 9076 6560
rect 9012 6500 9016 6556
rect 9016 6500 9072 6556
rect 9072 6500 9076 6556
rect 9012 6496 9076 6500
rect 9092 6556 9156 6560
rect 9092 6500 9096 6556
rect 9096 6500 9152 6556
rect 9152 6500 9156 6556
rect 9092 6496 9156 6500
rect 9172 6556 9236 6560
rect 9172 6500 9176 6556
rect 9176 6500 9232 6556
rect 9232 6500 9236 6556
rect 9172 6496 9236 6500
rect 9252 6556 9316 6560
rect 9252 6500 9256 6556
rect 9256 6500 9312 6556
rect 9312 6500 9316 6556
rect 9252 6496 9316 6500
rect 15012 6556 15076 6560
rect 15012 6500 15016 6556
rect 15016 6500 15072 6556
rect 15072 6500 15076 6556
rect 15012 6496 15076 6500
rect 15092 6556 15156 6560
rect 15092 6500 15096 6556
rect 15096 6500 15152 6556
rect 15152 6500 15156 6556
rect 15092 6496 15156 6500
rect 15172 6556 15236 6560
rect 15172 6500 15176 6556
rect 15176 6500 15232 6556
rect 15232 6500 15236 6556
rect 15172 6496 15236 6500
rect 15252 6556 15316 6560
rect 15252 6500 15256 6556
rect 15256 6500 15312 6556
rect 15312 6500 15316 6556
rect 15252 6496 15316 6500
rect 21012 6556 21076 6560
rect 21012 6500 21016 6556
rect 21016 6500 21072 6556
rect 21072 6500 21076 6556
rect 21012 6496 21076 6500
rect 21092 6556 21156 6560
rect 21092 6500 21096 6556
rect 21096 6500 21152 6556
rect 21152 6500 21156 6556
rect 21092 6496 21156 6500
rect 21172 6556 21236 6560
rect 21172 6500 21176 6556
rect 21176 6500 21232 6556
rect 21232 6500 21236 6556
rect 21172 6496 21236 6500
rect 21252 6556 21316 6560
rect 21252 6500 21256 6556
rect 21256 6500 21312 6556
rect 21312 6500 21316 6556
rect 21252 6496 21316 6500
rect 27012 6556 27076 6560
rect 27012 6500 27016 6556
rect 27016 6500 27072 6556
rect 27072 6500 27076 6556
rect 27012 6496 27076 6500
rect 27092 6556 27156 6560
rect 27092 6500 27096 6556
rect 27096 6500 27152 6556
rect 27152 6500 27156 6556
rect 27092 6496 27156 6500
rect 27172 6556 27236 6560
rect 27172 6500 27176 6556
rect 27176 6500 27232 6556
rect 27232 6500 27236 6556
rect 27172 6496 27236 6500
rect 27252 6556 27316 6560
rect 27252 6500 27256 6556
rect 27256 6500 27312 6556
rect 27312 6500 27316 6556
rect 27252 6496 27316 6500
rect 1952 6012 2016 6016
rect 1952 5956 1956 6012
rect 1956 5956 2012 6012
rect 2012 5956 2016 6012
rect 1952 5952 2016 5956
rect 2032 6012 2096 6016
rect 2032 5956 2036 6012
rect 2036 5956 2092 6012
rect 2092 5956 2096 6012
rect 2032 5952 2096 5956
rect 2112 6012 2176 6016
rect 2112 5956 2116 6012
rect 2116 5956 2172 6012
rect 2172 5956 2176 6012
rect 2112 5952 2176 5956
rect 2192 6012 2256 6016
rect 2192 5956 2196 6012
rect 2196 5956 2252 6012
rect 2252 5956 2256 6012
rect 2192 5952 2256 5956
rect 7952 6012 8016 6016
rect 7952 5956 7956 6012
rect 7956 5956 8012 6012
rect 8012 5956 8016 6012
rect 7952 5952 8016 5956
rect 8032 6012 8096 6016
rect 8032 5956 8036 6012
rect 8036 5956 8092 6012
rect 8092 5956 8096 6012
rect 8032 5952 8096 5956
rect 8112 6012 8176 6016
rect 8112 5956 8116 6012
rect 8116 5956 8172 6012
rect 8172 5956 8176 6012
rect 8112 5952 8176 5956
rect 8192 6012 8256 6016
rect 8192 5956 8196 6012
rect 8196 5956 8252 6012
rect 8252 5956 8256 6012
rect 8192 5952 8256 5956
rect 13952 6012 14016 6016
rect 13952 5956 13956 6012
rect 13956 5956 14012 6012
rect 14012 5956 14016 6012
rect 13952 5952 14016 5956
rect 14032 6012 14096 6016
rect 14032 5956 14036 6012
rect 14036 5956 14092 6012
rect 14092 5956 14096 6012
rect 14032 5952 14096 5956
rect 14112 6012 14176 6016
rect 14112 5956 14116 6012
rect 14116 5956 14172 6012
rect 14172 5956 14176 6012
rect 14112 5952 14176 5956
rect 14192 6012 14256 6016
rect 14192 5956 14196 6012
rect 14196 5956 14252 6012
rect 14252 5956 14256 6012
rect 14192 5952 14256 5956
rect 19952 6012 20016 6016
rect 19952 5956 19956 6012
rect 19956 5956 20012 6012
rect 20012 5956 20016 6012
rect 19952 5952 20016 5956
rect 20032 6012 20096 6016
rect 20032 5956 20036 6012
rect 20036 5956 20092 6012
rect 20092 5956 20096 6012
rect 20032 5952 20096 5956
rect 20112 6012 20176 6016
rect 20112 5956 20116 6012
rect 20116 5956 20172 6012
rect 20172 5956 20176 6012
rect 20112 5952 20176 5956
rect 20192 6012 20256 6016
rect 20192 5956 20196 6012
rect 20196 5956 20252 6012
rect 20252 5956 20256 6012
rect 20192 5952 20256 5956
rect 25952 6012 26016 6016
rect 25952 5956 25956 6012
rect 25956 5956 26012 6012
rect 26012 5956 26016 6012
rect 25952 5952 26016 5956
rect 26032 6012 26096 6016
rect 26032 5956 26036 6012
rect 26036 5956 26092 6012
rect 26092 5956 26096 6012
rect 26032 5952 26096 5956
rect 26112 6012 26176 6016
rect 26112 5956 26116 6012
rect 26116 5956 26172 6012
rect 26172 5956 26176 6012
rect 26112 5952 26176 5956
rect 26192 6012 26256 6016
rect 26192 5956 26196 6012
rect 26196 5956 26252 6012
rect 26252 5956 26256 6012
rect 26192 5952 26256 5956
rect 31952 6012 32016 6016
rect 31952 5956 31956 6012
rect 31956 5956 32012 6012
rect 32012 5956 32016 6012
rect 31952 5952 32016 5956
rect 32032 6012 32096 6016
rect 32032 5956 32036 6012
rect 32036 5956 32092 6012
rect 32092 5956 32096 6012
rect 32032 5952 32096 5956
rect 32112 6012 32176 6016
rect 32112 5956 32116 6012
rect 32116 5956 32172 6012
rect 32172 5956 32176 6012
rect 32112 5952 32176 5956
rect 32192 6012 32256 6016
rect 32192 5956 32196 6012
rect 32196 5956 32252 6012
rect 32252 5956 32256 6012
rect 32192 5952 32256 5956
rect 3012 5468 3076 5472
rect 3012 5412 3016 5468
rect 3016 5412 3072 5468
rect 3072 5412 3076 5468
rect 3012 5408 3076 5412
rect 3092 5468 3156 5472
rect 3092 5412 3096 5468
rect 3096 5412 3152 5468
rect 3152 5412 3156 5468
rect 3092 5408 3156 5412
rect 3172 5468 3236 5472
rect 3172 5412 3176 5468
rect 3176 5412 3232 5468
rect 3232 5412 3236 5468
rect 3172 5408 3236 5412
rect 3252 5468 3316 5472
rect 3252 5412 3256 5468
rect 3256 5412 3312 5468
rect 3312 5412 3316 5468
rect 3252 5408 3316 5412
rect 9012 5468 9076 5472
rect 9012 5412 9016 5468
rect 9016 5412 9072 5468
rect 9072 5412 9076 5468
rect 9012 5408 9076 5412
rect 9092 5468 9156 5472
rect 9092 5412 9096 5468
rect 9096 5412 9152 5468
rect 9152 5412 9156 5468
rect 9092 5408 9156 5412
rect 9172 5468 9236 5472
rect 9172 5412 9176 5468
rect 9176 5412 9232 5468
rect 9232 5412 9236 5468
rect 9172 5408 9236 5412
rect 9252 5468 9316 5472
rect 9252 5412 9256 5468
rect 9256 5412 9312 5468
rect 9312 5412 9316 5468
rect 9252 5408 9316 5412
rect 15012 5468 15076 5472
rect 15012 5412 15016 5468
rect 15016 5412 15072 5468
rect 15072 5412 15076 5468
rect 15012 5408 15076 5412
rect 15092 5468 15156 5472
rect 15092 5412 15096 5468
rect 15096 5412 15152 5468
rect 15152 5412 15156 5468
rect 15092 5408 15156 5412
rect 15172 5468 15236 5472
rect 15172 5412 15176 5468
rect 15176 5412 15232 5468
rect 15232 5412 15236 5468
rect 15172 5408 15236 5412
rect 15252 5468 15316 5472
rect 15252 5412 15256 5468
rect 15256 5412 15312 5468
rect 15312 5412 15316 5468
rect 15252 5408 15316 5412
rect 21012 5468 21076 5472
rect 21012 5412 21016 5468
rect 21016 5412 21072 5468
rect 21072 5412 21076 5468
rect 21012 5408 21076 5412
rect 21092 5468 21156 5472
rect 21092 5412 21096 5468
rect 21096 5412 21152 5468
rect 21152 5412 21156 5468
rect 21092 5408 21156 5412
rect 21172 5468 21236 5472
rect 21172 5412 21176 5468
rect 21176 5412 21232 5468
rect 21232 5412 21236 5468
rect 21172 5408 21236 5412
rect 21252 5468 21316 5472
rect 21252 5412 21256 5468
rect 21256 5412 21312 5468
rect 21312 5412 21316 5468
rect 21252 5408 21316 5412
rect 27012 5468 27076 5472
rect 27012 5412 27016 5468
rect 27016 5412 27072 5468
rect 27072 5412 27076 5468
rect 27012 5408 27076 5412
rect 27092 5468 27156 5472
rect 27092 5412 27096 5468
rect 27096 5412 27152 5468
rect 27152 5412 27156 5468
rect 27092 5408 27156 5412
rect 27172 5468 27236 5472
rect 27172 5412 27176 5468
rect 27176 5412 27232 5468
rect 27232 5412 27236 5468
rect 27172 5408 27236 5412
rect 27252 5468 27316 5472
rect 27252 5412 27256 5468
rect 27256 5412 27312 5468
rect 27312 5412 27316 5468
rect 27252 5408 27316 5412
rect 1952 4924 2016 4928
rect 1952 4868 1956 4924
rect 1956 4868 2012 4924
rect 2012 4868 2016 4924
rect 1952 4864 2016 4868
rect 2032 4924 2096 4928
rect 2032 4868 2036 4924
rect 2036 4868 2092 4924
rect 2092 4868 2096 4924
rect 2032 4864 2096 4868
rect 2112 4924 2176 4928
rect 2112 4868 2116 4924
rect 2116 4868 2172 4924
rect 2172 4868 2176 4924
rect 2112 4864 2176 4868
rect 2192 4924 2256 4928
rect 2192 4868 2196 4924
rect 2196 4868 2252 4924
rect 2252 4868 2256 4924
rect 2192 4864 2256 4868
rect 7952 4924 8016 4928
rect 7952 4868 7956 4924
rect 7956 4868 8012 4924
rect 8012 4868 8016 4924
rect 7952 4864 8016 4868
rect 8032 4924 8096 4928
rect 8032 4868 8036 4924
rect 8036 4868 8092 4924
rect 8092 4868 8096 4924
rect 8032 4864 8096 4868
rect 8112 4924 8176 4928
rect 8112 4868 8116 4924
rect 8116 4868 8172 4924
rect 8172 4868 8176 4924
rect 8112 4864 8176 4868
rect 8192 4924 8256 4928
rect 8192 4868 8196 4924
rect 8196 4868 8252 4924
rect 8252 4868 8256 4924
rect 8192 4864 8256 4868
rect 13952 4924 14016 4928
rect 13952 4868 13956 4924
rect 13956 4868 14012 4924
rect 14012 4868 14016 4924
rect 13952 4864 14016 4868
rect 14032 4924 14096 4928
rect 14032 4868 14036 4924
rect 14036 4868 14092 4924
rect 14092 4868 14096 4924
rect 14032 4864 14096 4868
rect 14112 4924 14176 4928
rect 14112 4868 14116 4924
rect 14116 4868 14172 4924
rect 14172 4868 14176 4924
rect 14112 4864 14176 4868
rect 14192 4924 14256 4928
rect 14192 4868 14196 4924
rect 14196 4868 14252 4924
rect 14252 4868 14256 4924
rect 14192 4864 14256 4868
rect 19952 4924 20016 4928
rect 19952 4868 19956 4924
rect 19956 4868 20012 4924
rect 20012 4868 20016 4924
rect 19952 4864 20016 4868
rect 20032 4924 20096 4928
rect 20032 4868 20036 4924
rect 20036 4868 20092 4924
rect 20092 4868 20096 4924
rect 20032 4864 20096 4868
rect 20112 4924 20176 4928
rect 20112 4868 20116 4924
rect 20116 4868 20172 4924
rect 20172 4868 20176 4924
rect 20112 4864 20176 4868
rect 20192 4924 20256 4928
rect 20192 4868 20196 4924
rect 20196 4868 20252 4924
rect 20252 4868 20256 4924
rect 20192 4864 20256 4868
rect 25952 4924 26016 4928
rect 25952 4868 25956 4924
rect 25956 4868 26012 4924
rect 26012 4868 26016 4924
rect 25952 4864 26016 4868
rect 26032 4924 26096 4928
rect 26032 4868 26036 4924
rect 26036 4868 26092 4924
rect 26092 4868 26096 4924
rect 26032 4864 26096 4868
rect 26112 4924 26176 4928
rect 26112 4868 26116 4924
rect 26116 4868 26172 4924
rect 26172 4868 26176 4924
rect 26112 4864 26176 4868
rect 26192 4924 26256 4928
rect 26192 4868 26196 4924
rect 26196 4868 26252 4924
rect 26252 4868 26256 4924
rect 26192 4864 26256 4868
rect 31952 4924 32016 4928
rect 31952 4868 31956 4924
rect 31956 4868 32012 4924
rect 32012 4868 32016 4924
rect 31952 4864 32016 4868
rect 32032 4924 32096 4928
rect 32032 4868 32036 4924
rect 32036 4868 32092 4924
rect 32092 4868 32096 4924
rect 32032 4864 32096 4868
rect 32112 4924 32176 4928
rect 32112 4868 32116 4924
rect 32116 4868 32172 4924
rect 32172 4868 32176 4924
rect 32112 4864 32176 4868
rect 32192 4924 32256 4928
rect 32192 4868 32196 4924
rect 32196 4868 32252 4924
rect 32252 4868 32256 4924
rect 32192 4864 32256 4868
rect 3012 4380 3076 4384
rect 3012 4324 3016 4380
rect 3016 4324 3072 4380
rect 3072 4324 3076 4380
rect 3012 4320 3076 4324
rect 3092 4380 3156 4384
rect 3092 4324 3096 4380
rect 3096 4324 3152 4380
rect 3152 4324 3156 4380
rect 3092 4320 3156 4324
rect 3172 4380 3236 4384
rect 3172 4324 3176 4380
rect 3176 4324 3232 4380
rect 3232 4324 3236 4380
rect 3172 4320 3236 4324
rect 3252 4380 3316 4384
rect 3252 4324 3256 4380
rect 3256 4324 3312 4380
rect 3312 4324 3316 4380
rect 3252 4320 3316 4324
rect 9012 4380 9076 4384
rect 9012 4324 9016 4380
rect 9016 4324 9072 4380
rect 9072 4324 9076 4380
rect 9012 4320 9076 4324
rect 9092 4380 9156 4384
rect 9092 4324 9096 4380
rect 9096 4324 9152 4380
rect 9152 4324 9156 4380
rect 9092 4320 9156 4324
rect 9172 4380 9236 4384
rect 9172 4324 9176 4380
rect 9176 4324 9232 4380
rect 9232 4324 9236 4380
rect 9172 4320 9236 4324
rect 9252 4380 9316 4384
rect 9252 4324 9256 4380
rect 9256 4324 9312 4380
rect 9312 4324 9316 4380
rect 9252 4320 9316 4324
rect 15012 4380 15076 4384
rect 15012 4324 15016 4380
rect 15016 4324 15072 4380
rect 15072 4324 15076 4380
rect 15012 4320 15076 4324
rect 15092 4380 15156 4384
rect 15092 4324 15096 4380
rect 15096 4324 15152 4380
rect 15152 4324 15156 4380
rect 15092 4320 15156 4324
rect 15172 4380 15236 4384
rect 15172 4324 15176 4380
rect 15176 4324 15232 4380
rect 15232 4324 15236 4380
rect 15172 4320 15236 4324
rect 15252 4380 15316 4384
rect 15252 4324 15256 4380
rect 15256 4324 15312 4380
rect 15312 4324 15316 4380
rect 15252 4320 15316 4324
rect 21012 4380 21076 4384
rect 21012 4324 21016 4380
rect 21016 4324 21072 4380
rect 21072 4324 21076 4380
rect 21012 4320 21076 4324
rect 21092 4380 21156 4384
rect 21092 4324 21096 4380
rect 21096 4324 21152 4380
rect 21152 4324 21156 4380
rect 21092 4320 21156 4324
rect 21172 4380 21236 4384
rect 21172 4324 21176 4380
rect 21176 4324 21232 4380
rect 21232 4324 21236 4380
rect 21172 4320 21236 4324
rect 21252 4380 21316 4384
rect 21252 4324 21256 4380
rect 21256 4324 21312 4380
rect 21312 4324 21316 4380
rect 21252 4320 21316 4324
rect 27012 4380 27076 4384
rect 27012 4324 27016 4380
rect 27016 4324 27072 4380
rect 27072 4324 27076 4380
rect 27012 4320 27076 4324
rect 27092 4380 27156 4384
rect 27092 4324 27096 4380
rect 27096 4324 27152 4380
rect 27152 4324 27156 4380
rect 27092 4320 27156 4324
rect 27172 4380 27236 4384
rect 27172 4324 27176 4380
rect 27176 4324 27232 4380
rect 27232 4324 27236 4380
rect 27172 4320 27236 4324
rect 27252 4380 27316 4384
rect 27252 4324 27256 4380
rect 27256 4324 27312 4380
rect 27312 4324 27316 4380
rect 27252 4320 27316 4324
rect 1952 3836 2016 3840
rect 1952 3780 1956 3836
rect 1956 3780 2012 3836
rect 2012 3780 2016 3836
rect 1952 3776 2016 3780
rect 2032 3836 2096 3840
rect 2032 3780 2036 3836
rect 2036 3780 2092 3836
rect 2092 3780 2096 3836
rect 2032 3776 2096 3780
rect 2112 3836 2176 3840
rect 2112 3780 2116 3836
rect 2116 3780 2172 3836
rect 2172 3780 2176 3836
rect 2112 3776 2176 3780
rect 2192 3836 2256 3840
rect 2192 3780 2196 3836
rect 2196 3780 2252 3836
rect 2252 3780 2256 3836
rect 2192 3776 2256 3780
rect 7952 3836 8016 3840
rect 7952 3780 7956 3836
rect 7956 3780 8012 3836
rect 8012 3780 8016 3836
rect 7952 3776 8016 3780
rect 8032 3836 8096 3840
rect 8032 3780 8036 3836
rect 8036 3780 8092 3836
rect 8092 3780 8096 3836
rect 8032 3776 8096 3780
rect 8112 3836 8176 3840
rect 8112 3780 8116 3836
rect 8116 3780 8172 3836
rect 8172 3780 8176 3836
rect 8112 3776 8176 3780
rect 8192 3836 8256 3840
rect 8192 3780 8196 3836
rect 8196 3780 8252 3836
rect 8252 3780 8256 3836
rect 8192 3776 8256 3780
rect 13952 3836 14016 3840
rect 13952 3780 13956 3836
rect 13956 3780 14012 3836
rect 14012 3780 14016 3836
rect 13952 3776 14016 3780
rect 14032 3836 14096 3840
rect 14032 3780 14036 3836
rect 14036 3780 14092 3836
rect 14092 3780 14096 3836
rect 14032 3776 14096 3780
rect 14112 3836 14176 3840
rect 14112 3780 14116 3836
rect 14116 3780 14172 3836
rect 14172 3780 14176 3836
rect 14112 3776 14176 3780
rect 14192 3836 14256 3840
rect 14192 3780 14196 3836
rect 14196 3780 14252 3836
rect 14252 3780 14256 3836
rect 14192 3776 14256 3780
rect 19952 3836 20016 3840
rect 19952 3780 19956 3836
rect 19956 3780 20012 3836
rect 20012 3780 20016 3836
rect 19952 3776 20016 3780
rect 20032 3836 20096 3840
rect 20032 3780 20036 3836
rect 20036 3780 20092 3836
rect 20092 3780 20096 3836
rect 20032 3776 20096 3780
rect 20112 3836 20176 3840
rect 20112 3780 20116 3836
rect 20116 3780 20172 3836
rect 20172 3780 20176 3836
rect 20112 3776 20176 3780
rect 20192 3836 20256 3840
rect 20192 3780 20196 3836
rect 20196 3780 20252 3836
rect 20252 3780 20256 3836
rect 20192 3776 20256 3780
rect 25952 3836 26016 3840
rect 25952 3780 25956 3836
rect 25956 3780 26012 3836
rect 26012 3780 26016 3836
rect 25952 3776 26016 3780
rect 26032 3836 26096 3840
rect 26032 3780 26036 3836
rect 26036 3780 26092 3836
rect 26092 3780 26096 3836
rect 26032 3776 26096 3780
rect 26112 3836 26176 3840
rect 26112 3780 26116 3836
rect 26116 3780 26172 3836
rect 26172 3780 26176 3836
rect 26112 3776 26176 3780
rect 26192 3836 26256 3840
rect 26192 3780 26196 3836
rect 26196 3780 26252 3836
rect 26252 3780 26256 3836
rect 26192 3776 26256 3780
rect 31952 3836 32016 3840
rect 31952 3780 31956 3836
rect 31956 3780 32012 3836
rect 32012 3780 32016 3836
rect 31952 3776 32016 3780
rect 32032 3836 32096 3840
rect 32032 3780 32036 3836
rect 32036 3780 32092 3836
rect 32092 3780 32096 3836
rect 32032 3776 32096 3780
rect 32112 3836 32176 3840
rect 32112 3780 32116 3836
rect 32116 3780 32172 3836
rect 32172 3780 32176 3836
rect 32112 3776 32176 3780
rect 32192 3836 32256 3840
rect 32192 3780 32196 3836
rect 32196 3780 32252 3836
rect 32252 3780 32256 3836
rect 32192 3776 32256 3780
rect 3012 3292 3076 3296
rect 3012 3236 3016 3292
rect 3016 3236 3072 3292
rect 3072 3236 3076 3292
rect 3012 3232 3076 3236
rect 3092 3292 3156 3296
rect 3092 3236 3096 3292
rect 3096 3236 3152 3292
rect 3152 3236 3156 3292
rect 3092 3232 3156 3236
rect 3172 3292 3236 3296
rect 3172 3236 3176 3292
rect 3176 3236 3232 3292
rect 3232 3236 3236 3292
rect 3172 3232 3236 3236
rect 3252 3292 3316 3296
rect 3252 3236 3256 3292
rect 3256 3236 3312 3292
rect 3312 3236 3316 3292
rect 3252 3232 3316 3236
rect 9012 3292 9076 3296
rect 9012 3236 9016 3292
rect 9016 3236 9072 3292
rect 9072 3236 9076 3292
rect 9012 3232 9076 3236
rect 9092 3292 9156 3296
rect 9092 3236 9096 3292
rect 9096 3236 9152 3292
rect 9152 3236 9156 3292
rect 9092 3232 9156 3236
rect 9172 3292 9236 3296
rect 9172 3236 9176 3292
rect 9176 3236 9232 3292
rect 9232 3236 9236 3292
rect 9172 3232 9236 3236
rect 9252 3292 9316 3296
rect 9252 3236 9256 3292
rect 9256 3236 9312 3292
rect 9312 3236 9316 3292
rect 9252 3232 9316 3236
rect 15012 3292 15076 3296
rect 15012 3236 15016 3292
rect 15016 3236 15072 3292
rect 15072 3236 15076 3292
rect 15012 3232 15076 3236
rect 15092 3292 15156 3296
rect 15092 3236 15096 3292
rect 15096 3236 15152 3292
rect 15152 3236 15156 3292
rect 15092 3232 15156 3236
rect 15172 3292 15236 3296
rect 15172 3236 15176 3292
rect 15176 3236 15232 3292
rect 15232 3236 15236 3292
rect 15172 3232 15236 3236
rect 15252 3292 15316 3296
rect 15252 3236 15256 3292
rect 15256 3236 15312 3292
rect 15312 3236 15316 3292
rect 15252 3232 15316 3236
rect 21012 3292 21076 3296
rect 21012 3236 21016 3292
rect 21016 3236 21072 3292
rect 21072 3236 21076 3292
rect 21012 3232 21076 3236
rect 21092 3292 21156 3296
rect 21092 3236 21096 3292
rect 21096 3236 21152 3292
rect 21152 3236 21156 3292
rect 21092 3232 21156 3236
rect 21172 3292 21236 3296
rect 21172 3236 21176 3292
rect 21176 3236 21232 3292
rect 21232 3236 21236 3292
rect 21172 3232 21236 3236
rect 21252 3292 21316 3296
rect 21252 3236 21256 3292
rect 21256 3236 21312 3292
rect 21312 3236 21316 3292
rect 21252 3232 21316 3236
rect 27012 3292 27076 3296
rect 27012 3236 27016 3292
rect 27016 3236 27072 3292
rect 27072 3236 27076 3292
rect 27012 3232 27076 3236
rect 27092 3292 27156 3296
rect 27092 3236 27096 3292
rect 27096 3236 27152 3292
rect 27152 3236 27156 3292
rect 27092 3232 27156 3236
rect 27172 3292 27236 3296
rect 27172 3236 27176 3292
rect 27176 3236 27232 3292
rect 27232 3236 27236 3292
rect 27172 3232 27236 3236
rect 27252 3292 27316 3296
rect 27252 3236 27256 3292
rect 27256 3236 27312 3292
rect 27312 3236 27316 3292
rect 27252 3232 27316 3236
rect 1952 2748 2016 2752
rect 1952 2692 1956 2748
rect 1956 2692 2012 2748
rect 2012 2692 2016 2748
rect 1952 2688 2016 2692
rect 2032 2748 2096 2752
rect 2032 2692 2036 2748
rect 2036 2692 2092 2748
rect 2092 2692 2096 2748
rect 2032 2688 2096 2692
rect 2112 2748 2176 2752
rect 2112 2692 2116 2748
rect 2116 2692 2172 2748
rect 2172 2692 2176 2748
rect 2112 2688 2176 2692
rect 2192 2748 2256 2752
rect 2192 2692 2196 2748
rect 2196 2692 2252 2748
rect 2252 2692 2256 2748
rect 2192 2688 2256 2692
rect 7952 2748 8016 2752
rect 7952 2692 7956 2748
rect 7956 2692 8012 2748
rect 8012 2692 8016 2748
rect 7952 2688 8016 2692
rect 8032 2748 8096 2752
rect 8032 2692 8036 2748
rect 8036 2692 8092 2748
rect 8092 2692 8096 2748
rect 8032 2688 8096 2692
rect 8112 2748 8176 2752
rect 8112 2692 8116 2748
rect 8116 2692 8172 2748
rect 8172 2692 8176 2748
rect 8112 2688 8176 2692
rect 8192 2748 8256 2752
rect 8192 2692 8196 2748
rect 8196 2692 8252 2748
rect 8252 2692 8256 2748
rect 8192 2688 8256 2692
rect 13952 2748 14016 2752
rect 13952 2692 13956 2748
rect 13956 2692 14012 2748
rect 14012 2692 14016 2748
rect 13952 2688 14016 2692
rect 14032 2748 14096 2752
rect 14032 2692 14036 2748
rect 14036 2692 14092 2748
rect 14092 2692 14096 2748
rect 14032 2688 14096 2692
rect 14112 2748 14176 2752
rect 14112 2692 14116 2748
rect 14116 2692 14172 2748
rect 14172 2692 14176 2748
rect 14112 2688 14176 2692
rect 14192 2748 14256 2752
rect 14192 2692 14196 2748
rect 14196 2692 14252 2748
rect 14252 2692 14256 2748
rect 14192 2688 14256 2692
rect 19952 2748 20016 2752
rect 19952 2692 19956 2748
rect 19956 2692 20012 2748
rect 20012 2692 20016 2748
rect 19952 2688 20016 2692
rect 20032 2748 20096 2752
rect 20032 2692 20036 2748
rect 20036 2692 20092 2748
rect 20092 2692 20096 2748
rect 20032 2688 20096 2692
rect 20112 2748 20176 2752
rect 20112 2692 20116 2748
rect 20116 2692 20172 2748
rect 20172 2692 20176 2748
rect 20112 2688 20176 2692
rect 20192 2748 20256 2752
rect 20192 2692 20196 2748
rect 20196 2692 20252 2748
rect 20252 2692 20256 2748
rect 20192 2688 20256 2692
rect 25952 2748 26016 2752
rect 25952 2692 25956 2748
rect 25956 2692 26012 2748
rect 26012 2692 26016 2748
rect 25952 2688 26016 2692
rect 26032 2748 26096 2752
rect 26032 2692 26036 2748
rect 26036 2692 26092 2748
rect 26092 2692 26096 2748
rect 26032 2688 26096 2692
rect 26112 2748 26176 2752
rect 26112 2692 26116 2748
rect 26116 2692 26172 2748
rect 26172 2692 26176 2748
rect 26112 2688 26176 2692
rect 26192 2748 26256 2752
rect 26192 2692 26196 2748
rect 26196 2692 26252 2748
rect 26252 2692 26256 2748
rect 26192 2688 26256 2692
rect 31952 2748 32016 2752
rect 31952 2692 31956 2748
rect 31956 2692 32012 2748
rect 32012 2692 32016 2748
rect 31952 2688 32016 2692
rect 32032 2748 32096 2752
rect 32032 2692 32036 2748
rect 32036 2692 32092 2748
rect 32092 2692 32096 2748
rect 32032 2688 32096 2692
rect 32112 2748 32176 2752
rect 32112 2692 32116 2748
rect 32116 2692 32172 2748
rect 32172 2692 32176 2748
rect 32112 2688 32176 2692
rect 32192 2748 32256 2752
rect 32192 2692 32196 2748
rect 32196 2692 32252 2748
rect 32252 2692 32256 2748
rect 32192 2688 32256 2692
rect 3012 2204 3076 2208
rect 3012 2148 3016 2204
rect 3016 2148 3072 2204
rect 3072 2148 3076 2204
rect 3012 2144 3076 2148
rect 3092 2204 3156 2208
rect 3092 2148 3096 2204
rect 3096 2148 3152 2204
rect 3152 2148 3156 2204
rect 3092 2144 3156 2148
rect 3172 2204 3236 2208
rect 3172 2148 3176 2204
rect 3176 2148 3232 2204
rect 3232 2148 3236 2204
rect 3172 2144 3236 2148
rect 3252 2204 3316 2208
rect 3252 2148 3256 2204
rect 3256 2148 3312 2204
rect 3312 2148 3316 2204
rect 3252 2144 3316 2148
rect 9012 2204 9076 2208
rect 9012 2148 9016 2204
rect 9016 2148 9072 2204
rect 9072 2148 9076 2204
rect 9012 2144 9076 2148
rect 9092 2204 9156 2208
rect 9092 2148 9096 2204
rect 9096 2148 9152 2204
rect 9152 2148 9156 2204
rect 9092 2144 9156 2148
rect 9172 2204 9236 2208
rect 9172 2148 9176 2204
rect 9176 2148 9232 2204
rect 9232 2148 9236 2204
rect 9172 2144 9236 2148
rect 9252 2204 9316 2208
rect 9252 2148 9256 2204
rect 9256 2148 9312 2204
rect 9312 2148 9316 2204
rect 9252 2144 9316 2148
rect 15012 2204 15076 2208
rect 15012 2148 15016 2204
rect 15016 2148 15072 2204
rect 15072 2148 15076 2204
rect 15012 2144 15076 2148
rect 15092 2204 15156 2208
rect 15092 2148 15096 2204
rect 15096 2148 15152 2204
rect 15152 2148 15156 2204
rect 15092 2144 15156 2148
rect 15172 2204 15236 2208
rect 15172 2148 15176 2204
rect 15176 2148 15232 2204
rect 15232 2148 15236 2204
rect 15172 2144 15236 2148
rect 15252 2204 15316 2208
rect 15252 2148 15256 2204
rect 15256 2148 15312 2204
rect 15312 2148 15316 2204
rect 15252 2144 15316 2148
rect 21012 2204 21076 2208
rect 21012 2148 21016 2204
rect 21016 2148 21072 2204
rect 21072 2148 21076 2204
rect 21012 2144 21076 2148
rect 21092 2204 21156 2208
rect 21092 2148 21096 2204
rect 21096 2148 21152 2204
rect 21152 2148 21156 2204
rect 21092 2144 21156 2148
rect 21172 2204 21236 2208
rect 21172 2148 21176 2204
rect 21176 2148 21232 2204
rect 21232 2148 21236 2204
rect 21172 2144 21236 2148
rect 21252 2204 21316 2208
rect 21252 2148 21256 2204
rect 21256 2148 21312 2204
rect 21312 2148 21316 2204
rect 21252 2144 21316 2148
rect 27012 2204 27076 2208
rect 27012 2148 27016 2204
rect 27016 2148 27072 2204
rect 27072 2148 27076 2204
rect 27012 2144 27076 2148
rect 27092 2204 27156 2208
rect 27092 2148 27096 2204
rect 27096 2148 27152 2204
rect 27152 2148 27156 2204
rect 27092 2144 27156 2148
rect 27172 2204 27236 2208
rect 27172 2148 27176 2204
rect 27176 2148 27232 2204
rect 27232 2148 27236 2204
rect 27172 2144 27236 2148
rect 27252 2204 27316 2208
rect 27252 2148 27256 2204
rect 27256 2148 27312 2204
rect 27312 2148 27316 2204
rect 27252 2144 27316 2148
<< metal4 >>
rect 1944 8192 2264 11250
rect 1944 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2264 8192
rect 1944 7104 2264 8128
rect 1944 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2264 7104
rect 1944 6016 2264 7040
rect 1944 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2264 6016
rect 1944 4928 2264 5952
rect 1944 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2264 4928
rect 1944 3840 2264 4864
rect 1944 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2264 3840
rect 1944 2752 2264 3776
rect 1944 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2264 2752
rect 1944 0 2264 2688
rect 3004 8736 3324 11250
rect 3004 8672 3012 8736
rect 3076 8672 3092 8736
rect 3156 8672 3172 8736
rect 3236 8672 3252 8736
rect 3316 8672 3324 8736
rect 3004 7648 3324 8672
rect 3004 7584 3012 7648
rect 3076 7584 3092 7648
rect 3156 7584 3172 7648
rect 3236 7584 3252 7648
rect 3316 7584 3324 7648
rect 3004 6560 3324 7584
rect 3004 6496 3012 6560
rect 3076 6496 3092 6560
rect 3156 6496 3172 6560
rect 3236 6496 3252 6560
rect 3316 6496 3324 6560
rect 3004 5472 3324 6496
rect 3004 5408 3012 5472
rect 3076 5408 3092 5472
rect 3156 5408 3172 5472
rect 3236 5408 3252 5472
rect 3316 5408 3324 5472
rect 3004 4384 3324 5408
rect 3004 4320 3012 4384
rect 3076 4320 3092 4384
rect 3156 4320 3172 4384
rect 3236 4320 3252 4384
rect 3316 4320 3324 4384
rect 3004 3296 3324 4320
rect 3004 3232 3012 3296
rect 3076 3232 3092 3296
rect 3156 3232 3172 3296
rect 3236 3232 3252 3296
rect 3316 3232 3324 3296
rect 3004 2208 3324 3232
rect 3004 2144 3012 2208
rect 3076 2144 3092 2208
rect 3156 2144 3172 2208
rect 3236 2144 3252 2208
rect 3316 2144 3324 2208
rect 3004 0 3324 2144
rect 7944 8192 8264 11250
rect 7944 8128 7952 8192
rect 8016 8128 8032 8192
rect 8096 8128 8112 8192
rect 8176 8128 8192 8192
rect 8256 8128 8264 8192
rect 7944 7104 8264 8128
rect 7944 7040 7952 7104
rect 8016 7040 8032 7104
rect 8096 7040 8112 7104
rect 8176 7040 8192 7104
rect 8256 7040 8264 7104
rect 7944 6016 8264 7040
rect 7944 5952 7952 6016
rect 8016 5952 8032 6016
rect 8096 5952 8112 6016
rect 8176 5952 8192 6016
rect 8256 5952 8264 6016
rect 7944 4928 8264 5952
rect 7944 4864 7952 4928
rect 8016 4864 8032 4928
rect 8096 4864 8112 4928
rect 8176 4864 8192 4928
rect 8256 4864 8264 4928
rect 7944 3840 8264 4864
rect 7944 3776 7952 3840
rect 8016 3776 8032 3840
rect 8096 3776 8112 3840
rect 8176 3776 8192 3840
rect 8256 3776 8264 3840
rect 7944 2752 8264 3776
rect 7944 2688 7952 2752
rect 8016 2688 8032 2752
rect 8096 2688 8112 2752
rect 8176 2688 8192 2752
rect 8256 2688 8264 2752
rect 7944 0 8264 2688
rect 9004 8736 9324 11250
rect 9004 8672 9012 8736
rect 9076 8672 9092 8736
rect 9156 8672 9172 8736
rect 9236 8672 9252 8736
rect 9316 8672 9324 8736
rect 9004 7648 9324 8672
rect 9004 7584 9012 7648
rect 9076 7584 9092 7648
rect 9156 7584 9172 7648
rect 9236 7584 9252 7648
rect 9316 7584 9324 7648
rect 9004 6560 9324 7584
rect 9004 6496 9012 6560
rect 9076 6496 9092 6560
rect 9156 6496 9172 6560
rect 9236 6496 9252 6560
rect 9316 6496 9324 6560
rect 9004 5472 9324 6496
rect 9004 5408 9012 5472
rect 9076 5408 9092 5472
rect 9156 5408 9172 5472
rect 9236 5408 9252 5472
rect 9316 5408 9324 5472
rect 9004 4384 9324 5408
rect 9004 4320 9012 4384
rect 9076 4320 9092 4384
rect 9156 4320 9172 4384
rect 9236 4320 9252 4384
rect 9316 4320 9324 4384
rect 9004 3296 9324 4320
rect 9004 3232 9012 3296
rect 9076 3232 9092 3296
rect 9156 3232 9172 3296
rect 9236 3232 9252 3296
rect 9316 3232 9324 3296
rect 9004 2208 9324 3232
rect 9004 2144 9012 2208
rect 9076 2144 9092 2208
rect 9156 2144 9172 2208
rect 9236 2144 9252 2208
rect 9316 2144 9324 2208
rect 9004 0 9324 2144
rect 13944 8192 14264 11250
rect 13944 8128 13952 8192
rect 14016 8128 14032 8192
rect 14096 8128 14112 8192
rect 14176 8128 14192 8192
rect 14256 8128 14264 8192
rect 13944 7104 14264 8128
rect 13944 7040 13952 7104
rect 14016 7040 14032 7104
rect 14096 7040 14112 7104
rect 14176 7040 14192 7104
rect 14256 7040 14264 7104
rect 13944 6016 14264 7040
rect 13944 5952 13952 6016
rect 14016 5952 14032 6016
rect 14096 5952 14112 6016
rect 14176 5952 14192 6016
rect 14256 5952 14264 6016
rect 13944 4928 14264 5952
rect 13944 4864 13952 4928
rect 14016 4864 14032 4928
rect 14096 4864 14112 4928
rect 14176 4864 14192 4928
rect 14256 4864 14264 4928
rect 13944 3840 14264 4864
rect 13944 3776 13952 3840
rect 14016 3776 14032 3840
rect 14096 3776 14112 3840
rect 14176 3776 14192 3840
rect 14256 3776 14264 3840
rect 13944 2752 14264 3776
rect 13944 2688 13952 2752
rect 14016 2688 14032 2752
rect 14096 2688 14112 2752
rect 14176 2688 14192 2752
rect 14256 2688 14264 2752
rect 13944 0 14264 2688
rect 15004 8736 15324 11250
rect 15004 8672 15012 8736
rect 15076 8672 15092 8736
rect 15156 8672 15172 8736
rect 15236 8672 15252 8736
rect 15316 8672 15324 8736
rect 15004 7648 15324 8672
rect 15004 7584 15012 7648
rect 15076 7584 15092 7648
rect 15156 7584 15172 7648
rect 15236 7584 15252 7648
rect 15316 7584 15324 7648
rect 15004 6560 15324 7584
rect 15004 6496 15012 6560
rect 15076 6496 15092 6560
rect 15156 6496 15172 6560
rect 15236 6496 15252 6560
rect 15316 6496 15324 6560
rect 15004 5472 15324 6496
rect 15004 5408 15012 5472
rect 15076 5408 15092 5472
rect 15156 5408 15172 5472
rect 15236 5408 15252 5472
rect 15316 5408 15324 5472
rect 15004 4384 15324 5408
rect 15004 4320 15012 4384
rect 15076 4320 15092 4384
rect 15156 4320 15172 4384
rect 15236 4320 15252 4384
rect 15316 4320 15324 4384
rect 15004 3296 15324 4320
rect 15004 3232 15012 3296
rect 15076 3232 15092 3296
rect 15156 3232 15172 3296
rect 15236 3232 15252 3296
rect 15316 3232 15324 3296
rect 15004 2208 15324 3232
rect 15004 2144 15012 2208
rect 15076 2144 15092 2208
rect 15156 2144 15172 2208
rect 15236 2144 15252 2208
rect 15316 2144 15324 2208
rect 15004 0 15324 2144
rect 19944 8192 20264 11250
rect 19944 8128 19952 8192
rect 20016 8128 20032 8192
rect 20096 8128 20112 8192
rect 20176 8128 20192 8192
rect 20256 8128 20264 8192
rect 19944 7104 20264 8128
rect 19944 7040 19952 7104
rect 20016 7040 20032 7104
rect 20096 7040 20112 7104
rect 20176 7040 20192 7104
rect 20256 7040 20264 7104
rect 19944 6016 20264 7040
rect 19944 5952 19952 6016
rect 20016 5952 20032 6016
rect 20096 5952 20112 6016
rect 20176 5952 20192 6016
rect 20256 5952 20264 6016
rect 19944 4928 20264 5952
rect 19944 4864 19952 4928
rect 20016 4864 20032 4928
rect 20096 4864 20112 4928
rect 20176 4864 20192 4928
rect 20256 4864 20264 4928
rect 19944 3840 20264 4864
rect 19944 3776 19952 3840
rect 20016 3776 20032 3840
rect 20096 3776 20112 3840
rect 20176 3776 20192 3840
rect 20256 3776 20264 3840
rect 19944 2752 20264 3776
rect 19944 2688 19952 2752
rect 20016 2688 20032 2752
rect 20096 2688 20112 2752
rect 20176 2688 20192 2752
rect 20256 2688 20264 2752
rect 19944 0 20264 2688
rect 21004 8736 21324 11250
rect 21004 8672 21012 8736
rect 21076 8672 21092 8736
rect 21156 8672 21172 8736
rect 21236 8672 21252 8736
rect 21316 8672 21324 8736
rect 21004 7648 21324 8672
rect 21004 7584 21012 7648
rect 21076 7584 21092 7648
rect 21156 7584 21172 7648
rect 21236 7584 21252 7648
rect 21316 7584 21324 7648
rect 21004 6560 21324 7584
rect 21004 6496 21012 6560
rect 21076 6496 21092 6560
rect 21156 6496 21172 6560
rect 21236 6496 21252 6560
rect 21316 6496 21324 6560
rect 21004 5472 21324 6496
rect 21004 5408 21012 5472
rect 21076 5408 21092 5472
rect 21156 5408 21172 5472
rect 21236 5408 21252 5472
rect 21316 5408 21324 5472
rect 21004 4384 21324 5408
rect 21004 4320 21012 4384
rect 21076 4320 21092 4384
rect 21156 4320 21172 4384
rect 21236 4320 21252 4384
rect 21316 4320 21324 4384
rect 21004 3296 21324 4320
rect 21004 3232 21012 3296
rect 21076 3232 21092 3296
rect 21156 3232 21172 3296
rect 21236 3232 21252 3296
rect 21316 3232 21324 3296
rect 21004 2208 21324 3232
rect 21004 2144 21012 2208
rect 21076 2144 21092 2208
rect 21156 2144 21172 2208
rect 21236 2144 21252 2208
rect 21316 2144 21324 2208
rect 21004 0 21324 2144
rect 25944 8192 26264 11250
rect 25944 8128 25952 8192
rect 26016 8128 26032 8192
rect 26096 8128 26112 8192
rect 26176 8128 26192 8192
rect 26256 8128 26264 8192
rect 25944 7104 26264 8128
rect 25944 7040 25952 7104
rect 26016 7040 26032 7104
rect 26096 7040 26112 7104
rect 26176 7040 26192 7104
rect 26256 7040 26264 7104
rect 25944 6016 26264 7040
rect 25944 5952 25952 6016
rect 26016 5952 26032 6016
rect 26096 5952 26112 6016
rect 26176 5952 26192 6016
rect 26256 5952 26264 6016
rect 25944 4928 26264 5952
rect 25944 4864 25952 4928
rect 26016 4864 26032 4928
rect 26096 4864 26112 4928
rect 26176 4864 26192 4928
rect 26256 4864 26264 4928
rect 25944 3840 26264 4864
rect 25944 3776 25952 3840
rect 26016 3776 26032 3840
rect 26096 3776 26112 3840
rect 26176 3776 26192 3840
rect 26256 3776 26264 3840
rect 25944 2752 26264 3776
rect 25944 2688 25952 2752
rect 26016 2688 26032 2752
rect 26096 2688 26112 2752
rect 26176 2688 26192 2752
rect 26256 2688 26264 2752
rect 25944 0 26264 2688
rect 27004 8736 27324 11250
rect 27004 8672 27012 8736
rect 27076 8672 27092 8736
rect 27156 8672 27172 8736
rect 27236 8672 27252 8736
rect 27316 8672 27324 8736
rect 27004 7648 27324 8672
rect 27004 7584 27012 7648
rect 27076 7584 27092 7648
rect 27156 7584 27172 7648
rect 27236 7584 27252 7648
rect 27316 7584 27324 7648
rect 27004 6560 27324 7584
rect 27004 6496 27012 6560
rect 27076 6496 27092 6560
rect 27156 6496 27172 6560
rect 27236 6496 27252 6560
rect 27316 6496 27324 6560
rect 27004 5472 27324 6496
rect 27004 5408 27012 5472
rect 27076 5408 27092 5472
rect 27156 5408 27172 5472
rect 27236 5408 27252 5472
rect 27316 5408 27324 5472
rect 27004 4384 27324 5408
rect 27004 4320 27012 4384
rect 27076 4320 27092 4384
rect 27156 4320 27172 4384
rect 27236 4320 27252 4384
rect 27316 4320 27324 4384
rect 27004 3296 27324 4320
rect 27004 3232 27012 3296
rect 27076 3232 27092 3296
rect 27156 3232 27172 3296
rect 27236 3232 27252 3296
rect 27316 3232 27324 3296
rect 27004 2208 27324 3232
rect 27004 2144 27012 2208
rect 27076 2144 27092 2208
rect 27156 2144 27172 2208
rect 27236 2144 27252 2208
rect 27316 2144 27324 2208
rect 27004 0 27324 2144
rect 31944 8192 32264 11250
rect 31944 8128 31952 8192
rect 32016 8128 32032 8192
rect 32096 8128 32112 8192
rect 32176 8128 32192 8192
rect 32256 8128 32264 8192
rect 31944 7104 32264 8128
rect 31944 7040 31952 7104
rect 32016 7040 32032 7104
rect 32096 7040 32112 7104
rect 32176 7040 32192 7104
rect 32256 7040 32264 7104
rect 31944 6016 32264 7040
rect 31944 5952 31952 6016
rect 32016 5952 32032 6016
rect 32096 5952 32112 6016
rect 32176 5952 32192 6016
rect 32256 5952 32264 6016
rect 31944 4928 32264 5952
rect 31944 4864 31952 4928
rect 32016 4864 32032 4928
rect 32096 4864 32112 4928
rect 32176 4864 32192 4928
rect 32256 4864 32264 4928
rect 31944 3840 32264 4864
rect 31944 3776 31952 3840
rect 32016 3776 32032 3840
rect 32096 3776 32112 3840
rect 32176 3776 32192 3840
rect 32256 3776 32264 3840
rect 31944 2752 32264 3776
rect 31944 2688 31952 2752
rect 32016 2688 32032 2752
rect 32096 2688 32112 2752
rect 32176 2688 32192 2752
rect 32256 2688 32264 2752
rect 31944 0 32264 2688
use sky130_fd_sc_hd__buf_1  _00_
timestamp -3599
transform 1 0 17572 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _01_
timestamp -3599
transform 1 0 20608 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _02_
timestamp -3599
transform -1 0 21988 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _03_
timestamp -3599
transform -1 0 21712 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _04_
timestamp -3599
transform 1 0 19688 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _05_
timestamp -3599
transform -1 0 26680 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _06_
timestamp -3599
transform -1 0 26220 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _07_
timestamp -3599
transform -1 0 25668 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _08_
timestamp -3599
transform -1 0 25576 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _09_
timestamp -3599
transform 1 0 18216 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _10_
timestamp -3599
transform -1 0 23552 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _11_
timestamp -3599
transform 1 0 21160 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _12_
timestamp -3599
transform 1 0 19504 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _13_
timestamp -3599
transform 1 0 17204 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _14_
timestamp -3599
transform 1 0 11868 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _15_
timestamp -3599
transform 1 0 12880 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _16_
timestamp -3599
transform 1 0 14996 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _17_
timestamp -3599
transform 1 0 17940 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _18_
timestamp -3599
transform 1 0 9292 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _19_
timestamp -3599
transform 1 0 13708 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _20_
timestamp -3599
transform -1 0 9016 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _21_
timestamp -3599
transform 1 0 6532 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _22_
timestamp -3599
transform 1 0 16652 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _23_
timestamp -3599
transform 1 0 6808 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _24_
timestamp -3599
transform 1 0 14720 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _25_
timestamp -3599
transform 1 0 13984 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _26_
timestamp -3599
transform 1 0 16192 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _27_
timestamp -3599
transform 1 0 12144 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _28_
timestamp -3599
transform 1 0 12420 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _29_
timestamp -3599
transform 1 0 5704 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _30_
timestamp -3599
transform -1 0 9292 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _31_
timestamp -3599
transform 1 0 17296 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _32_
timestamp -3599
transform -1 0 24472 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _33_
timestamp -3599
transform -1 0 20976 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _34_
timestamp -3599
transform -1 0 20516 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _35_
timestamp -3599
transform 1 0 14260 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _36_
timestamp -3599
transform -1 0 19964 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _37_
timestamp -3599
transform -1 0 23184 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _38_
timestamp -3599
transform -1 0 25576 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _39_
timestamp -3599
transform -1 0 25392 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _40_
timestamp -3599
transform 1 0 23644 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _41_
timestamp -3599
transform 1 0 21896 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _42_
timestamp -3599
transform 1 0 20424 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _43_
timestamp -3599
transform 1 0 20976 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _44_
timestamp -3599
transform 1 0 22172 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _45_
timestamp -3599
transform 1 0 23092 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _46_
timestamp -3599
transform -1 0 23736 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _47_
timestamp -3599
transform -1 0 24104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _48_
timestamp -3599
transform -1 0 25116 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _49_
timestamp -3599
transform -1 0 27232 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _50_
timestamp -3599
transform -1 0 29256 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _51_
timestamp -3599
transform -1 0 30912 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _52_
timestamp -3599
transform -1 0 10856 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _53_
timestamp -3599
transform -1 0 8280 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _54_
timestamp -3599
transform -1 0 7452 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _55_
timestamp -3599
transform 1 0 5428 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _56_
timestamp -3599
transform -1 0 13064 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _57_
timestamp -3599
transform -1 0 12604 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _58_
timestamp -3599
transform -1 0 11776 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _59_
timestamp -3599
transform -1 0 9200 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _60_
timestamp -3599
transform 1 0 7452 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _61_
timestamp -3599
transform 1 0 5704 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _62_
timestamp -3599
transform 1 0 3772 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _63_
timestamp -3599
transform 1 0 2576 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _64_
timestamp -3599
transform -1 0 14076 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _65_
timestamp -3599
transform -1 0 13800 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _66_
timestamp -3599
transform -1 0 11224 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _67_
timestamp -3599
transform 1 0 9752 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _68_
timestamp -3599
transform 1 0 8372 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _69_
timestamp -3599
transform 1 0 7176 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _70_
timestamp -3599
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _71_
timestamp -3599
transform 1 0 4692 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _72_
timestamp -3599
transform -1 0 12696 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _73_
timestamp -3599
transform -1 0 12420 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _74_
timestamp -3599
transform -1 0 12696 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _75_
timestamp -3599
transform -1 0 12972 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _76_
timestamp -3599
transform -1 0 13340 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _77_
timestamp -3599
transform -1 0 14720 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _78_
timestamp -3599
transform -1 0 14444 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _79_
timestamp -3599
transform -1 0 14444 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _80_
timestamp -3599
transform -1 0 15364 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _81_
timestamp -3599
transform -1 0 16008 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _82_
timestamp -3599
transform -1 0 16928 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _83_
timestamp -3599
transform -1 0 17388 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _84_
timestamp -3599
transform -1 0 18308 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _85_
timestamp -3599
transform -1 0 19688 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _86_
timestamp -3599
transform -1 0 20056 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _87_
timestamp -3599
transform -1 0 20332 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _88_
timestamp -3599
transform 1 0 24932 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp -3599
transform 1 0 17388 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp -3599
transform 1 0 23092 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp -3599
transform 1 0 20976 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp -3599
transform -1 0 19504 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp -3599
transform -1 0 17204 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp -3599
transform 1 0 12696 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp -3599
transform -1 0 15456 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp -3599
transform 1 0 17756 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp -3599
transform 1 0 13524 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp -3599
transform -1 0 20608 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp -3599
transform -1 0 17112 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp -3599
transform -1 0 14720 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp -3599
transform -1 0 13524 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp -3599
transform -1 0 16192 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp -3599
transform -1 0 22172 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp -3599
transform -1 0 17296 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp -3599
transform -1 0 21436 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp -3599
transform 1 0 18952 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp -3599
transform -1 0 26404 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp -3599
transform -1 0 25944 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp -3599
transform -1 0 25392 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_22
timestamp -3599
transform -1 0 25300 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_23
timestamp -3599
transform -1 0 18216 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_24
timestamp -3599
transform -1 0 13340 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_25
timestamp -3599
transform 1 0 19228 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3
timestamp 1636964856
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1636964856
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27
timestamp -3599
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1636964856
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1636964856
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53
timestamp -3599
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1636964856
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1636964856
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp -3599
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1636964856
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1636964856
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp -3599
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1636964856
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_125
timestamp -3599
transform 1 0 12604 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_133
timestamp -3599
transform 1 0 13340 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_141
timestamp -3599
transform 1 0 14076 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_169
timestamp -3599
transform 1 0 16652 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_182
timestamp -3599
transform 1 0 17848 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp -3599
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp -3599
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_257
timestamp 1636964856
transform 1 0 24748 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_269
timestamp -3599
transform 1 0 25852 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp -3599
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_281
timestamp 1636964856
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_293
timestamp 1636964856
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp -3599
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_309
timestamp -3599
transform 1 0 29532 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_317
timestamp -3599
transform 1 0 30268 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_337
timestamp -3599
transform 1 0 32108 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1636964856
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1636964856
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1636964856
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1636964856
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp -3599
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp -3599
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1636964856
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1636964856
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1636964856
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1636964856
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp -3599
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp -3599
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1636964856
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1636964856
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_137
timestamp -3599
transform 1 0 13708 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_149
timestamp -3599
transform 1 0 14812 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_153
timestamp -3599
transform 1 0 15180 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_158
timestamp -3599
transform 1 0 15640 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_162
timestamp -3599
transform 1 0 16008 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp -3599
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1636964856
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1636964856
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_193
timestamp -3599
transform 1 0 18860 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_203
timestamp -3599
transform 1 0 19780 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_219
timestamp -3599
transform 1 0 21252 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp -3599
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_229
timestamp -3599
transform 1 0 22172 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_239
timestamp -3599
transform 1 0 23092 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_245
timestamp -3599
transform 1 0 23644 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_251
timestamp 1636964856
transform 1 0 24196 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_263
timestamp 1636964856
transform 1 0 25300 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_275
timestamp -3599
transform 1 0 26404 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp -3599
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1636964856
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_293
timestamp 1636964856
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_305
timestamp 1636964856
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_317
timestamp -3599
transform 1 0 30268 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_325
timestamp -3599
transform 1 0 31004 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_337
timestamp -3599
transform 1 0 32108 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1636964856
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1636964856
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp -3599
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1636964856
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1636964856
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1636964856
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1636964856
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp -3599
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp -3599
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1636964856
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1636964856
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1636964856
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_121
timestamp -3599
transform 1 0 12236 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_126
timestamp 1636964856
transform 1 0 12696 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp -3599
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1636964856
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1636964856
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1636964856
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1636964856
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp -3599
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp -3599
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_197
timestamp -3599
transform 1 0 19228 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_209
timestamp -3599
transform 1 0 20332 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_215
timestamp -3599
transform 1 0 20884 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_229
timestamp 1636964856
transform 1 0 22172 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_241
timestamp -3599
transform 1 0 23276 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_249
timestamp -3599
transform 1 0 24012 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_253
timestamp -3599
transform 1 0 24380 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_261
timestamp -3599
transform 1 0 25116 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_267
timestamp -3599
transform 1 0 25668 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_278
timestamp 1636964856
transform 1 0 26680 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_290
timestamp 1636964856
transform 1 0 27784 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_302
timestamp -3599
transform 1 0 28888 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1636964856
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_321
timestamp -3599
transform 1 0 30636 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_329
timestamp -3599
transform 1 0 31372 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1636964856
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1636964856
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1636964856
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1636964856
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp -3599
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp -3599
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1636964856
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1636964856
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1636964856
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1636964856
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp -3599
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp -3599
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_113
timestamp -3599
transform 1 0 11500 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_119
timestamp -3599
transform 1 0 12052 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_129
timestamp -3599
transform 1 0 12972 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_133
timestamp -3599
transform 1 0 13340 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_141
timestamp -3599
transform 1 0 14076 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_148
timestamp -3599
transform 1 0 14720 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_155
timestamp -3599
transform 1 0 15364 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_162
timestamp -3599
transform 1 0 16008 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_3_172
timestamp -3599
transform 1 0 16928 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_182
timestamp -3599
transform 1 0 17848 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_187
timestamp -3599
transform 1 0 18308 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_193
timestamp -3599
transform 1 0 18860 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_196
timestamp -3599
transform 1 0 19136 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1636964856
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp -3599
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp -3599
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_225
timestamp -3599
transform 1 0 21804 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_232
timestamp -3599
transform 1 0 22448 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_238
timestamp -3599
transform 1 0 23000 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_242
timestamp -3599
transform 1 0 23368 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_246
timestamp -3599
transform 1 0 23736 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_250
timestamp 1636964856
transform 1 0 24104 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_262
timestamp 1636964856
transform 1 0 25208 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_274
timestamp -3599
transform 1 0 26312 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1636964856
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1636964856
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1636964856
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_317
timestamp -3599
transform 1 0 30268 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_325
timestamp -3599
transform 1 0 31004 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_337
timestamp -3599
transform 1 0 32108 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1636964856
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_15
timestamp -3599
transform 1 0 2484 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_19
timestamp -3599
transform 1 0 2852 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp -3599
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1636964856
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1636964856
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1636964856
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1636964856
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp -3599
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp -3599
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1636964856
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1636964856
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_109
timestamp -3599
transform 1 0 11132 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_116
timestamp -3599
transform 1 0 11776 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_125
timestamp -3599
transform 1 0 12604 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_130
timestamp -3599
transform 1 0 13064 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_138
timestamp -3599
transform 1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_141
timestamp -3599
transform 1 0 14076 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_145
timestamp 1636964856
transform 1 0 14444 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_157
timestamp 1636964856
transform 1 0 15548 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_169
timestamp 1636964856
transform 1 0 16652 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_181
timestamp 1636964856
transform 1 0 17756 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_193
timestamp -3599
transform 1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1636964856
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1636964856
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1636964856
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1636964856
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp -3599
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp -3599
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_253
timestamp -3599
transform 1 0 24380 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_257
timestamp -3599
transform 1 0 24748 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_266
timestamp 1636964856
transform 1 0 25576 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_278
timestamp 1636964856
transform 1 0 26680 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_290
timestamp 1636964856
transform 1 0 27784 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_302
timestamp -3599
transform 1 0 28888 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1636964856
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_321
timestamp -3599
transform 1 0 30636 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_329
timestamp -3599
transform 1 0 31372 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1636964856
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1636964856
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1636964856
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_39
timestamp -3599
transform 1 0 4692 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_5_50
timestamp -3599
transform 1 0 5704 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1636964856
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1636964856
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1636964856
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_93
timestamp -3599
transform 1 0 9660 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_101
timestamp -3599
transform 1 0 10396 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_106
timestamp -3599
transform 1 0 10856 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1636964856
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1636964856
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1636964856
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1636964856
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp -3599
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp -3599
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1636964856
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1636964856
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1636964856
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1636964856
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp -3599
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp -3599
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1636964856
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_237
timestamp -3599
transform 1 0 22908 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_244
timestamp -3599
transform 1 0 23552 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_248
timestamp 1636964856
transform 1 0 23920 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_260
timestamp 1636964856
transform 1 0 25024 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_272
timestamp -3599
transform 1 0 26128 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_5_284
timestamp 1636964856
transform 1 0 27232 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_296
timestamp 1636964856
transform 1 0 28336 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_308
timestamp 1636964856
transform 1 0 29440 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_320
timestamp -3599
transform 1 0 30544 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_337
timestamp -3599
transform 1 0 32108 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1636964856
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1636964856
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp -3599
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_32
timestamp 1636964856
transform 1 0 4048 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_44
timestamp 1636964856
transform 1 0 5152 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_56
timestamp 1636964856
transform 1 0 6256 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_68
timestamp 1636964856
transform 1 0 7360 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_80
timestamp -3599
transform 1 0 8464 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1636964856
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_97
timestamp -3599
transform 1 0 10028 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_105
timestamp -3599
transform 1 0 10764 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_110
timestamp 1636964856
transform 1 0 11224 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_122
timestamp 1636964856
transform 1 0 12328 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_134
timestamp -3599
transform 1 0 13432 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1636964856
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1636964856
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1636964856
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_177
timestamp -3599
transform 1 0 17388 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_183
timestamp -3599
transform 1 0 17940 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp -3599
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp -3599
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1636964856
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_209
timestamp -3599
transform 1 0 20332 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_215
timestamp -3599
transform 1 0 20884 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_219
timestamp -3599
transform 1 0 21252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_225
timestamp -3599
transform 1 0 21804 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_229
timestamp 1636964856
transform 1 0 22172 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_241
timestamp -3599
transform 1 0 23276 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_249
timestamp -3599
transform 1 0 24012 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1636964856
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1636964856
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1636964856
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1636964856
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_301
timestamp -3599
transform 1 0 28796 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_306
timestamp -3599
transform 1 0 29256 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1636964856
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_324
timestamp -3599
transform 1 0 30912 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1636964856
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1636964856
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1636964856
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1636964856
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp -3599
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp -3599
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_57
timestamp -3599
transform 1 0 6348 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_65
timestamp -3599
transform 1 0 7084 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1636964856
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1636964856
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_93
timestamp -3599
transform 1 0 9660 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_97
timestamp 1636964856
transform 1 0 10028 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_109
timestamp -3599
transform 1 0 11132 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1636964856
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1636964856
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1636964856
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1636964856
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp -3599
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp -3599
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1636964856
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1636964856
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1636964856
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_205
timestamp -3599
transform 1 0 19964 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_209
timestamp -3599
transform 1 0 20332 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_213
timestamp -3599
transform 1 0 20700 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_221
timestamp -3599
transform 1 0 21436 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1636964856
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1636964856
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1636964856
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1636964856
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp -3599
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp -3599
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1636964856
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1636964856
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1636964856
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_317
timestamp -3599
transform 1 0 30268 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_325
timestamp -3599
transform 1 0 31004 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_337
timestamp -3599
transform 1 0 32108 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1636964856
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1636964856
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp -3599
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1636964856
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_41
timestamp -3599
transform 1 0 4876 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_49
timestamp -3599
transform 1 0 5612 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1636964856
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_65
timestamp -3599
transform 1 0 7084 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_73
timestamp -3599
transform 1 0 7820 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_78
timestamp -3599
transform 1 0 8280 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_82
timestamp -3599
transform 1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_88
timestamp 1636964856
transform 1 0 9200 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_100
timestamp 1636964856
transform 1 0 10304 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_112
timestamp 1636964856
transform 1 0 11408 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_124
timestamp 1636964856
transform 1 0 12512 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_136
timestamp -3599
transform 1 0 13616 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1636964856
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1636964856
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_165
timestamp -3599
transform 1 0 16284 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_8_178
timestamp 1636964856
transform 1 0 17480 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_190
timestamp -3599
transform 1 0 18584 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_197
timestamp -3599
transform 1 0 19228 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_203
timestamp 1636964856
transform 1 0 19780 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_215
timestamp 1636964856
transform 1 0 20884 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_227
timestamp 1636964856
transform 1 0 21988 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_239
timestamp 1636964856
transform 1 0 23092 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp -3599
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_253
timestamp -3599
transform 1 0 24380 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_8_264
timestamp 1636964856
transform 1 0 25392 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_276
timestamp 1636964856
transform 1 0 26496 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_288
timestamp 1636964856
transform 1 0 27600 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_300
timestamp -3599
transform 1 0 28704 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1636964856
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_321
timestamp -3599
transform 1 0 30636 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1636964856
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1636964856
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1636964856
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_42
timestamp -3599
transform 1 0 4968 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_57
timestamp -3599
transform 1 0 6348 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_65
timestamp -3599
transform 1 0 7084 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_72
timestamp -3599
transform 1 0 7728 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_80
timestamp -3599
transform 1 0 8464 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_92
timestamp 1636964856
transform 1 0 9568 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_104
timestamp -3599
transform 1 0 10672 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_113
timestamp -3599
transform 1 0 11500 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_156
timestamp -3599
transform 1 0 15456 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp -3599
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_179
timestamp -3599
transform 1 0 17572 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_186
timestamp 1636964856
transform 1 0 18216 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_198
timestamp -3599
transform 1 0 19320 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_9_205
timestamp -3599
transform 1 0 19964 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_211
timestamp -3599
transform 1 0 20516 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_216
timestamp -3599
transform 1 0 20976 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1636964856
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_240
timestamp -3599
transform 1 0 23184 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_248
timestamp -3599
transform 1 0 23920 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_254
timestamp -3599
transform 1 0 24472 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_258
timestamp -3599
transform 1 0 24840 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_266
timestamp 1636964856
transform 1 0 25576 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_278
timestamp -3599
transform 1 0 26680 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1636964856
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1636964856
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1636964856
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_317
timestamp -3599
transform 1 0 30268 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_325
timestamp -3599
transform 1 0 31004 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_337
timestamp -3599
transform 1 0 32108 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1636964856
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1636964856
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp -3599
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1636964856
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1636964856
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1636964856
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1636964856
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp -3599
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp -3599
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1636964856
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1636964856
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1636964856
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1636964856
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp -3599
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp -3599
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1636964856
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1636964856
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1636964856
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1636964856
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp -3599
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp -3599
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1636964856
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1636964856
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1636964856
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_233
timestamp 1636964856
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp -3599
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp -3599
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1636964856
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1636964856
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1636964856
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_289
timestamp 1636964856
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp -3599
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp -3599
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_309
timestamp -3599
transform 1 0 29532 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_317
timestamp -3599
transform 1 0 30268 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_6
timestamp 1636964856
transform 1 0 1656 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_18
timestamp -3599
transform 1 0 2760 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_23
timestamp -3599
transform 1 0 3220 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_27
timestamp -3599
transform 1 0 3588 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_29
timestamp -3599
transform 1 0 3772 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_35
timestamp -3599
transform 1 0 4324 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_40
timestamp 1636964856
transform 1 0 4784 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_52
timestamp -3599
transform 1 0 5888 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_61
timestamp -3599
transform 1 0 6716 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_69
timestamp -3599
transform 1 0 7452 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_74
timestamp -3599
transform 1 0 7912 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_82
timestamp -3599
transform 1 0 8648 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_85
timestamp -3599
transform 1 0 8924 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_91
timestamp 1636964856
transform 1 0 9476 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_103
timestamp -3599
transform 1 0 10580 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_108
timestamp -3599
transform 1 0 11040 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_113
timestamp -3599
transform 1 0 11500 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1636964856
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_137
timestamp -3599
transform 1 0 13708 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_145
timestamp -3599
transform 1 0 14444 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_153
timestamp -3599
transform 1 0 15180 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_159
timestamp -3599
transform 1 0 15732 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp -3599
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_169
timestamp -3599
transform 1 0 16652 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_176
timestamp 1636964856
transform 1 0 17296 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_188
timestamp -3599
transform 1 0 18400 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_193
timestamp -3599
transform 1 0 18860 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_197
timestamp -3599
transform 1 0 19228 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_205
timestamp -3599
transform 1 0 19964 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_210
timestamp 1636964856
transform 1 0 20424 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_222
timestamp -3599
transform 1 0 21528 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_229
timestamp -3599
transform 1 0 22172 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_237
timestamp -3599
transform 1 0 22908 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_244
timestamp -3599
transform 1 0 23552 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_253
timestamp -3599
transform 1 0 24380 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_261
timestamp 1636964856
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_273
timestamp -3599
transform 1 0 26220 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_278
timestamp -3599
transform 1 0 26680 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_281
timestamp -3599
transform 1 0 26956 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_289
timestamp -3599
transform 1 0 27692 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_295
timestamp 1636964856
transform 1 0 28244 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_307
timestamp -3599
transform 1 0 29348 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_329
timestamp -3599
transform 1 0 31372 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_337
timestamp -3599
transform 1 0 32108 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  output1
timestamp -3599
transform 1 0 31280 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output2
timestamp -3599
transform 1 0 31556 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output3
timestamp -3599
transform 1 0 31924 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output4
timestamp -3599
transform 1 0 31280 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output5
timestamp -3599
transform 1 0 31648 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output6
timestamp -3599
transform 1 0 31188 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output7
timestamp -3599
transform 1 0 31556 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output8
timestamp -3599
transform 1 0 31924 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output9
timestamp -3599
transform 1 0 31280 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp -3599
transform 1 0 31648 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp -3599
transform 1 0 31188 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp -3599
transform 1 0 30912 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp -3599
transform 1 0 31556 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp -3599
transform 1 0 31648 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output15
timestamp -3599
transform 1 0 31556 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output16
timestamp -3599
transform 1 0 31924 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output17
timestamp -3599
transform 1 0 31648 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output18
timestamp -3599
transform 1 0 30636 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output19
timestamp -3599
transform 1 0 31188 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output20
timestamp -3599
transform 1 0 30820 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output21
timestamp -3599
transform 1 0 30268 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output22
timestamp -3599
transform 1 0 31280 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output23
timestamp -3599
transform 1 0 30544 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output24
timestamp -3599
transform 1 0 30452 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output25
timestamp -3599
transform 1 0 29900 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output26
timestamp -3599
transform 1 0 31648 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output27
timestamp -3599
transform 1 0 31280 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output28
timestamp -3599
transform 1 0 31648 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output29
timestamp -3599
transform 1 0 31556 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output30
timestamp -3599
transform 1 0 31924 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output31
timestamp -3599
transform 1 0 31280 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output32
timestamp -3599
transform 1 0 31648 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output33
timestamp -3599
transform -1 0 3220 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output34
timestamp -3599
transform -1 0 18860 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output35
timestamp -3599
transform -1 0 20424 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output36
timestamp -3599
transform -1 0 22172 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output37
timestamp -3599
transform 1 0 23184 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output38
timestamp -3599
transform 1 0 24748 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output39
timestamp -3599
transform 1 0 26312 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output40
timestamp -3599
transform 1 0 27876 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output41
timestamp -3599
transform 1 0 29532 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output42
timestamp -3599
transform 1 0 31004 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output43
timestamp -3599
transform 1 0 31924 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output44
timestamp -3599
transform -1 0 4784 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output45
timestamp -3599
transform -1 0 6716 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output46
timestamp -3599
transform -1 0 7912 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output47
timestamp -3599
transform -1 0 9476 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output48
timestamp -3599
transform -1 0 11040 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output49
timestamp -3599
transform -1 0 12604 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output50
timestamp -3599
transform -1 0 14444 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output51
timestamp -3599
transform -1 0 15732 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output52
timestamp -3599
transform -1 0 17296 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output53
timestamp -3599
transform 1 0 13616 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output54
timestamp -3599
transform 1 0 14444 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output55
timestamp -3599
transform 1 0 14352 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output56
timestamp -3599
transform 1 0 14720 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output57
timestamp -3599
transform 1 0 15272 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output58
timestamp -3599
transform 1 0 15088 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output59
timestamp -3599
transform 1 0 15456 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output60
timestamp -3599
transform 1 0 16100 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output61
timestamp -3599
transform 1 0 15824 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp -3599
transform 1 0 16192 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output63
timestamp -3599
transform 1 0 16744 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp -3599
transform 1 0 17112 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp -3599
transform 1 0 17480 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp -3599
transform 1 0 18400 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp -3599
transform 1 0 18032 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp -3599
transform 1 0 18768 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp -3599
transform 1 0 19228 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp -3599
transform 1 0 19596 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp -3599
transform 1 0 19964 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp -3599
transform 1 0 19412 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp -3599
transform 1 0 20332 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp -3599
transform 1 0 23276 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp -3599
transform 1 0 22724 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp -3599
transform 1 0 23644 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp -3599
transform 1 0 23276 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp -3599
transform 1 0 24380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp -3599
transform 1 0 23828 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp -3599
transform 1 0 20700 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp -3599
transform 1 0 21068 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp -3599
transform 1 0 20516 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp -3599
transform 1 0 20884 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp -3599
transform 1 0 21804 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp -3599
transform 1 0 22172 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp -3599
transform 1 0 21804 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp -3599
transform 1 0 22540 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp -3599
transform 1 0 22908 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  output89
timestamp -3599
transform -1 0 1656 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_12
timestamp -3599
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp -3599
transform -1 0 32568 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_13
timestamp -3599
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp -3599
transform -1 0 32568 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_14
timestamp -3599
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp -3599
transform -1 0 32568 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_15
timestamp -3599
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp -3599
transform -1 0 32568 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_16
timestamp -3599
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp -3599
transform -1 0 32568 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_17
timestamp -3599
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp -3599
transform -1 0 32568 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_18
timestamp -3599
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp -3599
transform -1 0 32568 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_19
timestamp -3599
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp -3599
transform -1 0 32568 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_20
timestamp -3599
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp -3599
transform -1 0 32568 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_21
timestamp -3599
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp -3599
transform -1 0 32568 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_22
timestamp -3599
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp -3599
transform -1 0 32568 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_23
timestamp -3599
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp -3599
transform -1 0 32568 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_24
timestamp -3599
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_25
timestamp -3599
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_26
timestamp -3599
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_27
timestamp -3599
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_28
timestamp -3599
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_29
timestamp -3599
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_30
timestamp -3599
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_31
timestamp -3599
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_32
timestamp -3599
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_33
timestamp -3599
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_34
timestamp -3599
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_35
timestamp -3599
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_36
timestamp -3599
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_37
timestamp -3599
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_38
timestamp -3599
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_39
timestamp -3599
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_40
timestamp -3599
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_41
timestamp -3599
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_42
timestamp -3599
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_43
timestamp -3599
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_44
timestamp -3599
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_45
timestamp -3599
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_46
timestamp -3599
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_47
timestamp -3599
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_48
timestamp -3599
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_49
timestamp -3599
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_50
timestamp -3599
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_51
timestamp -3599
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_52
timestamp -3599
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_53
timestamp -3599
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_54
timestamp -3599
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_55
timestamp -3599
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_56
timestamp -3599
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_57
timestamp -3599
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_58
timestamp -3599
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_59
timestamp -3599
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_60
timestamp -3599
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_61
timestamp -3599
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_62
timestamp -3599
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_63
timestamp -3599
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_64
timestamp -3599
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_65
timestamp -3599
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_66
timestamp -3599
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_67
timestamp -3599
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_68
timestamp -3599
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_69
timestamp -3599
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_70
timestamp -3599
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_71
timestamp -3599
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_72
timestamp -3599
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_73
timestamp -3599
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_74
timestamp -3599
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_75
timestamp -3599
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_76
timestamp -3599
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_77
timestamp -3599
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_78
timestamp -3599
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_79
timestamp -3599
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_80
timestamp -3599
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_81
timestamp -3599
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_82
timestamp -3599
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_83
timestamp -3599
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_84
timestamp -3599
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_85
timestamp -3599
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_86
timestamp -3599
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_87
timestamp -3599
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_88
timestamp -3599
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_89
timestamp -3599
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_90
timestamp -3599
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_91
timestamp -3599
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_92
timestamp -3599
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_93
timestamp -3599
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_94
timestamp -3599
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_95
timestamp -3599
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_96
timestamp -3599
transform 1 0 3680 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_97
timestamp -3599
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_98
timestamp -3599
transform 1 0 8832 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_99
timestamp -3599
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_100
timestamp -3599
transform 1 0 13984 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_101
timestamp -3599
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_102
timestamp -3599
transform 1 0 19136 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_103
timestamp -3599
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_104
timestamp -3599
transform 1 0 24288 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_105
timestamp -3599
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_106
timestamp -3599
transform 1 0 29440 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_107
timestamp -3599
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
<< labels >>
flabel metal3 s 0 1368 120 1488 0 FreeSans 480 0 0 0 FrameData[0]
port 0 nsew signal input
flabel metal3 s 0 4088 120 4208 0 FreeSans 480 0 0 0 FrameData[10]
port 1 nsew signal input
flabel metal3 s 0 4360 120 4480 0 FreeSans 480 0 0 0 FrameData[11]
port 2 nsew signal input
flabel metal3 s 0 4632 120 4752 0 FreeSans 480 0 0 0 FrameData[12]
port 3 nsew signal input
flabel metal3 s 0 4904 120 5024 0 FreeSans 480 0 0 0 FrameData[13]
port 4 nsew signal input
flabel metal3 s 0 5176 120 5296 0 FreeSans 480 0 0 0 FrameData[14]
port 5 nsew signal input
flabel metal3 s 0 5448 120 5568 0 FreeSans 480 0 0 0 FrameData[15]
port 6 nsew signal input
flabel metal3 s 0 5720 120 5840 0 FreeSans 480 0 0 0 FrameData[16]
port 7 nsew signal input
flabel metal3 s 0 5992 120 6112 0 FreeSans 480 0 0 0 FrameData[17]
port 8 nsew signal input
flabel metal3 s 0 6264 120 6384 0 FreeSans 480 0 0 0 FrameData[18]
port 9 nsew signal input
flabel metal3 s 0 6536 120 6656 0 FreeSans 480 0 0 0 FrameData[19]
port 10 nsew signal input
flabel metal3 s 0 1640 120 1760 0 FreeSans 480 0 0 0 FrameData[1]
port 11 nsew signal input
flabel metal3 s 0 6808 120 6928 0 FreeSans 480 0 0 0 FrameData[20]
port 12 nsew signal input
flabel metal3 s 0 7080 120 7200 0 FreeSans 480 0 0 0 FrameData[21]
port 13 nsew signal input
flabel metal3 s 0 7352 120 7472 0 FreeSans 480 0 0 0 FrameData[22]
port 14 nsew signal input
flabel metal3 s 0 7624 120 7744 0 FreeSans 480 0 0 0 FrameData[23]
port 15 nsew signal input
flabel metal3 s 0 7896 120 8016 0 FreeSans 480 0 0 0 FrameData[24]
port 16 nsew signal input
flabel metal3 s 0 8168 120 8288 0 FreeSans 480 0 0 0 FrameData[25]
port 17 nsew signal input
flabel metal3 s 0 8440 120 8560 0 FreeSans 480 0 0 0 FrameData[26]
port 18 nsew signal input
flabel metal3 s 0 8712 120 8832 0 FreeSans 480 0 0 0 FrameData[27]
port 19 nsew signal input
flabel metal3 s 0 8984 120 9104 0 FreeSans 480 0 0 0 FrameData[28]
port 20 nsew signal input
flabel metal3 s 0 9256 120 9376 0 FreeSans 480 0 0 0 FrameData[29]
port 21 nsew signal input
flabel metal3 s 0 1912 120 2032 0 FreeSans 480 0 0 0 FrameData[2]
port 22 nsew signal input
flabel metal3 s 0 9528 120 9648 0 FreeSans 480 0 0 0 FrameData[30]
port 23 nsew signal input
flabel metal3 s 0 9800 120 9920 0 FreeSans 480 0 0 0 FrameData[31]
port 24 nsew signal input
flabel metal3 s 0 2184 120 2304 0 FreeSans 480 0 0 0 FrameData[3]
port 25 nsew signal input
flabel metal3 s 0 2456 120 2576 0 FreeSans 480 0 0 0 FrameData[4]
port 26 nsew signal input
flabel metal3 s 0 2728 120 2848 0 FreeSans 480 0 0 0 FrameData[5]
port 27 nsew signal input
flabel metal3 s 0 3000 120 3120 0 FreeSans 480 0 0 0 FrameData[6]
port 28 nsew signal input
flabel metal3 s 0 3272 120 3392 0 FreeSans 480 0 0 0 FrameData[7]
port 29 nsew signal input
flabel metal3 s 0 3544 120 3664 0 FreeSans 480 0 0 0 FrameData[8]
port 30 nsew signal input
flabel metal3 s 0 3816 120 3936 0 FreeSans 480 0 0 0 FrameData[9]
port 31 nsew signal input
flabel metal3 s 33630 1368 33750 1488 0 FreeSans 480 0 0 0 FrameData_O[0]
port 32 nsew signal output
flabel metal3 s 33630 4088 33750 4208 0 FreeSans 480 0 0 0 FrameData_O[10]
port 33 nsew signal output
flabel metal3 s 33630 4360 33750 4480 0 FreeSans 480 0 0 0 FrameData_O[11]
port 34 nsew signal output
flabel metal3 s 33630 4632 33750 4752 0 FreeSans 480 0 0 0 FrameData_O[12]
port 35 nsew signal output
flabel metal3 s 33630 4904 33750 5024 0 FreeSans 480 0 0 0 FrameData_O[13]
port 36 nsew signal output
flabel metal3 s 33630 5176 33750 5296 0 FreeSans 480 0 0 0 FrameData_O[14]
port 37 nsew signal output
flabel metal3 s 33630 5448 33750 5568 0 FreeSans 480 0 0 0 FrameData_O[15]
port 38 nsew signal output
flabel metal3 s 33630 5720 33750 5840 0 FreeSans 480 0 0 0 FrameData_O[16]
port 39 nsew signal output
flabel metal3 s 33630 5992 33750 6112 0 FreeSans 480 0 0 0 FrameData_O[17]
port 40 nsew signal output
flabel metal3 s 33630 6264 33750 6384 0 FreeSans 480 0 0 0 FrameData_O[18]
port 41 nsew signal output
flabel metal3 s 33630 6536 33750 6656 0 FreeSans 480 0 0 0 FrameData_O[19]
port 42 nsew signal output
flabel metal3 s 33630 1640 33750 1760 0 FreeSans 480 0 0 0 FrameData_O[1]
port 43 nsew signal output
flabel metal3 s 33630 6808 33750 6928 0 FreeSans 480 0 0 0 FrameData_O[20]
port 44 nsew signal output
flabel metal3 s 33630 7080 33750 7200 0 FreeSans 480 0 0 0 FrameData_O[21]
port 45 nsew signal output
flabel metal3 s 33630 7352 33750 7472 0 FreeSans 480 0 0 0 FrameData_O[22]
port 46 nsew signal output
flabel metal3 s 33630 7624 33750 7744 0 FreeSans 480 0 0 0 FrameData_O[23]
port 47 nsew signal output
flabel metal3 s 33630 7896 33750 8016 0 FreeSans 480 0 0 0 FrameData_O[24]
port 48 nsew signal output
flabel metal3 s 33630 8168 33750 8288 0 FreeSans 480 0 0 0 FrameData_O[25]
port 49 nsew signal output
flabel metal3 s 33630 8440 33750 8560 0 FreeSans 480 0 0 0 FrameData_O[26]
port 50 nsew signal output
flabel metal3 s 33630 8712 33750 8832 0 FreeSans 480 0 0 0 FrameData_O[27]
port 51 nsew signal output
flabel metal3 s 33630 8984 33750 9104 0 FreeSans 480 0 0 0 FrameData_O[28]
port 52 nsew signal output
flabel metal3 s 33630 9256 33750 9376 0 FreeSans 480 0 0 0 FrameData_O[29]
port 53 nsew signal output
flabel metal3 s 33630 1912 33750 2032 0 FreeSans 480 0 0 0 FrameData_O[2]
port 54 nsew signal output
flabel metal3 s 33630 9528 33750 9648 0 FreeSans 480 0 0 0 FrameData_O[30]
port 55 nsew signal output
flabel metal3 s 33630 9800 33750 9920 0 FreeSans 480 0 0 0 FrameData_O[31]
port 56 nsew signal output
flabel metal3 s 33630 2184 33750 2304 0 FreeSans 480 0 0 0 FrameData_O[3]
port 57 nsew signal output
flabel metal3 s 33630 2456 33750 2576 0 FreeSans 480 0 0 0 FrameData_O[4]
port 58 nsew signal output
flabel metal3 s 33630 2728 33750 2848 0 FreeSans 480 0 0 0 FrameData_O[5]
port 59 nsew signal output
flabel metal3 s 33630 3000 33750 3120 0 FreeSans 480 0 0 0 FrameData_O[6]
port 60 nsew signal output
flabel metal3 s 33630 3272 33750 3392 0 FreeSans 480 0 0 0 FrameData_O[7]
port 61 nsew signal output
flabel metal3 s 33630 3544 33750 3664 0 FreeSans 480 0 0 0 FrameData_O[8]
port 62 nsew signal output
flabel metal3 s 33630 3816 33750 3936 0 FreeSans 480 0 0 0 FrameData_O[9]
port 63 nsew signal output
flabel metal2 s 24306 0 24362 56 0 FreeSans 224 0 0 0 FrameStrobe[0]
port 64 nsew signal input
flabel metal2 s 27066 0 27122 56 0 FreeSans 224 0 0 0 FrameStrobe[10]
port 65 nsew signal input
flabel metal2 s 27342 0 27398 56 0 FreeSans 224 0 0 0 FrameStrobe[11]
port 66 nsew signal input
flabel metal2 s 27618 0 27674 56 0 FreeSans 224 0 0 0 FrameStrobe[12]
port 67 nsew signal input
flabel metal2 s 27894 0 27950 56 0 FreeSans 224 0 0 0 FrameStrobe[13]
port 68 nsew signal input
flabel metal2 s 28170 0 28226 56 0 FreeSans 224 0 0 0 FrameStrobe[14]
port 69 nsew signal input
flabel metal2 s 28446 0 28502 56 0 FreeSans 224 0 0 0 FrameStrobe[15]
port 70 nsew signal input
flabel metal2 s 28722 0 28778 56 0 FreeSans 224 0 0 0 FrameStrobe[16]
port 71 nsew signal input
flabel metal2 s 28998 0 29054 56 0 FreeSans 224 0 0 0 FrameStrobe[17]
port 72 nsew signal input
flabel metal2 s 29274 0 29330 56 0 FreeSans 224 0 0 0 FrameStrobe[18]
port 73 nsew signal input
flabel metal2 s 29550 0 29606 56 0 FreeSans 224 0 0 0 FrameStrobe[19]
port 74 nsew signal input
flabel metal2 s 24582 0 24638 56 0 FreeSans 224 0 0 0 FrameStrobe[1]
port 75 nsew signal input
flabel metal2 s 24858 0 24914 56 0 FreeSans 224 0 0 0 FrameStrobe[2]
port 76 nsew signal input
flabel metal2 s 25134 0 25190 56 0 FreeSans 224 0 0 0 FrameStrobe[3]
port 77 nsew signal input
flabel metal2 s 25410 0 25466 56 0 FreeSans 224 0 0 0 FrameStrobe[4]
port 78 nsew signal input
flabel metal2 s 25686 0 25742 56 0 FreeSans 224 0 0 0 FrameStrobe[5]
port 79 nsew signal input
flabel metal2 s 25962 0 26018 56 0 FreeSans 224 0 0 0 FrameStrobe[6]
port 80 nsew signal input
flabel metal2 s 26238 0 26294 56 0 FreeSans 224 0 0 0 FrameStrobe[7]
port 81 nsew signal input
flabel metal2 s 26514 0 26570 56 0 FreeSans 224 0 0 0 FrameStrobe[8]
port 82 nsew signal input
flabel metal2 s 26790 0 26846 56 0 FreeSans 224 0 0 0 FrameStrobe[9]
port 83 nsew signal input
flabel metal2 s 2778 11194 2834 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[0]
port 84 nsew signal output
flabel metal2 s 18418 11194 18474 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[10]
port 85 nsew signal output
flabel metal2 s 19982 11194 20038 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[11]
port 86 nsew signal output
flabel metal2 s 21546 11194 21602 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[12]
port 87 nsew signal output
flabel metal2 s 23110 11194 23166 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[13]
port 88 nsew signal output
flabel metal2 s 24674 11194 24730 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[14]
port 89 nsew signal output
flabel metal2 s 26238 11194 26294 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[15]
port 90 nsew signal output
flabel metal2 s 27802 11194 27858 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[16]
port 91 nsew signal output
flabel metal2 s 29366 11194 29422 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[17]
port 92 nsew signal output
flabel metal2 s 30930 11194 30986 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[18]
port 93 nsew signal output
flabel metal2 s 32494 11194 32550 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[19]
port 94 nsew signal output
flabel metal2 s 4342 11194 4398 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[1]
port 95 nsew signal output
flabel metal2 s 5906 11194 5962 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[2]
port 96 nsew signal output
flabel metal2 s 7470 11194 7526 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[3]
port 97 nsew signal output
flabel metal2 s 9034 11194 9090 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[4]
port 98 nsew signal output
flabel metal2 s 10598 11194 10654 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[5]
port 99 nsew signal output
flabel metal2 s 12162 11194 12218 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[6]
port 100 nsew signal output
flabel metal2 s 13726 11194 13782 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[7]
port 101 nsew signal output
flabel metal2 s 15290 11194 15346 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[8]
port 102 nsew signal output
flabel metal2 s 16854 11194 16910 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[9]
port 103 nsew signal output
flabel metal2 s 4158 0 4214 56 0 FreeSans 224 0 0 0 N1END[0]
port 104 nsew signal input
flabel metal2 s 4434 0 4490 56 0 FreeSans 224 0 0 0 N1END[1]
port 105 nsew signal input
flabel metal2 s 4710 0 4766 56 0 FreeSans 224 0 0 0 N1END[2]
port 106 nsew signal input
flabel metal2 s 4986 0 5042 56 0 FreeSans 224 0 0 0 N1END[3]
port 107 nsew signal input
flabel metal2 s 7470 0 7526 56 0 FreeSans 224 0 0 0 N2END[0]
port 108 nsew signal input
flabel metal2 s 7746 0 7802 56 0 FreeSans 224 0 0 0 N2END[1]
port 109 nsew signal input
flabel metal2 s 8022 0 8078 56 0 FreeSans 224 0 0 0 N2END[2]
port 110 nsew signal input
flabel metal2 s 8298 0 8354 56 0 FreeSans 224 0 0 0 N2END[3]
port 111 nsew signal input
flabel metal2 s 8574 0 8630 56 0 FreeSans 224 0 0 0 N2END[4]
port 112 nsew signal input
flabel metal2 s 8850 0 8906 56 0 FreeSans 224 0 0 0 N2END[5]
port 113 nsew signal input
flabel metal2 s 9126 0 9182 56 0 FreeSans 224 0 0 0 N2END[6]
port 114 nsew signal input
flabel metal2 s 9402 0 9458 56 0 FreeSans 224 0 0 0 N2END[7]
port 115 nsew signal input
flabel metal2 s 5262 0 5318 56 0 FreeSans 224 0 0 0 N2MID[0]
port 116 nsew signal input
flabel metal2 s 5538 0 5594 56 0 FreeSans 224 0 0 0 N2MID[1]
port 117 nsew signal input
flabel metal2 s 5814 0 5870 56 0 FreeSans 224 0 0 0 N2MID[2]
port 118 nsew signal input
flabel metal2 s 6090 0 6146 56 0 FreeSans 224 0 0 0 N2MID[3]
port 119 nsew signal input
flabel metal2 s 6366 0 6422 56 0 FreeSans 224 0 0 0 N2MID[4]
port 120 nsew signal input
flabel metal2 s 6642 0 6698 56 0 FreeSans 224 0 0 0 N2MID[5]
port 121 nsew signal input
flabel metal2 s 6918 0 6974 56 0 FreeSans 224 0 0 0 N2MID[6]
port 122 nsew signal input
flabel metal2 s 7194 0 7250 56 0 FreeSans 224 0 0 0 N2MID[7]
port 123 nsew signal input
flabel metal2 s 9678 0 9734 56 0 FreeSans 224 0 0 0 N4END[0]
port 124 nsew signal input
flabel metal2 s 12438 0 12494 56 0 FreeSans 224 0 0 0 N4END[10]
port 125 nsew signal input
flabel metal2 s 12714 0 12770 56 0 FreeSans 224 0 0 0 N4END[11]
port 126 nsew signal input
flabel metal2 s 12990 0 13046 56 0 FreeSans 224 0 0 0 N4END[12]
port 127 nsew signal input
flabel metal2 s 13266 0 13322 56 0 FreeSans 224 0 0 0 N4END[13]
port 128 nsew signal input
flabel metal2 s 13542 0 13598 56 0 FreeSans 224 0 0 0 N4END[14]
port 129 nsew signal input
flabel metal2 s 13818 0 13874 56 0 FreeSans 224 0 0 0 N4END[15]
port 130 nsew signal input
flabel metal2 s 9954 0 10010 56 0 FreeSans 224 0 0 0 N4END[1]
port 131 nsew signal input
flabel metal2 s 10230 0 10286 56 0 FreeSans 224 0 0 0 N4END[2]
port 132 nsew signal input
flabel metal2 s 10506 0 10562 56 0 FreeSans 224 0 0 0 N4END[3]
port 133 nsew signal input
flabel metal2 s 10782 0 10838 56 0 FreeSans 224 0 0 0 N4END[4]
port 134 nsew signal input
flabel metal2 s 11058 0 11114 56 0 FreeSans 224 0 0 0 N4END[5]
port 135 nsew signal input
flabel metal2 s 11334 0 11390 56 0 FreeSans 224 0 0 0 N4END[6]
port 136 nsew signal input
flabel metal2 s 11610 0 11666 56 0 FreeSans 224 0 0 0 N4END[7]
port 137 nsew signal input
flabel metal2 s 11886 0 11942 56 0 FreeSans 224 0 0 0 N4END[8]
port 138 nsew signal input
flabel metal2 s 12162 0 12218 56 0 FreeSans 224 0 0 0 N4END[9]
port 139 nsew signal input
flabel metal2 s 14094 0 14150 56 0 FreeSans 224 0 0 0 S1BEG[0]
port 140 nsew signal output
flabel metal2 s 14370 0 14426 56 0 FreeSans 224 0 0 0 S1BEG[1]
port 141 nsew signal output
flabel metal2 s 14646 0 14702 56 0 FreeSans 224 0 0 0 S1BEG[2]
port 142 nsew signal output
flabel metal2 s 14922 0 14978 56 0 FreeSans 224 0 0 0 S1BEG[3]
port 143 nsew signal output
flabel metal2 s 15198 0 15254 56 0 FreeSans 224 0 0 0 S2BEG[0]
port 144 nsew signal output
flabel metal2 s 15474 0 15530 56 0 FreeSans 224 0 0 0 S2BEG[1]
port 145 nsew signal output
flabel metal2 s 15750 0 15806 56 0 FreeSans 224 0 0 0 S2BEG[2]
port 146 nsew signal output
flabel metal2 s 16026 0 16082 56 0 FreeSans 224 0 0 0 S2BEG[3]
port 147 nsew signal output
flabel metal2 s 16302 0 16358 56 0 FreeSans 224 0 0 0 S2BEG[4]
port 148 nsew signal output
flabel metal2 s 16578 0 16634 56 0 FreeSans 224 0 0 0 S2BEG[5]
port 149 nsew signal output
flabel metal2 s 16854 0 16910 56 0 FreeSans 224 0 0 0 S2BEG[6]
port 150 nsew signal output
flabel metal2 s 17130 0 17186 56 0 FreeSans 224 0 0 0 S2BEG[7]
port 151 nsew signal output
flabel metal2 s 17406 0 17462 56 0 FreeSans 224 0 0 0 S2BEGb[0]
port 152 nsew signal output
flabel metal2 s 17682 0 17738 56 0 FreeSans 224 0 0 0 S2BEGb[1]
port 153 nsew signal output
flabel metal2 s 17958 0 18014 56 0 FreeSans 224 0 0 0 S2BEGb[2]
port 154 nsew signal output
flabel metal2 s 18234 0 18290 56 0 FreeSans 224 0 0 0 S2BEGb[3]
port 155 nsew signal output
flabel metal2 s 18510 0 18566 56 0 FreeSans 224 0 0 0 S2BEGb[4]
port 156 nsew signal output
flabel metal2 s 18786 0 18842 56 0 FreeSans 224 0 0 0 S2BEGb[5]
port 157 nsew signal output
flabel metal2 s 19062 0 19118 56 0 FreeSans 224 0 0 0 S2BEGb[6]
port 158 nsew signal output
flabel metal2 s 19338 0 19394 56 0 FreeSans 224 0 0 0 S2BEGb[7]
port 159 nsew signal output
flabel metal2 s 19614 0 19670 56 0 FreeSans 224 0 0 0 S4BEG[0]
port 160 nsew signal output
flabel metal2 s 22374 0 22430 56 0 FreeSans 224 0 0 0 S4BEG[10]
port 161 nsew signal output
flabel metal2 s 22650 0 22706 56 0 FreeSans 224 0 0 0 S4BEG[11]
port 162 nsew signal output
flabel metal2 s 22926 0 22982 56 0 FreeSans 224 0 0 0 S4BEG[12]
port 163 nsew signal output
flabel metal2 s 23202 0 23258 56 0 FreeSans 224 0 0 0 S4BEG[13]
port 164 nsew signal output
flabel metal2 s 23478 0 23534 56 0 FreeSans 224 0 0 0 S4BEG[14]
port 165 nsew signal output
flabel metal2 s 23754 0 23810 56 0 FreeSans 224 0 0 0 S4BEG[15]
port 166 nsew signal output
flabel metal2 s 19890 0 19946 56 0 FreeSans 224 0 0 0 S4BEG[1]
port 167 nsew signal output
flabel metal2 s 20166 0 20222 56 0 FreeSans 224 0 0 0 S4BEG[2]
port 168 nsew signal output
flabel metal2 s 20442 0 20498 56 0 FreeSans 224 0 0 0 S4BEG[3]
port 169 nsew signal output
flabel metal2 s 20718 0 20774 56 0 FreeSans 224 0 0 0 S4BEG[4]
port 170 nsew signal output
flabel metal2 s 20994 0 21050 56 0 FreeSans 224 0 0 0 S4BEG[5]
port 171 nsew signal output
flabel metal2 s 21270 0 21326 56 0 FreeSans 224 0 0 0 S4BEG[6]
port 172 nsew signal output
flabel metal2 s 21546 0 21602 56 0 FreeSans 224 0 0 0 S4BEG[7]
port 173 nsew signal output
flabel metal2 s 21822 0 21878 56 0 FreeSans 224 0 0 0 S4BEG[8]
port 174 nsew signal output
flabel metal2 s 22098 0 22154 56 0 FreeSans 224 0 0 0 S4BEG[9]
port 175 nsew signal output
flabel metal2 s 24030 0 24086 56 0 FreeSans 224 0 0 0 UserCLK
port 176 nsew signal input
flabel metal2 s 1214 11194 1270 11250 0 FreeSans 224 0 0 0 UserCLKo
port 177 nsew signal output
flabel metal4 s 3004 0 3324 11250 0 FreeSans 1920 90 0 0 VGND
port 178 nsew ground bidirectional
flabel metal4 s 3004 0 3324 60 0 FreeSans 480 0 0 0 VGND
port 178 nsew ground bidirectional
flabel metal4 s 3004 11190 3324 11250 0 FreeSans 480 0 0 0 VGND
port 178 nsew ground bidirectional
flabel metal4 s 9004 0 9324 11250 0 FreeSans 1920 90 0 0 VGND
port 178 nsew ground bidirectional
flabel metal4 s 9004 0 9324 60 0 FreeSans 480 0 0 0 VGND
port 178 nsew ground bidirectional
flabel metal4 s 9004 11190 9324 11250 0 FreeSans 480 0 0 0 VGND
port 178 nsew ground bidirectional
flabel metal4 s 15004 0 15324 11250 0 FreeSans 1920 90 0 0 VGND
port 178 nsew ground bidirectional
flabel metal4 s 15004 0 15324 60 0 FreeSans 480 0 0 0 VGND
port 178 nsew ground bidirectional
flabel metal4 s 15004 11190 15324 11250 0 FreeSans 480 0 0 0 VGND
port 178 nsew ground bidirectional
flabel metal4 s 21004 0 21324 11250 0 FreeSans 1920 90 0 0 VGND
port 178 nsew ground bidirectional
flabel metal4 s 21004 0 21324 60 0 FreeSans 480 0 0 0 VGND
port 178 nsew ground bidirectional
flabel metal4 s 21004 11190 21324 11250 0 FreeSans 480 0 0 0 VGND
port 178 nsew ground bidirectional
flabel metal4 s 27004 0 27324 11250 0 FreeSans 1920 90 0 0 VGND
port 178 nsew ground bidirectional
flabel metal4 s 27004 0 27324 60 0 FreeSans 480 0 0 0 VGND
port 178 nsew ground bidirectional
flabel metal4 s 27004 11190 27324 11250 0 FreeSans 480 0 0 0 VGND
port 178 nsew ground bidirectional
flabel metal4 s 1944 0 2264 11250 0 FreeSans 1920 90 0 0 VPWR
port 179 nsew power bidirectional
flabel metal4 s 1944 0 2264 60 0 FreeSans 480 0 0 0 VPWR
port 179 nsew power bidirectional
flabel metal4 s 1944 11190 2264 11250 0 FreeSans 480 0 0 0 VPWR
port 179 nsew power bidirectional
flabel metal4 s 7944 0 8264 11250 0 FreeSans 1920 90 0 0 VPWR
port 179 nsew power bidirectional
flabel metal4 s 7944 0 8264 60 0 FreeSans 480 0 0 0 VPWR
port 179 nsew power bidirectional
flabel metal4 s 7944 11190 8264 11250 0 FreeSans 480 0 0 0 VPWR
port 179 nsew power bidirectional
flabel metal4 s 13944 0 14264 11250 0 FreeSans 1920 90 0 0 VPWR
port 179 nsew power bidirectional
flabel metal4 s 13944 0 14264 60 0 FreeSans 480 0 0 0 VPWR
port 179 nsew power bidirectional
flabel metal4 s 13944 11190 14264 11250 0 FreeSans 480 0 0 0 VPWR
port 179 nsew power bidirectional
flabel metal4 s 19944 0 20264 11250 0 FreeSans 1920 90 0 0 VPWR
port 179 nsew power bidirectional
flabel metal4 s 19944 0 20264 60 0 FreeSans 480 0 0 0 VPWR
port 179 nsew power bidirectional
flabel metal4 s 19944 11190 20264 11250 0 FreeSans 480 0 0 0 VPWR
port 179 nsew power bidirectional
flabel metal4 s 25944 0 26264 11250 0 FreeSans 1920 90 0 0 VPWR
port 179 nsew power bidirectional
flabel metal4 s 25944 0 26264 60 0 FreeSans 480 0 0 0 VPWR
port 179 nsew power bidirectional
flabel metal4 s 25944 11190 26264 11250 0 FreeSans 480 0 0 0 VPWR
port 179 nsew power bidirectional
flabel metal4 s 31944 0 32264 11250 0 FreeSans 1920 90 0 0 VPWR
port 179 nsew power bidirectional
flabel metal4 s 31944 0 32264 60 0 FreeSans 480 0 0 0 VPWR
port 179 nsew power bidirectional
flabel metal4 s 31944 11190 32264 11250 0 FreeSans 480 0 0 0 VPWR
port 179 nsew power bidirectional
rlabel metal1 16836 8704 16836 8704 0 VGND
rlabel metal1 16836 8160 16836 8160 0 VPWR
rlabel metal2 17434 3553 17434 3553 0 FrameData[0]
rlabel metal1 23092 4998 23092 4998 0 FrameData[10]
rlabel metal3 1471 4420 1471 4420 0 FrameData[11]
rlabel metal2 19366 5661 19366 5661 0 FrameData[12]
rlabel metal3 919 4964 919 4964 0 FrameData[13]
rlabel metal3 6002 5236 6002 5236 0 FrameData[14]
rlabel metal3 1471 5508 1471 5508 0 FrameData[15]
rlabel metal3 6922 5780 6922 5780 0 FrameData[16]
rlabel metal3 919 6052 919 6052 0 FrameData[17]
rlabel metal3 2828 6324 2828 6324 0 FrameData[18]
rlabel metal3 1471 6596 1471 6596 0 FrameData[19]
rlabel metal2 20470 3196 20470 3196 0 FrameData[1]
rlabel metal3 3196 6868 3196 6868 0 FrameData[20]
rlabel metal3 919 7140 919 7140 0 FrameData[21]
rlabel metal1 16836 7378 16836 7378 0 FrameData[22]
rlabel metal3 1471 7684 1471 7684 0 FrameData[23]
rlabel metal2 14582 7667 14582 7667 0 FrameData[24]
rlabel metal3 919 8228 919 8228 0 FrameData[25]
rlabel metal3 735 8500 735 8500 0 FrameData[26]
rlabel metal3 1471 8772 1471 8772 0 FrameData[27]
rlabel metal2 12466 8211 12466 8211 0 FrameData[28]
rlabel metal3 2460 9316 2460 9316 0 FrameData[29]
rlabel metal1 21896 3502 21896 3502 0 FrameData[2]
rlabel metal2 7774 8381 7774 8381 0 FrameData[30]
rlabel metal2 17158 8653 17158 8653 0 FrameData[31]
rlabel metal3 1494 2244 1494 2244 0 FrameData[3]
rlabel metal1 19688 4114 19688 4114 0 FrameData[4]
rlabel metal3 919 2788 919 2788 0 FrameData[5]
rlabel metal2 25806 3213 25806 3213 0 FrameData[6]
rlabel metal3 1471 3332 1471 3332 0 FrameData[7]
rlabel metal2 13110 4029 13110 4029 0 FrameData[8]
rlabel metal3 919 3876 919 3876 0 FrameData[9]
rlabel metal3 32585 1428 32585 1428 0 FrameData_O[0]
rlabel metal3 32723 4148 32723 4148 0 FrameData_O[10]
rlabel metal3 32907 4420 32907 4420 0 FrameData_O[11]
rlabel metal2 31510 4845 31510 4845 0 FrameData_O[12]
rlabel metal3 33275 4964 33275 4964 0 FrameData_O[13]
rlabel metal3 32861 5236 32861 5236 0 FrameData_O[14]
rlabel metal3 32723 5508 32723 5508 0 FrameData_O[15]
rlabel metal3 32907 5780 32907 5780 0 FrameData_O[16]
rlabel metal3 33160 6052 33160 6052 0 FrameData_O[17]
rlabel metal3 32769 6324 32769 6324 0 FrameData_O[18]
rlabel via2 31418 6613 31418 6613 0 FrameData_O[19]
rlabel metal3 32401 1700 32401 1700 0 FrameData_O[1]
rlabel metal2 31786 6749 31786 6749 0 FrameData_O[20]
rlabel metal3 33229 7140 33229 7140 0 FrameData_O[21]
rlabel metal3 32723 7412 32723 7412 0 FrameData_O[22]
rlabel metal3 32907 7684 32907 7684 0 FrameData_O[23]
rlabel metal3 32769 7956 32769 7956 0 FrameData_O[24]
rlabel metal3 33045 8228 33045 8228 0 FrameData_O[25]
rlabel metal2 31418 8279 31418 8279 0 FrameData_O[26]
rlabel metal2 31050 8415 31050 8415 0 FrameData_O[27]
rlabel metal2 30498 8823 30498 8823 0 FrameData_O[28]
rlabel metal2 31510 8415 31510 8415 0 FrameData_O[29]
rlabel metal3 32217 1972 32217 1972 0 FrameData_O[2]
rlabel metal1 30774 8058 30774 8058 0 FrameData_O[30]
rlabel metal2 30130 9231 30130 9231 0 FrameData_O[31]
rlabel metal3 32769 2244 32769 2244 0 FrameData_O[3]
rlabel metal3 32723 2516 32723 2516 0 FrameData_O[4]
rlabel metal3 33275 2788 33275 2788 0 FrameData_O[5]
rlabel metal3 32723 3060 32723 3060 0 FrameData_O[6]
rlabel metal3 32907 3332 32907 3332 0 FrameData_O[7]
rlabel metal2 31510 3757 31510 3757 0 FrameData_O[8]
rlabel metal3 33275 3876 33275 3876 0 FrameData_O[9]
rlabel metal1 24380 7378 24380 7378 0 FrameStrobe[0]
rlabel metal1 20654 6256 20654 6256 0 FrameStrobe[10]
rlabel metal1 21206 5644 21206 5644 0 FrameStrobe[11]
rlabel metal1 25024 3570 25024 3570 0 FrameStrobe[12]
rlabel metal1 25622 3706 25622 3706 0 FrameStrobe[13]
rlabel metal1 25852 4046 25852 4046 0 FrameStrobe[14]
rlabel metal1 26174 4114 26174 4114 0 FrameStrobe[15]
rlabel metal1 26956 4522 26956 4522 0 FrameStrobe[16]
rlabel metal2 29026 1347 29026 1347 0 FrameStrobe[17]
rlabel metal1 29164 5678 29164 5678 0 FrameStrobe[18]
rlabel metal1 30130 5678 30130 5678 0 FrameStrobe[19]
rlabel metal2 20930 7140 20930 7140 0 FrameStrobe[1]
rlabel metal2 24886 1347 24886 1347 0 FrameStrobe[2]
rlabel metal1 20562 6188 20562 6188 0 FrameStrobe[3]
rlabel metal2 25438 684 25438 684 0 FrameStrobe[4]
rlabel metal1 24426 7446 24426 7446 0 FrameStrobe[5]
rlabel metal2 25990 735 25990 735 0 FrameStrobe[6]
rlabel metal2 26266 803 26266 803 0 FrameStrobe[7]
rlabel metal1 25208 5202 25208 5202 0 FrameStrobe[8]
rlabel metal1 26496 5542 26496 5542 0 FrameStrobe[9]
rlabel metal1 2898 8602 2898 8602 0 FrameStrobe_O[0]
rlabel metal1 18538 8602 18538 8602 0 FrameStrobe_O[10]
rlabel metal1 20102 8602 20102 8602 0 FrameStrobe_O[11]
rlabel metal1 21758 8602 21758 8602 0 FrameStrobe_O[12]
rlabel metal1 23276 8602 23276 8602 0 FrameStrobe_O[13]
rlabel metal1 24840 8602 24840 8602 0 FrameStrobe_O[14]
rlabel metal1 26404 8602 26404 8602 0 FrameStrobe_O[15]
rlabel metal1 27968 8602 27968 8602 0 FrameStrobe_O[16]
rlabel metal1 29578 8602 29578 8602 0 FrameStrobe_O[17]
rlabel metal1 31096 8602 31096 8602 0 FrameStrobe_O[18]
rlabel metal1 32246 6630 32246 6630 0 FrameStrobe_O[19]
rlabel metal1 4462 8602 4462 8602 0 FrameStrobe_O[1]
rlabel metal1 6210 8602 6210 8602 0 FrameStrobe_O[2]
rlabel metal1 7590 8602 7590 8602 0 FrameStrobe_O[3]
rlabel metal1 9062 8602 9062 8602 0 FrameStrobe_O[4]
rlabel metal1 10718 8602 10718 8602 0 FrameStrobe_O[5]
rlabel metal1 12282 8602 12282 8602 0 FrameStrobe_O[6]
rlabel metal1 13984 8602 13984 8602 0 FrameStrobe_O[7]
rlabel metal1 15456 8602 15456 8602 0 FrameStrobe_O[8]
rlabel metal1 16974 8602 16974 8602 0 FrameStrobe_O[9]
rlabel metal2 4186 2622 4186 2622 0 N1END[0]
rlabel metal2 4462 3166 4462 3166 0 N1END[1]
rlabel metal2 4738 3370 4738 3370 0 N1END[2]
rlabel metal2 5014 2588 5014 2588 0 N1END[3]
rlabel metal2 4738 7174 4738 7174 0 N2END[0]
rlabel metal1 6026 7344 6026 7344 0 N2END[1]
rlabel metal2 8050 55 8050 55 0 N2END[2]
rlabel metal2 8326 3404 8326 3404 0 N2END[3]
rlabel metal2 8602 3166 8602 3166 0 N2END[4]
rlabel metal2 8878 2860 8878 2860 0 N2END[5]
rlabel metal2 9154 55 9154 55 0 N2END[6]
rlabel metal2 9430 55 9430 55 0 N2END[7]
rlabel metal2 5290 2316 5290 2316 0 N2MID[0]
rlabel metal2 5566 2860 5566 2860 0 N2MID[1]
rlabel metal2 5842 3404 5842 3404 0 N2MID[2]
rlabel metal1 6394 7514 6394 7514 0 N2MID[3]
rlabel metal2 6394 3370 6394 3370 0 N2MID[4]
rlabel metal2 6670 2316 6670 2316 0 N2MID[5]
rlabel metal2 6946 2282 6946 2282 0 N2MID[6]
rlabel metal2 7222 2248 7222 2248 0 N2MID[7]
rlabel metal1 19826 3434 19826 3434 0 N4END[0]
rlabel metal1 13524 3434 13524 3434 0 N4END[10]
rlabel metal1 12926 3978 12926 3978 0 N4END[11]
rlabel metal1 12880 4114 12880 4114 0 N4END[12]
rlabel metal1 12880 2822 12880 2822 0 N4END[13]
rlabel metal1 13248 2890 13248 2890 0 N4END[14]
rlabel metal1 13156 3502 13156 3502 0 N4END[15]
rlabel metal2 19412 2924 19412 2924 0 N4END[1]
rlabel metal1 19136 3978 19136 3978 0 N4END[2]
rlabel metal2 10534 667 10534 667 0 N4END[3]
rlabel metal2 10810 1211 10810 1211 0 N4END[4]
rlabel metal2 11086 650 11086 650 0 N4END[5]
rlabel metal2 11362 1058 11362 1058 0 N4END[6]
rlabel metal2 11638 1568 11638 1568 0 N4END[7]
rlabel metal2 11914 2350 11914 2350 0 N4END[8]
rlabel metal2 12190 1806 12190 1806 0 N4END[9]
rlabel metal2 14122 1160 14122 1160 0 S1BEG[0]
rlabel metal1 14536 2822 14536 2822 0 S1BEG[1]
rlabel metal2 14674 1160 14674 1160 0 S1BEG[2]
rlabel metal2 14950 1160 14950 1160 0 S1BEG[3]
rlabel metal1 15456 2822 15456 2822 0 S2BEG[0]
rlabel metal2 15502 1160 15502 1160 0 S2BEG[1]
rlabel metal2 15778 1160 15778 1160 0 S2BEG[2]
rlabel metal1 16192 2822 16192 2822 0 S2BEG[3]
rlabel metal2 16330 1160 16330 1160 0 S2BEG[4]
rlabel metal2 16606 1160 16606 1160 0 S2BEG[5]
rlabel metal2 16882 1160 16882 1160 0 S2BEG[6]
rlabel metal2 17158 1160 17158 1160 0 S2BEG[7]
rlabel metal2 17434 1160 17434 1160 0 S2BEGb[0]
rlabel metal2 17710 1330 17710 1330 0 S2BEGb[1]
rlabel metal2 17986 1160 17986 1160 0 S2BEGb[2]
rlabel metal2 18262 1296 18262 1296 0 S2BEGb[3]
rlabel metal2 18538 1160 18538 1160 0 S2BEGb[4]
rlabel metal2 18814 55 18814 55 0 S2BEGb[5]
rlabel metal2 19090 718 19090 718 0 S2BEGb[6]
rlabel metal1 19504 2822 19504 2822 0 S2BEGb[7]
rlabel metal2 19642 1160 19642 1160 0 S4BEG[0]
rlabel metal2 22402 599 22402 599 0 S4BEG[10]
rlabel metal1 22816 2822 22816 2822 0 S4BEG[11]
rlabel metal2 22954 1296 22954 1296 0 S4BEG[12]
rlabel metal1 23368 2822 23368 2822 0 S4BEG[13]
rlabel metal2 23506 1160 23506 1160 0 S4BEG[14]
rlabel metal1 23920 2822 23920 2822 0 S4BEG[15]
rlabel metal2 19918 1296 19918 1296 0 S4BEG[1]
rlabel metal2 20194 599 20194 599 0 S4BEG[2]
rlabel metal1 20608 2822 20608 2822 0 S4BEG[3]
rlabel metal1 20976 2822 20976 2822 0 S4BEG[4]
rlabel metal2 21022 55 21022 55 0 S4BEG[5]
rlabel metal2 21298 55 21298 55 0 S4BEG[6]
rlabel metal1 21804 2822 21804 2822 0 S4BEG[7]
rlabel metal2 21850 1296 21850 1296 0 S4BEG[8]
rlabel metal2 22126 1160 22126 1160 0 S4BEG[9]
rlabel metal1 24518 7310 24518 7310 0 UserCLK
rlabel metal1 1334 8602 1334 8602 0 UserCLKo
rlabel metal1 18262 3910 18262 3910 0 net1
rlabel metal2 9522 6936 9522 6936 0 net10
rlabel metal1 17158 6800 17158 6800 0 net11
rlabel metal2 20838 3264 20838 3264 0 net12
rlabel metal2 17066 6596 17066 6596 0 net13
rlabel metal2 7590 7684 7590 7684 0 net14
rlabel metal2 16882 7446 16882 7446 0 net15
rlabel metal2 7038 7582 7038 7582 0 net16
rlabel metal1 21390 8432 21390 8432 0 net17
rlabel metal2 14214 7565 14214 7565 0 net18
rlabel metal2 16422 7718 16422 7718 0 net19
rlabel metal1 31602 4624 31602 4624 0 net2
rlabel metal2 12374 7072 12374 7072 0 net20
rlabel metal1 12604 7174 12604 7174 0 net21
rlabel via2 5934 7259 5934 7259 0 net22
rlabel metal1 30590 2482 30590 2482 0 net23
rlabel metal1 16560 7344 16560 7344 0 net24
rlabel metal2 17526 8058 17526 8058 0 net25
rlabel metal1 21666 3400 21666 3400 0 net26
rlabel metal2 31326 3468 31326 3468 0 net27
rlabel metal2 31694 3196 31694 3196 0 net28
rlabel metal1 31602 3468 31602 3468 0 net29
rlabel metal2 31878 5338 31878 5338 0 net3
rlabel metal1 31970 3570 31970 3570 0 net30
rlabel metal2 31326 4284 31326 4284 0 net31
rlabel metal2 19826 4777 19826 4777 0 net32
rlabel metal2 5014 8670 5014 8670 0 net33
rlabel metal1 19642 6154 19642 6154 0 net34
rlabel metal1 20700 5542 20700 5542 0 net35
rlabel metal2 22218 6222 22218 6222 0 net36
rlabel metal2 23138 6222 23138 6222 0 net37
rlabel metal2 23690 6222 23690 6222 0 net38
rlabel metal1 25254 3978 25254 3978 0 net39
rlabel metal2 19734 6528 19734 6528 0 net4
rlabel metal2 25070 6596 25070 6596 0 net40
rlabel metal1 28106 5338 28106 5338 0 net41
rlabel metal1 29854 5814 29854 5814 0 net42
rlabel metal1 31280 5542 31280 5542 0 net43
rlabel metal1 4738 8908 4738 8908 0 net44
rlabel metal2 20286 7752 20286 7752 0 net45
rlabel metal2 14306 7446 14306 7446 0 net46
rlabel metal1 19734 7480 19734 7480 0 net47
rlabel metal2 22954 8160 22954 8160 0 net48
rlabel metal2 17342 9248 17342 9248 0 net49
rlabel metal1 18354 6630 18354 6630 0 net5
rlabel metal2 16790 9112 16790 9112 0 net50
rlabel metal2 17066 8636 17066 8636 0 net51
rlabel metal1 21528 5542 21528 5542 0 net52
rlabel metal1 12236 4998 12236 4998 0 net53
rlabel metal2 8234 6528 8234 6528 0 net54
rlabel metal2 9614 4284 9614 4284 0 net55
rlabel metal2 9522 3808 9522 3808 0 net56
rlabel metal1 15364 3026 15364 3026 0 net57
rlabel metal1 13754 4794 13754 4794 0 net58
rlabel metal1 12282 4726 12282 4726 0 net59
rlabel metal2 12098 6528 12098 6528 0 net6
rlabel metal1 12650 6630 12650 6630 0 net60
rlabel metal2 12788 5372 12788 5372 0 net61
rlabel metal2 5934 6426 5934 6426 0 net62
rlabel metal1 5451 5542 5451 5542 0 net63
rlabel metal2 7130 4352 7130 4352 0 net64
rlabel metal2 14306 3740 14306 3740 0 net65
rlabel metal1 14628 3706 14628 3706 0 net66
rlabel metal1 14582 5542 14582 5542 0 net67
rlabel metal2 17802 4454 17802 4454 0 net68
rlabel metal1 8832 6630 8832 6630 0 net69
rlabel metal2 13110 6460 13110 6460 0 net7
rlabel metal1 7912 5542 7912 5542 0 net70
rlabel metal2 6210 4556 6210 4556 0 net71
rlabel metal2 19458 4012 19458 4012 0 net72
rlabel metal1 14306 3366 14306 3366 0 net73
rlabel metal2 23322 2210 23322 2210 0 net74
rlabel metal2 17342 3808 17342 3808 0 net75
rlabel metal2 23690 2244 23690 2244 0 net76
rlabel metal2 19826 3434 19826 3434 0 net77
rlabel metal1 24104 2414 24104 2414 0 net78
rlabel metal2 20286 3230 20286 3230 0 net79
rlabel metal1 15318 7242 15318 7242 0 net8
rlabel metal1 20562 2380 20562 2380 0 net80
rlabel metal2 19918 3264 19918 3264 0 net81
rlabel metal2 18538 3536 18538 3536 0 net82
rlabel metal1 18814 3978 18814 3978 0 net83
rlabel metal2 14674 3672 14674 3672 0 net84
rlabel metal2 14398 3536 14398 3536 0 net85
rlabel metal2 20378 3944 20378 3944 0 net86
rlabel metal1 19274 3536 19274 3536 0 net87
rlabel metal2 17250 3536 17250 3536 0 net88
rlabel via2 1610 8483 1610 8483 0 net89
rlabel metal2 18170 7684 18170 7684 0 net9
<< properties >>
string FIXED_BBOX 0 0 33750 11250
<< end >>
