module LUT4AB (Ci,
    Co,
    UserCLK,
    UserCLKo,
    E1BEG,
    E1END,
    E2BEG,
    E2BEGb,
    E2END,
    E2MID,
    E6BEG,
    E6END,
    EE4BEG,
    EE4END,
    FrameData,
    FrameData_O,
    FrameStrobe,
    FrameStrobe_O,
    N1BEG,
    N1END,
    N2BEG,
    N2BEGb,
    N2END,
    N2MID,
    N4BEG,
    N4END,
    NN4BEG,
    NN4END,
    S1BEG,
    S1END,
    S2BEG,
    S2BEGb,
    S2END,
    S2MID,
    S4BEG,
    S4END,
    SS4BEG,
    SS4END,
    W1BEG,
    W1END,
    W2BEG,
    W2BEGb,
    W2END,
    W2MID,
    W6BEG,
    W6END,
    WW4BEG,
    WW4END);
 input Ci;
 output Co;
 input UserCLK;
 output UserCLKo;
 output [3:0] E1BEG;
 input [3:0] E1END;
 output [7:0] E2BEG;
 output [7:0] E2BEGb;
 input [7:0] E2END;
 input [7:0] E2MID;
 output [11:0] E6BEG;
 input [11:0] E6END;
 output [15:0] EE4BEG;
 input [15:0] EE4END;
 input [31:0] FrameData;
 output [31:0] FrameData_O;
 input [19:0] FrameStrobe;
 output [19:0] FrameStrobe_O;
 output [3:0] N1BEG;
 input [3:0] N1END;
 output [7:0] N2BEG;
 output [7:0] N2BEGb;
 input [7:0] N2END;
 input [7:0] N2MID;
 output [15:0] N4BEG;
 input [15:0] N4END;
 output [15:0] NN4BEG;
 input [15:0] NN4END;
 output [3:0] S1BEG;
 input [3:0] S1END;
 output [7:0] S2BEG;
 output [7:0] S2BEGb;
 input [7:0] S2END;
 input [7:0] S2MID;
 output [15:0] S4BEG;
 input [15:0] S4END;
 output [15:0] SS4BEG;
 input [15:0] SS4END;
 output [3:0] W1BEG;
 input [3:0] W1END;
 output [7:0] W2BEG;
 output [7:0] W2BEGb;
 input [7:0] W2END;
 input [7:0] W2MID;
 output [11:0] W6BEG;
 input [11:0] W6END;
 output [15:0] WW4BEG;
 input [15:0] WW4END;

 wire A;
 wire B;
 wire C;
 wire net112;
 wire D;
 wire E;
 wire net113;
 wire net114;
 wire net397;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net123;
 wire net396;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net386;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net392;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire F;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire G;
 wire H;
 wire \Inst_LA_LUT4c_frame_config_dffesr.LUT_flop ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.c_I0mux ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.c_out_mux ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.c_reset_value ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.LUT_flop ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.c_I0mux ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.c_out_mux ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.c_reset_value ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.LUT_flop ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.c_I0mux ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.c_out_mux ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.c_reset_value ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.LUT_flop ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.c_I0mux ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.c_out_mux ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.c_reset_value ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.LUT_flop ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.c_I0mux ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.c_out_mux ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.c_reset_value ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.LUT_flop ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.c_I0mux ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.c_out_mux ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.c_reset_value ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.LUT_flop ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.c_I0mux ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.c_out_mux ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.c_reset_value ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.LUT_flop ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.c_I0mux ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.c_out_mux ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.c_reset_value ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit9.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit9.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit9.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit9.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit9.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit9.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit9.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit9.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit9.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit9.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit9.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit9.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit9.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit9.Q ;
 wire \Inst_LUT4AB_switch_matrix.E1BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.E1BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.E1BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.E1BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.E2BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.E2BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.E2BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.E2BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.E2BEG4 ;
 wire \Inst_LUT4AB_switch_matrix.E2BEG5 ;
 wire \Inst_LUT4AB_switch_matrix.E2BEG6 ;
 wire \Inst_LUT4AB_switch_matrix.E2BEG7 ;
 wire \Inst_LUT4AB_switch_matrix.E6BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.E6BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.EE4BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.EE4BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.EE4BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.EE4BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.JN2BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.JN2BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.JN2BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.JN2BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.JN2BEG4 ;
 wire \Inst_LUT4AB_switch_matrix.JN2BEG5 ;
 wire \Inst_LUT4AB_switch_matrix.JN2BEG6 ;
 wire \Inst_LUT4AB_switch_matrix.JN2BEG7 ;
 wire \Inst_LUT4AB_switch_matrix.JS2BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.JS2BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.JS2BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.JS2BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.JS2BEG4 ;
 wire \Inst_LUT4AB_switch_matrix.JS2BEG5 ;
 wire \Inst_LUT4AB_switch_matrix.JS2BEG6 ;
 wire \Inst_LUT4AB_switch_matrix.JS2BEG7 ;
 wire \Inst_LUT4AB_switch_matrix.JW2BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.JW2BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.JW2BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.JW2BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.JW2BEG4 ;
 wire \Inst_LUT4AB_switch_matrix.JW2BEG5 ;
 wire \Inst_LUT4AB_switch_matrix.JW2BEG6 ;
 wire \Inst_LUT4AB_switch_matrix.JW2BEG7 ;
 wire \Inst_LUT4AB_switch_matrix.M_AB ;
 wire \Inst_LUT4AB_switch_matrix.M_AD ;
 wire \Inst_LUT4AB_switch_matrix.M_AH ;
 wire \Inst_LUT4AB_switch_matrix.M_EF ;
 wire \Inst_LUT4AB_switch_matrix.N1BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.N1BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.N1BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.N1BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.N4BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.N4BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.N4BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.N4BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.NN4BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.NN4BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.NN4BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.NN4BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.S1BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.S1BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.S1BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.S1BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.S4BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.S4BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.S4BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.S4BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.SS4BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.SS4BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.SS4BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.SS4BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.W1BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.W1BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.W1BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.W1BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.W6BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.W6BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.WW4BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.WW4BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.WW4BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.WW4BEG3 ;
 wire net214;
 wire net395;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net391;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net393;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net394;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net390;
 wire net305;
 wire net306;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net380;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net366;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net387;
 wire net388;
 wire net389;

 sg13g2_inv_1 _1179_ (.Y(_1012_),
    .A(net51));
 sg13g2_inv_1 _1180_ (.Y(_1013_),
    .A(net4));
 sg13g2_inv_1 _1181_ (.Y(_1014_),
    .A(net1213));
 sg13g2_inv_1 _1182_ (.Y(_1015_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit8.Q ));
 sg13g2_inv_1 _1183_ (.Y(_1016_),
    .A(net1217));
 sg13g2_inv_1 _1184_ (.Y(_1017_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit7.Q ));
 sg13g2_inv_1 _1185_ (.Y(_1018_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit8.Q ));
 sg13g2_inv_1 _1186_ (.Y(_1019_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit9.Q ));
 sg13g2_inv_1 _1187_ (.Y(_1020_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit0.Q ));
 sg13g2_inv_1 _1188_ (.Y(_1021_),
    .A(net47));
 sg13g2_inv_1 _1189_ (.Y(_1022_),
    .A(net79));
 sg13g2_inv_1 _1190_ (.Y(_1023_),
    .A(net110));
 sg13g2_inv_1 _1191_ (.Y(_1024_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit8.Q ));
 sg13g2_inv_1 _1192_ (.Y(_1025_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit9.Q ));
 sg13g2_inv_1 _1193_ (.Y(_1026_),
    .A(net102));
 sg13g2_inv_1 _1194_ (.Y(_1027_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit0.Q ));
 sg13g2_inv_1 _1195_ (.Y(_1028_),
    .A(net107));
 sg13g2_inv_1 _1196_ (.Y(_1029_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit9.Q ));
 sg13g2_inv_1 _1197_ (.Y(_1030_),
    .A(net109));
 sg13g2_inv_1 _1198_ (.Y(_1031_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit4.Q ));
 sg13g2_inv_1 _1199_ (.Y(_1032_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit4.Q ));
 sg13g2_inv_1 _1200_ (.Y(_1033_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit5.Q ));
 sg13g2_inv_1 _1201_ (.Y(_1034_),
    .A(net75));
 sg13g2_inv_1 _1202_ (.Y(_1035_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit13.Q ));
 sg13g2_inv_1 _1203_ (.Y(_1036_),
    .A(net80));
 sg13g2_inv_1 _1204_ (.Y(_1037_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit4.Q ));
 sg13g2_inv_1 _1205_ (.Y(_1038_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit5.Q ));
 sg13g2_inv_1 _1206_ (.Y(_1039_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit12.Q ));
 sg13g2_inv_1 _1207_ (.Y(_1040_),
    .A(net25));
 sg13g2_inv_1 _1208_ (.Y(_1041_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit13.Q ));
 sg13g2_inv_1 _1209_ (.Y(_1042_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit16.Q ));
 sg13g2_inv_1 _1210_ (.Y(_1043_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit18.Q ));
 sg13g2_inv_1 _1211_ (.Y(_1044_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit20.Q ));
 sg13g2_inv_1 _1212_ (.Y(_1045_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit24.Q ));
 sg13g2_inv_1 _1213_ (.Y(_1046_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit25.Q ));
 sg13g2_inv_1 _1214_ (.Y(_1047_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit21.Q ));
 sg13g2_inv_1 _1215_ (.Y(_1048_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit19.Q ));
 sg13g2_inv_1 _1216_ (.Y(_1049_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit8.Q ));
 sg13g2_inv_1 _1217_ (.Y(_1050_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit7.Q ));
 sg13g2_inv_16 _1218_ (.A(net951),
    .Y(_1051_));
 sg13g2_inv_1 _1219_ (.Y(_1052_),
    .A(net935));
 sg13g2_mux4_1 _1220_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit30.Q ),
    .A0(net957),
    .A1(net950),
    .A2(net935),
    .A3(net930),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit31.Q ),
    .X(_1053_));
 sg13g2_mux4_1 _1221_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit31.Q ),
    .A0(net975),
    .A1(net945),
    .A2(net940),
    .A3(net962),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit30.Q ),
    .X(_1054_));
 sg13g2_mux2_1 _1222_ (.A0(_1053_),
    .A1(_1054_),
    .S(_1020_),
    .X(_1055_));
 sg13g2_nand2_2 _1223_ (.Y(_1056_),
    .A(_1055_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit1.Q ));
 sg13g2_mux4_1 _1224_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit30.Q ),
    .A0(net31),
    .A1(net37),
    .A2(net53),
    .A3(net8),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit31.Q ),
    .X(_1057_));
 sg13g2_nor2_1 _1225_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit0.Q ),
    .B(_1057_),
    .Y(_1058_));
 sg13g2_mux2_1 _1226_ (.A0(net1212),
    .A1(net65),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit30.Q ),
    .X(_1059_));
 sg13g2_nand2b_1 _1227_ (.Y(_1060_),
    .B(_1059_),
    .A_N(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit31.Q ));
 sg13g2_mux2_1 _1228_ (.A0(net92),
    .A1(net111),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit30.Q ),
    .X(_1061_));
 sg13g2_a21oi_1 _1229_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit31.Q ),
    .A2(_1061_),
    .Y(_1062_),
    .B1(_1020_));
 sg13g2_a21o_1 _1230_ (.A2(_1062_),
    .A1(_1060_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit1.Q ),
    .X(_1063_));
 sg13g2_o21ai_1 _1231_ (.B1(_1056_),
    .Y(\Inst_LUT4AB_switch_matrix.E2BEG1 ),
    .A1(_1058_),
    .A2(_1063_));
 sg13g2_inv_1 _1232_ (.Y(_1064_),
    .A(net383));
 sg13g2_mux4_1 _1233_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit28.Q ),
    .A0(net24),
    .A1(net81),
    .A2(net97),
    .A3(\Inst_LUT4AB_switch_matrix.E2BEG1 ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit29.Q ),
    .X(_1065_));
 sg13g2_mux4_1 _1234_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit29.Q ),
    .A0(net55),
    .A1(net65),
    .A2(net8),
    .A3(net92),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit28.Q ),
    .X(_1066_));
 sg13g2_mux2_1 _1235_ (.A0(net934),
    .A1(net928),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit6.Q ),
    .X(_1067_));
 sg13g2_nand2_2 _1236_ (.Y(_1068_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit7.Q ),
    .B(_1067_));
 sg13g2_mux2_1 _1237_ (.A0(net956),
    .A1(net950),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit6.Q ),
    .X(_1069_));
 sg13g2_a21oi_1 _1238_ (.A1(_1017_),
    .A2(_1069_),
    .Y(_1070_),
    .B1(_1018_));
 sg13g2_mux2_1 _1239_ (.A0(net939),
    .A1(net961),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit6.Q ),
    .X(_1071_));
 sg13g2_nand2_1 _1240_ (.Y(_1072_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit7.Q ),
    .B(_1071_));
 sg13g2_mux2_1 _1241_ (.A0(net974),
    .A1(net968),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit6.Q ),
    .X(_1073_));
 sg13g2_a21oi_1 _1242_ (.A1(_1017_),
    .A2(_1073_),
    .Y(_1074_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit8.Q ));
 sg13g2_a221oi_1 _1243_ (.B2(_1074_),
    .C1(_1019_),
    .B1(_1072_),
    .A1(_1070_),
    .Y(_1075_),
    .A2(_1068_));
 sg13g2_mux4_1 _1244_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit6.Q ),
    .A0(net1008),
    .A1(net39),
    .A2(net51),
    .A3(net10),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit7.Q ),
    .X(_1076_));
 sg13g2_nor2_1 _1245_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit8.Q ),
    .B(_1076_),
    .Y(_1077_));
 sg13g2_mux2_1 _1246_ (.A0(net94),
    .A1(net106),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit6.Q ),
    .X(_1078_));
 sg13g2_mux2_1 _1247_ (.A0(net1212),
    .A1(net67),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit6.Q ),
    .X(_1079_));
 sg13g2_nand2_1 _1248_ (.Y(_1080_),
    .A(_1017_),
    .B(_1079_));
 sg13g2_a21oi_1 _1249_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit7.Q ),
    .A2(_1078_),
    .Y(_1081_),
    .B1(_1018_));
 sg13g2_a21oi_1 _1250_ (.A1(_1080_),
    .A2(_1081_),
    .Y(_1082_),
    .B1(_1077_));
 sg13g2_a21o_2 _1251_ (.A2(_1082_),
    .A1(_1019_),
    .B1(_1075_),
    .X(\Inst_LUT4AB_switch_matrix.E2BEG3 ));
 sg13g2_mux4_1 _1252_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit28.Q ),
    .A0(net16),
    .A1(net73),
    .A2(net100),
    .A3(\Inst_LUT4AB_switch_matrix.E2BEG3 ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit29.Q ),
    .X(_1083_));
 sg13g2_mux4_1 _1253_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit28.Q ),
    .A0(net46),
    .A1(net17),
    .A2(net74),
    .A3(net101),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit29.Q ),
    .X(_1084_));
 sg13g2_mux4_1 _1254_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit5.Q ),
    .A0(_1083_),
    .A1(_1084_),
    .A2(_1066_),
    .A3(_1065_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit6.Q ),
    .X(_1085_));
 sg13g2_mux4_1 _1255_ (.S0(net1000),
    .A0(net974),
    .A1(net968),
    .A2(net938),
    .A3(net961),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit7.Q ),
    .X(_1086_));
 sg13g2_nor2_1 _1256_ (.A(net1000),
    .B(net955),
    .Y(_1087_));
 sg13g2_a21oi_2 _1257_ (.B1(_1087_),
    .Y(_1088_),
    .A2(_1051_),
    .A1(net1000));
 sg13g2_nand2b_1 _1258_ (.Y(_1089_),
    .B(net1000),
    .A_N(net929));
 sg13g2_o21ai_1 _1259_ (.B1(_1089_),
    .Y(_1090_),
    .A1(net1000),
    .A2(net934));
 sg13g2_o21ai_1 _1260_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit8.Q ),
    .Y(_1091_),
    .A1(_1088_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit7.Q ));
 sg13g2_a21oi_2 _1261_ (.B1(_1091_),
    .Y(_1092_),
    .A2(_1090_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit7.Q ));
 sg13g2_nand2b_1 _1262_ (.Y(_1093_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit9.Q ),
    .A_N(_1092_));
 sg13g2_a21oi_2 _1263_ (.B1(_1093_),
    .Y(_1094_),
    .A2(_1086_),
    .A1(_1015_));
 sg13g2_mux2_1 _1264_ (.A0(net1212),
    .A1(net67),
    .S(net1000),
    .X(_1095_));
 sg13g2_mux2_1 _1265_ (.A0(net94),
    .A1(net106),
    .S(net1000),
    .X(_1096_));
 sg13g2_mux2_1 _1266_ (.A0(net1215),
    .A1(net10),
    .S(net1000),
    .X(_1097_));
 sg13g2_nor2_1 _1267_ (.A(net39),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit6.Q ),
    .Y(_1098_));
 sg13g2_a21oi_1 _1268_ (.A1(_1012_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit6.Q ),
    .Y(_1099_),
    .B1(_1098_));
 sg13g2_mux4_1 _1269_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit7.Q ),
    .A0(_1095_),
    .A1(_1096_),
    .A2(_1099_),
    .A3(_1097_),
    .S1(_1015_),
    .X(_1100_));
 sg13g2_nor2_1 _1270_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit9.Q ),
    .B(_1100_),
    .Y(_1101_));
 sg13g2_nor2_2 _1271_ (.A(_1101_),
    .B(_1094_),
    .Y(\Inst_LUT4AB_switch_matrix.JN2BEG3 ));
 sg13g2_mux4_1 _1272_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit26.Q ),
    .A0(net49),
    .A1(net77),
    .A2(net104),
    .A3(\Inst_LUT4AB_switch_matrix.JN2BEG3 ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit27.Q ),
    .X(_1102_));
 sg13g2_mux4_1 _1273_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit26.Q ),
    .A0(net50),
    .A1(net21),
    .A2(net78),
    .A3(net105),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit27.Q ),
    .X(_1103_));
 sg13g2_inv_1 _1274_ (.Y(_1104_),
    .A(_1103_));
 sg13g2_mux4_1 _1275_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit30.Q ),
    .A0(net957),
    .A1(net951),
    .A2(net935),
    .A3(net931),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit31.Q ),
    .X(_1105_));
 sg13g2_mux4_1 _1276_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit31.Q ),
    .A0(net975),
    .A1(D),
    .A2(net940),
    .A3(net963),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit30.Q ),
    .X(_1106_));
 sg13g2_nand2b_1 _1277_ (.Y(_1107_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit0.Q ),
    .A_N(_1105_));
 sg13g2_o21ai_1 _1278_ (.B1(_1107_),
    .Y(_1108_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit0.Q ),
    .A2(_1106_));
 sg13g2_mux4_1 _1279_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit31.Q ),
    .A0(net37),
    .A1(net2),
    .A2(net53),
    .A3(net8),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit30.Q ),
    .X(_1109_));
 sg13g2_nand2b_1 _1280_ (.Y(_1110_),
    .B(_1109_),
    .A_N(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit0.Q ));
 sg13g2_nand2_1 _1281_ (.Y(_1111_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit30.Q ),
    .B(net65));
 sg13g2_o21ai_1 _1282_ (.B1(_1111_),
    .Y(_1112_),
    .A1(_1014_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit30.Q ));
 sg13g2_nand2b_1 _1283_ (.Y(_1113_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit30.Q ),
    .A_N(net106));
 sg13g2_o21ai_1 _1284_ (.B1(_1113_),
    .Y(_1114_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit30.Q ),
    .A2(net92));
 sg13g2_o21ai_1 _1285_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit0.Q ),
    .Y(_1115_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit31.Q ),
    .A2(_1112_));
 sg13g2_a21oi_1 _1286_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit31.Q ),
    .A2(_1114_),
    .Y(_1116_),
    .B1(_1115_));
 sg13g2_nor2_1 _1287_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit1.Q ),
    .B(_1116_),
    .Y(_1117_));
 sg13g2_a22oi_1 _1288_ (.Y(\Inst_LUT4AB_switch_matrix.JN2BEG1 ),
    .B1(_1110_),
    .B2(_1117_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit1.Q ),
    .A1(_1108_));
 sg13g2_mux4_1 _1289_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit27.Q ),
    .A0(net58),
    .A1(net108),
    .A2(net82),
    .A3(\Inst_LUT4AB_switch_matrix.JN2BEG1 ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit26.Q ),
    .X(_1118_));
 sg13g2_mux4_1 _1290_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit27.Q ),
    .A0(net41),
    .A1(net86),
    .A2(net12),
    .A3(net96),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit26.Q ),
    .X(_1119_));
 sg13g2_mux4_1 _1291_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit3.Q ),
    .A0(_1102_),
    .A1(_1103_),
    .A2(_1119_),
    .A3(_1118_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit4.Q ),
    .X(_1120_));
 sg13g2_mux2_2 _1292_ (.A0(_1120_),
    .A1(net1),
    .S(\Inst_LA_LUT4c_frame_config_dffesr.c_I0mux ),
    .X(_1121_));
 sg13g2_nand2b_1 _1293_ (.Y(_1122_),
    .B(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ),
    .A_N(net982));
 sg13g2_nand2_1 _1294_ (.Y(_1123_),
    .A(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ),
    .B(net982));
 sg13g2_nand3_1 _1295_ (.B(_1122_),
    .C(_1123_),
    .A(_1085_),
    .Y(_1124_));
 sg13g2_nor2b_1 _1296_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit30.Q ),
    .B_N(net956),
    .Y(_1125_));
 sg13g2_a21oi_1 _1297_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit30.Q ),
    .A2(net951),
    .Y(_1126_),
    .B1(_1125_));
 sg13g2_mux2_1 _1298_ (.A0(net935),
    .A1(net929),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit30.Q ),
    .X(_1127_));
 sg13g2_a21oi_1 _1299_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit31.Q ),
    .A2(_1127_),
    .Y(_1128_),
    .B1(_1027_));
 sg13g2_o21ai_1 _1300_ (.B1(_1128_),
    .Y(_1129_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit31.Q ),
    .A2(_1126_));
 sg13g2_mux4_1 _1301_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit31.Q ),
    .A0(net975),
    .A1(net944),
    .A2(net939),
    .A3(net962),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit30.Q ),
    .X(_1130_));
 sg13g2_nor2_1 _1302_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit0.Q ),
    .B(_1130_),
    .Y(_1131_));
 sg13g2_nor2b_1 _1303_ (.A(_1131_),
    .B_N(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit1.Q ),
    .Y(_1132_));
 sg13g2_mux4_1 _1304_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit31.Q ),
    .A0(net57),
    .A1(net24),
    .A2(net1217),
    .A3(net1212),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit30.Q ),
    .X(_1133_));
 sg13g2_inv_1 _1305_ (.Y(_1134_),
    .A(_1133_));
 sg13g2_mux2_1 _1306_ (.A0(net81),
    .A1(net85),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit30.Q ),
    .X(_1135_));
 sg13g2_nand2b_1 _1307_ (.Y(_1136_),
    .B(_1135_),
    .A_N(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit31.Q ));
 sg13g2_mux2_1 _1308_ (.A0(net92),
    .A1(net106),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit30.Q ),
    .X(_1137_));
 sg13g2_a21oi_1 _1309_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit31.Q ),
    .A2(_1137_),
    .Y(_1138_),
    .B1(_1027_));
 sg13g2_a221oi_1 _1310_ (.B2(_1138_),
    .C1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit1.Q ),
    .B1(_1136_),
    .A1(_1027_),
    .Y(_1139_),
    .A2(_1134_));
 sg13g2_a21o_1 _1311_ (.A2(_1132_),
    .A1(_1129_),
    .B1(_1139_),
    .X(\Inst_LUT4AB_switch_matrix.JS2BEG1 ));
 sg13g2_mux4_1 _1312_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit30.Q ),
    .A0(net52),
    .A1(net1210),
    .A2(net107),
    .A3(\Inst_LUT4AB_switch_matrix.JS2BEG1 ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit31.Q ),
    .X(_1140_));
 sg13g2_mux4_1 _1313_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit31.Q ),
    .A0(net39),
    .A1(net67),
    .A2(net22),
    .A3(net94),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit30.Q ),
    .X(_1141_));
 sg13g2_mux4_1 _1314_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit6.Q ),
    .A0(net974),
    .A1(net968),
    .A2(net938),
    .A3(net961),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit7.Q ),
    .X(_1142_));
 sg13g2_inv_1 _1315_ (.Y(_1143_),
    .A(_1142_));
 sg13g2_mux2_1 _1316_ (.A0(net955),
    .A1(net950),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit6.Q ),
    .X(_1144_));
 sg13g2_nand2b_1 _1317_ (.Y(_1145_),
    .B(_1144_),
    .A_N(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit7.Q ));
 sg13g2_mux2_1 _1318_ (.A0(net934),
    .A1(net931),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit6.Q ),
    .X(_1146_));
 sg13g2_a21oi_1 _1319_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit7.Q ),
    .A2(_1146_),
    .Y(_1147_),
    .B1(_1024_));
 sg13g2_a221oi_1 _1320_ (.B2(_1147_),
    .C1(_1025_),
    .B1(_1145_),
    .A1(_1024_),
    .Y(_1148_),
    .A2(_1143_));
 sg13g2_nor2b_1 _1321_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit6.Q ),
    .B_N(net67),
    .Y(_1149_));
 sg13g2_a21oi_1 _1322_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit6.Q ),
    .A2(net79),
    .Y(_1150_),
    .B1(_1149_));
 sg13g2_mux2_1 _1323_ (.A0(net94),
    .A1(net110),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit6.Q ),
    .X(_1151_));
 sg13g2_a21oi_1 _1324_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit7.Q ),
    .A2(_1151_),
    .Y(_1152_),
    .B1(_1024_));
 sg13g2_o21ai_1 _1325_ (.B1(_1152_),
    .Y(_1153_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit7.Q ),
    .A2(_1150_));
 sg13g2_mux4_1 _1326_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit6.Q ),
    .A0(net39),
    .A1(net1215),
    .A2(net10),
    .A3(net1212),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit7.Q ),
    .X(_1154_));
 sg13g2_nor2_1 _1327_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit8.Q ),
    .B(_1154_),
    .Y(_1155_));
 sg13g2_nor2_1 _1328_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit9.Q ),
    .B(_1155_),
    .Y(_1156_));
 sg13g2_a21o_2 _1329_ (.A2(_1156_),
    .A1(_1153_),
    .B1(_1148_),
    .X(\Inst_LUT4AB_switch_matrix.JS2BEG3 ));
 sg13g2_mux4_1 _1330_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit30.Q ),
    .A0(net47),
    .A1(net18),
    .A2(net102),
    .A3(\Inst_LUT4AB_switch_matrix.JS2BEG3 ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit31.Q ),
    .X(_1157_));
 sg13g2_inv_1 _1331_ (.Y(_1158_),
    .A(_1157_));
 sg13g2_mux4_1 _1332_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit30.Q ),
    .A0(net48),
    .A1(net19),
    .A2(net76),
    .A3(net103),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit31.Q ),
    .X(_1159_));
 sg13g2_mux4_1 _1333_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit7.Q ),
    .A0(_1157_),
    .A1(_1159_),
    .A2(_1141_),
    .A3(_1140_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit8.Q ),
    .X(_1160_));
 sg13g2_mux2_1 _1334_ (.A0(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ),
    .A1(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ),
    .S(net982),
    .X(_1161_));
 sg13g2_nor2_1 _1335_ (.A(_1085_),
    .B(_1161_),
    .Y(_1162_));
 sg13g2_nor2_1 _1336_ (.A(_1160_),
    .B(_1162_),
    .Y(_0008_));
 sg13g2_mux4_1 _1337_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit30.Q ),
    .A0(net955),
    .A1(net950),
    .A2(net934),
    .A3(net928),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit31.Q ),
    .X(_0009_));
 sg13g2_mux4_1 _1338_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit31.Q ),
    .A0(net974),
    .A1(net944),
    .A2(net938),
    .A3(net962),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit30.Q ),
    .X(_0010_));
 sg13g2_nand2b_1 _1339_ (.Y(_0011_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit0.Q ),
    .A_N(_0009_));
 sg13g2_o21ai_1 _1340_ (.B1(_0011_),
    .Y(_0012_),
    .A1(_0010_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit0.Q ));
 sg13g2_mux4_1 _1341_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit31.Q ),
    .A0(net1010),
    .A1(net8),
    .A2(net37),
    .A3(net1212),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit30.Q ),
    .X(_0013_));
 sg13g2_nor2b_1 _1342_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit0.Q ),
    .B_N(_0013_),
    .Y(_0014_));
 sg13g2_mux2_1 _1343_ (.A0(net65),
    .A1(net81),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit30.Q ),
    .X(_0015_));
 sg13g2_nand2b_1 _1344_ (.Y(_0016_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit30.Q ),
    .A_N(net106));
 sg13g2_o21ai_1 _1345_ (.B1(_0016_),
    .Y(_0017_),
    .A1(net92),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit30.Q ));
 sg13g2_o21ai_1 _1346_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit0.Q ),
    .Y(_0018_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit31.Q ),
    .A2(_0015_));
 sg13g2_a21oi_1 _1347_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit31.Q ),
    .A2(_0017_),
    .Y(_0019_),
    .B1(_0018_));
 sg13g2_nor3_1 _1348_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit1.Q ),
    .B(_0014_),
    .C(_0019_),
    .Y(_0020_));
 sg13g2_a21o_2 _1349_ (.A2(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit1.Q ),
    .A1(_0012_),
    .B1(_0020_),
    .X(_0021_));
 sg13g2_inv_1 _1350_ (.Y(\Inst_LUT4AB_switch_matrix.JW2BEG1 ),
    .A(_0021_));
 sg13g2_mux4_1 _1351_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit0.Q ),
    .A0(_1012_),
    .A1(_1014_),
    .A2(_1022_),
    .A3(_0021_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit1.Q ),
    .X(_0022_));
 sg13g2_mux4_1 _1352_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit1.Q ),
    .A0(net35),
    .A1(net63),
    .A2(net6),
    .A3(net111),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit0.Q ),
    .X(_0023_));
 sg13g2_mux4_1 _1353_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit6.Q ),
    .A0(net974),
    .A1(net968),
    .A2(net938),
    .A3(net961),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit7.Q ),
    .X(_0024_));
 sg13g2_mux4_1 _1354_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit6.Q ),
    .A0(net955),
    .A1(net950),
    .A2(net934),
    .A3(net930),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit7.Q ),
    .X(_0025_));
 sg13g2_nand2b_1 _1355_ (.Y(_0026_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit8.Q ),
    .A_N(_0025_));
 sg13g2_o21ai_1 _1356_ (.B1(_0026_),
    .Y(_0027_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit8.Q ),
    .A2(_0024_));
 sg13g2_mux4_1 _1357_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit7.Q ),
    .A0(net1008),
    .A1(net10),
    .A2(net39),
    .A3(net1212),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit6.Q ),
    .X(_0028_));
 sg13g2_nor2b_1 _1358_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit8.Q ),
    .B_N(_0028_),
    .Y(_0029_));
 sg13g2_nor2_1 _1359_ (.A(net67),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit6.Q ),
    .Y(_0030_));
 sg13g2_a21oi_1 _1360_ (.A1(_1022_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit6.Q ),
    .Y(_0031_),
    .B1(_0030_));
 sg13g2_nand2_1 _1361_ (.Y(_0032_),
    .A(_1023_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit6.Q ));
 sg13g2_o21ai_1 _1362_ (.B1(_0032_),
    .Y(_0033_),
    .A1(net94),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit6.Q ));
 sg13g2_o21ai_1 _1363_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit8.Q ),
    .Y(_0034_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit7.Q ),
    .A2(_0031_));
 sg13g2_a21oi_1 _1364_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit7.Q ),
    .A2(_0033_),
    .Y(_0035_),
    .B1(_0034_));
 sg13g2_nor3_1 _1365_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit9.Q ),
    .B(_0029_),
    .C(_0035_),
    .Y(_0036_));
 sg13g2_a21o_2 _1366_ (.A2(_0027_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit9.Q ),
    .B1(_0036_),
    .X(_0037_));
 sg13g2_inv_1 _1367_ (.Y(\Inst_LUT4AB_switch_matrix.JW2BEG3 ),
    .A(_0037_));
 sg13g2_o21ai_1 _1368_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit1.Q ),
    .Y(_0038_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit0.Q ),
    .A2(net71));
 sg13g2_a21oi_1 _1369_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit0.Q ),
    .A2(_0037_),
    .Y(_0039_),
    .B1(_0038_));
 sg13g2_nor2b_1 _1370_ (.A(net14),
    .B_N(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit0.Q ),
    .Y(_0040_));
 sg13g2_nor2_1 _1371_ (.A(net43),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit0.Q ),
    .Y(_0041_));
 sg13g2_nor3_1 _1372_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit1.Q ),
    .B(_0040_),
    .C(_0041_),
    .Y(_0042_));
 sg13g2_nor2_1 _1373_ (.A(_0039_),
    .B(_0042_),
    .Y(_0043_));
 sg13g2_mux2_1 _1374_ (.A0(net44),
    .A1(net15),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit0.Q ),
    .X(_0044_));
 sg13g2_nand2b_1 _1375_ (.Y(_0045_),
    .B(net72),
    .A_N(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit0.Q ));
 sg13g2_nand2_1 _1376_ (.Y(_0046_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit0.Q ),
    .B(net99));
 sg13g2_nand3_1 _1377_ (.B(_0045_),
    .C(_0046_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit1.Q ),
    .Y(_0047_));
 sg13g2_o21ai_1 _1378_ (.B1(_0047_),
    .Y(_0048_),
    .A1(_0044_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit1.Q ));
 sg13g2_nand2_2 _1379_ (.Y(_0049_),
    .A(_0048_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit9.Q ));
 sg13g2_a21oi_1 _1380_ (.A1(_1029_),
    .A2(_0043_),
    .Y(_0050_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit10.Q ));
 sg13g2_o21ai_1 _1381_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit10.Q ),
    .Y(_0051_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit9.Q ),
    .A2(_0023_));
 sg13g2_a21oi_1 _1382_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit9.Q ),
    .A2(_0022_),
    .Y(_0052_),
    .B1(_0051_));
 sg13g2_a21oi_1 _1383_ (.A1(_0049_),
    .A2(_0050_),
    .Y(_0053_),
    .B1(_0052_));
 sg13g2_mux2_1 _1384_ (.A0(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ),
    .A1(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ),
    .S(net982),
    .X(_0054_));
 sg13g2_mux2_1 _1385_ (.A0(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ),
    .A1(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ),
    .S(net982),
    .X(_0055_));
 sg13g2_mux2_1 _1386_ (.A0(_0055_),
    .A1(_0054_),
    .S(_1085_),
    .X(_0056_));
 sg13g2_a221oi_1 _1387_ (.B2(_1160_),
    .C1(_0053_),
    .B1(_0056_),
    .A1(_1124_),
    .Y(_0057_),
    .A2(_0008_));
 sg13g2_mux2_1 _1388_ (.A0(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ),
    .A1(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ),
    .S(_1121_),
    .X(_0058_));
 sg13g2_mux2_1 _1389_ (.A0(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ),
    .A1(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ),
    .S(net982),
    .X(_0059_));
 sg13g2_mux2_1 _1390_ (.A0(_0059_),
    .A1(_0058_),
    .S(_1085_),
    .X(_0060_));
 sg13g2_nand2b_1 _1391_ (.Y(_0061_),
    .B(_0060_),
    .A_N(_1160_));
 sg13g2_nand2b_1 _1392_ (.Y(_0062_),
    .B(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ),
    .A_N(_1121_));
 sg13g2_a21oi_1 _1393_ (.A1(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ),
    .A2(_1121_),
    .Y(_0063_),
    .B1(_1085_));
 sg13g2_nand2_1 _1394_ (.Y(_0064_),
    .A(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ),
    .B(net982));
 sg13g2_nand2b_1 _1395_ (.Y(_0065_),
    .B(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ),
    .A_N(net982));
 sg13g2_and2_1 _1396_ (.A(_1085_),
    .B(_0065_),
    .X(_0066_));
 sg13g2_a22oi_1 _1397_ (.Y(_0067_),
    .B1(_0064_),
    .B2(_0066_),
    .A2(_0063_),
    .A1(_0062_));
 sg13g2_a221oi_1 _1398_ (.B2(_1160_),
    .C1(_0052_),
    .B1(_0067_),
    .A1(_0050_),
    .Y(_0068_),
    .A2(_0049_));
 sg13g2_a21oi_2 _1399_ (.B1(_0057_),
    .Y(_0069_),
    .A2(_0061_),
    .A1(_0068_));
 sg13g2_mux2_2 _1400_ (.A0(_0069_),
    .A1(\Inst_LA_LUT4c_frame_config_dffesr.LUT_flop ),
    .S(\Inst_LA_LUT4c_frame_config_dffesr.c_out_mux ),
    .X(A));
 sg13g2_o21ai_1 _1401_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit20.Q ),
    .Y(_0070_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit19.Q ),
    .A2(_0023_));
 sg13g2_a21o_1 _1402_ (.A2(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit19.Q ),
    .A1(_0022_),
    .B1(_0070_),
    .X(_0071_));
 sg13g2_mux2_1 _1403_ (.A0(_0043_),
    .A1(_0048_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit19.Q ),
    .X(_0072_));
 sg13g2_o21ai_1 _1404_ (.B1(_0071_),
    .Y(_0073_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit20.Q ),
    .A2(_0072_));
 sg13g2_mux4_1 _1405_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit15.Q ),
    .A0(_1083_),
    .A1(_1084_),
    .A2(_1066_),
    .A3(_1065_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit16.Q ),
    .X(_0074_));
 sg13g2_mux4_1 _1406_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit17.Q ),
    .A0(_1157_),
    .A1(_1159_),
    .A2(_1141_),
    .A3(_1140_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit18.Q ),
    .X(_0075_));
 sg13g2_nand2b_1 _1407_ (.Y(_0076_),
    .B(_0075_),
    .A_N(_0074_));
 sg13g2_o21ai_1 _1408_ (.B1(_0073_),
    .Y(_0077_),
    .A1(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ),
    .A2(_0076_));
 sg13g2_nor2b_1 _1409_ (.A(_0075_),
    .B_N(_0074_),
    .Y(_0078_));
 sg13g2_nor2b_1 _1410_ (.A(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ),
    .B_N(_0078_),
    .Y(_0079_));
 sg13g2_and2_1 _1411_ (.A(_0074_),
    .B(_0075_),
    .X(_0080_));
 sg13g2_nand2_1 _1412_ (.Y(_0081_),
    .A(_0074_),
    .B(_0075_));
 sg13g2_nor2_1 _1413_ (.A(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ),
    .B(_0081_),
    .Y(_0082_));
 sg13g2_or2_1 _1414_ (.X(_0083_),
    .B(_0075_),
    .A(_0074_));
 sg13g2_nor2_1 _1415_ (.A(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ),
    .B(_0083_),
    .Y(_0084_));
 sg13g2_or4_1 _1416_ (.A(_0084_),
    .B(_0079_),
    .C(_0082_),
    .D(_0077_),
    .X(_0085_));
 sg13g2_mux4_1 _1417_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit13.Q ),
    .A0(_1102_),
    .A1(_1103_),
    .A2(_1119_),
    .A3(_1118_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit14.Q ),
    .X(_0086_));
 sg13g2_nand2_1 _1418_ (.Y(_0087_),
    .A(net1),
    .B(_1160_));
 sg13g2_o21ai_1 _1419_ (.B1(_1085_),
    .Y(_0088_),
    .A1(net1),
    .A2(_1160_));
 sg13g2_nand2_2 _1420_ (.Y(_0089_),
    .A(_0088_),
    .B(_0087_));
 sg13g2_nor2b_1 _1421_ (.A(\Inst_LB_LUT4c_frame_config_dffesr.c_I0mux ),
    .B_N(_0086_),
    .Y(_0090_));
 sg13g2_a21oi_1 _1422_ (.A1(\Inst_LB_LUT4c_frame_config_dffesr.c_I0mux ),
    .A2(_0089_),
    .Y(_0091_),
    .B1(_0090_));
 sg13g2_nor2b_1 _1423_ (.A(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ),
    .B_N(_0078_),
    .Y(_0092_));
 sg13g2_nor2_1 _1424_ (.A(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ),
    .B(_0081_),
    .Y(_0093_));
 sg13g2_or2_1 _1425_ (.X(_0094_),
    .B(_0076_),
    .A(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ));
 sg13g2_o21ai_1 _1426_ (.B1(_0094_),
    .Y(_0095_),
    .A1(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ),
    .A2(_0083_));
 sg13g2_or4_1 _1427_ (.A(_0073_),
    .B(_0092_),
    .C(_0093_),
    .D(_0095_),
    .X(_0096_));
 sg13g2_and2_1 _1428_ (.A(_0091_),
    .B(_0096_),
    .X(_0097_));
 sg13g2_o21ai_1 _1429_ (.B1(_0073_),
    .Y(_0098_),
    .A1(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ),
    .A2(_0081_));
 sg13g2_nor2_1 _1430_ (.A(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ),
    .B(_0083_),
    .Y(_0099_));
 sg13g2_nand2b_1 _1431_ (.Y(_0100_),
    .B(_0078_),
    .A_N(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ));
 sg13g2_o21ai_1 _1432_ (.B1(_0100_),
    .Y(_0101_),
    .A1(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ),
    .A2(_0076_));
 sg13g2_nor3_1 _1433_ (.A(_0098_),
    .B(_0099_),
    .C(_0101_),
    .Y(_0102_));
 sg13g2_nor2_1 _1434_ (.A(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ),
    .B(_0076_),
    .Y(_0103_));
 sg13g2_nor2_1 _1435_ (.A(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ),
    .B(_0081_),
    .Y(_0104_));
 sg13g2_nand2b_1 _1436_ (.Y(_0105_),
    .B(_0078_),
    .A_N(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ));
 sg13g2_o21ai_1 _1437_ (.B1(_0105_),
    .Y(_0106_),
    .A1(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ),
    .A2(_0083_));
 sg13g2_nor4_1 _1438_ (.A(_0073_),
    .B(_0103_),
    .C(_0104_),
    .D(_0106_),
    .Y(_0107_));
 sg13g2_nor3_1 _1439_ (.A(_0091_),
    .B(_0102_),
    .C(_0107_),
    .Y(_0108_));
 sg13g2_a21oi_2 _1440_ (.B1(_0108_),
    .Y(_0109_),
    .A2(_0085_),
    .A1(_0097_));
 sg13g2_mux2_1 _1441_ (.A0(_0109_),
    .A1(\Inst_LB_LUT4c_frame_config_dffesr.LUT_flop ),
    .S(\Inst_LB_LUT4c_frame_config_dffesr.c_out_mux ),
    .X(B));
 sg13g2_nand2b_1 _1442_ (.Y(_0110_),
    .B(net993),
    .A_N(net931));
 sg13g2_o21ai_1 _1443_ (.B1(_0110_),
    .Y(_0111_),
    .A1(net993),
    .A2(net935));
 sg13g2_mux2_1 _1444_ (.A0(net957),
    .A1(net952),
    .S(net993),
    .X(_0112_));
 sg13g2_o21ai_1 _1445_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit4.Q ),
    .Y(_0113_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit3.Q ),
    .A2(_0112_));
 sg13g2_a21oi_1 _1446_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit3.Q ),
    .A2(_0111_),
    .Y(_0114_),
    .B1(_0113_));
 sg13g2_nand2b_1 _1447_ (.Y(_0115_),
    .B(net993),
    .A_N(net964));
 sg13g2_o21ai_1 _1448_ (.B1(_0115_),
    .Y(_0116_),
    .A1(net993),
    .A2(net945));
 sg13g2_mux2_1 _1449_ (.A0(net975),
    .A1(net970),
    .S(net993),
    .X(_0117_));
 sg13g2_o21ai_1 _1450_ (.B1(_1032_),
    .Y(_0118_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit3.Q ),
    .A2(_0117_));
 sg13g2_a21oi_1 _1451_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit3.Q ),
    .A2(_0116_),
    .Y(_0119_),
    .B1(_0118_));
 sg13g2_nor3_1 _1452_ (.A(_1033_),
    .B(_0114_),
    .C(_0119_),
    .Y(_0120_));
 sg13g2_mux4_1 _1453_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit3.Q ),
    .A0(net1009),
    .A1(net54),
    .A2(net38),
    .A3(net9),
    .S1(net993),
    .X(_0121_));
 sg13g2_nand2_1 _1454_ (.Y(_0122_),
    .A(_1032_),
    .B(_0121_));
 sg13g2_nand2b_1 _1455_ (.Y(_0123_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit2.Q ),
    .A_N(net107));
 sg13g2_o21ai_1 _1456_ (.B1(_0123_),
    .Y(_0124_),
    .A1(net93),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit2.Q ));
 sg13g2_mux2_1 _1457_ (.A0(net1210),
    .A1(net66),
    .S(net993),
    .X(_0125_));
 sg13g2_o21ai_1 _1458_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit4.Q ),
    .Y(_0126_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit3.Q ),
    .A2(_0125_));
 sg13g2_a21oi_1 _1459_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit3.Q ),
    .A2(_0124_),
    .Y(_0127_),
    .B1(_0126_));
 sg13g2_nor2_1 _1460_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit5.Q ),
    .B(_0127_),
    .Y(_0128_));
 sg13g2_a21oi_1 _1461_ (.A1(_0122_),
    .A2(_0128_),
    .Y(\Inst_LUT4AB_switch_matrix.E2BEG2 ),
    .B1(_0120_));
 sg13g2_mux4_1 _1462_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit4.Q ),
    .A0(net53),
    .A1(net8),
    .A2(net97),
    .A3(\Inst_LUT4AB_switch_matrix.E2BEG2 ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit5.Q ),
    .X(_0129_));
 sg13g2_mux4_1 _1463_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit4.Q ),
    .A0(net37),
    .A1(net8),
    .A2(net65),
    .A3(net110),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit5.Q ),
    .X(_0130_));
 sg13g2_mux4_1 _1464_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit10.Q ),
    .A0(net976),
    .A1(net972),
    .A2(net942),
    .A3(net947),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit11.Q ),
    .X(_0131_));
 sg13g2_nand2b_1 _1465_ (.Y(_0132_),
    .B(_0131_),
    .A_N(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit12.Q ));
 sg13g2_mux2_1 _1466_ (.A0(net959),
    .A1(net954),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit10.Q ),
    .X(_0133_));
 sg13g2_nand2b_1 _1467_ (.Y(_0134_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit10.Q ),
    .A_N(\Inst_LUT4AB_switch_matrix.M_EF ));
 sg13g2_o21ai_1 _1468_ (.B1(_0134_),
    .Y(_0135_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit10.Q ),
    .A2(net936));
 sg13g2_o21ai_1 _1469_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit12.Q ),
    .Y(_0136_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit11.Q ),
    .A2(_0133_));
 sg13g2_a21oi_2 _1470_ (.B1(_0136_),
    .Y(_0137_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit11.Q ),
    .A1(_0135_));
 sg13g2_nor2b_1 _1471_ (.A(_0137_),
    .B_N(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit13.Q ),
    .Y(_0138_));
 sg13g2_mux4_1 _1472_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit10.Q ),
    .A0(net32),
    .A1(net40),
    .A2(net1216),
    .A3(net11),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit11.Q ),
    .X(_0139_));
 sg13g2_nand2b_1 _1473_ (.Y(_0140_),
    .B(_0139_),
    .A_N(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit12.Q ));
 sg13g2_nand2b_1 _1474_ (.Y(_0141_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit10.Q ),
    .A_N(net1006));
 sg13g2_o21ai_1 _1475_ (.B1(_0141_),
    .Y(_0142_),
    .A1(net68),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit10.Q ));
 sg13g2_mux2_1 _1476_ (.A0(net60),
    .A1(net62),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit10.Q ),
    .X(_0143_));
 sg13g2_o21ai_1 _1477_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit12.Q ),
    .Y(_0144_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit11.Q ),
    .A2(_0143_));
 sg13g2_a21oi_1 _1478_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit11.Q ),
    .A2(_0142_),
    .Y(_0145_),
    .B1(_0144_));
 sg13g2_nor2_1 _1479_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit13.Q ),
    .B(_0145_),
    .Y(_0146_));
 sg13g2_a22oi_1 _1480_ (.Y(\Inst_LUT4AB_switch_matrix.E2BEG4 ),
    .B1(_0140_),
    .B2(_0146_),
    .A2(_0132_),
    .A1(_0138_));
 sg13g2_mux4_1 _1481_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit5.Q ),
    .A0(net45),
    .A1(net100),
    .A2(net16),
    .A3(\Inst_LUT4AB_switch_matrix.E2BEG4 ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit4.Q ),
    .X(_0147_));
 sg13g2_mux4_1 _1482_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit4.Q ),
    .A0(net46),
    .A1(net17),
    .A2(net74),
    .A3(net101),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit5.Q ),
    .X(_0148_));
 sg13g2_mux4_1 _1483_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit3.Q ),
    .A0(_0147_),
    .A1(_0148_),
    .A2(_0130_),
    .A3(_0129_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit4.Q ),
    .X(_0149_));
 sg13g2_nand2b_1 _1484_ (.Y(_0150_),
    .B(net990),
    .A_N(net966));
 sg13g2_o21ai_1 _1485_ (.B1(_0150_),
    .Y(_0151_),
    .A1(net990),
    .A2(net947));
 sg13g2_mux2_1 _1486_ (.A0(net978),
    .A1(net972),
    .S(net990),
    .X(_0152_));
 sg13g2_o21ai_1 _1487_ (.B1(_1037_),
    .Y(_0153_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit3.Q ),
    .A2(_0152_));
 sg13g2_a21oi_1 _1488_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit3.Q ),
    .A2(_0151_),
    .Y(_0154_),
    .B1(_0153_));
 sg13g2_nor2_1 _1489_ (.A(net990),
    .B(net959),
    .Y(_0155_));
 sg13g2_a21oi_1 _1490_ (.A1(net990),
    .A2(_1051_),
    .Y(_0156_),
    .B1(_0155_));
 sg13g2_nand2b_1 _1491_ (.Y(_0157_),
    .B(net990),
    .A_N(\Inst_LUT4AB_switch_matrix.M_AB ));
 sg13g2_o21ai_1 _1492_ (.B1(_0157_),
    .Y(_0158_),
    .A1(net990),
    .A2(net937));
 sg13g2_a21oi_2 _1493_ (.B1(_1037_),
    .Y(_0159_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit3.Q ),
    .A1(_0158_));
 sg13g2_o21ai_1 _1494_ (.B1(_0159_),
    .Y(_0160_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit3.Q ),
    .A2(_0156_));
 sg13g2_nor2_1 _1495_ (.A(_1038_),
    .B(_0154_),
    .Y(_0161_));
 sg13g2_mux4_1 _1496_ (.S0(net990),
    .A0(net58),
    .A1(net1216),
    .A2(net9),
    .A3(net1211),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit3.Q ),
    .X(_0162_));
 sg13g2_nand2b_1 _1497_ (.Y(_0163_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit2.Q ),
    .A_N(net107));
 sg13g2_o21ai_1 _1498_ (.B1(_0163_),
    .Y(_0164_),
    .A1(net93),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit2.Q ));
 sg13g2_mux2_1 _1499_ (.A0(net66),
    .A1(net82),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit2.Q ),
    .X(_0165_));
 sg13g2_o21ai_1 _1500_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit4.Q ),
    .Y(_0166_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit3.Q ),
    .A2(_0165_));
 sg13g2_a21oi_1 _1501_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit3.Q ),
    .A2(_0164_),
    .Y(_0167_),
    .B1(_0166_));
 sg13g2_a21oi_1 _1502_ (.A1(_1037_),
    .A2(_0162_),
    .Y(_0168_),
    .B1(_0167_));
 sg13g2_a22oi_1 _1503_ (.Y(\Inst_LUT4AB_switch_matrix.JS2BEG2 ),
    .B1(_0168_),
    .B2(_1038_),
    .A2(_0160_),
    .A1(_0161_));
 sg13g2_mux4_1 _1504_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit6.Q ),
    .A0(net56),
    .A1(net23),
    .A2(net80),
    .A3(\Inst_LUT4AB_switch_matrix.JS2BEG2 ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit7.Q ),
    .X(_0169_));
 sg13g2_mux4_1 _1505_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit6.Q ),
    .A0(net39),
    .A1(net10),
    .A2(net85),
    .A3(net94),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit7.Q ),
    .X(_0170_));
 sg13g2_inv_1 _1506_ (.Y(_0171_),
    .A(_0170_));
 sg13g2_nand2b_1 _1507_ (.Y(_0172_),
    .B(net989),
    .A_N(net946));
 sg13g2_o21ai_1 _1508_ (.B1(_0172_),
    .Y(_0173_),
    .A1(net989),
    .A2(net941));
 sg13g2_mux2_1 _1509_ (.A0(net976),
    .A1(net971),
    .S(net989),
    .X(_0174_));
 sg13g2_a21oi_2 _1510_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit12.Q ),
    .Y(_0175_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit11.Q ),
    .A1(_0173_));
 sg13g2_o21ai_1 _1511_ (.B1(_0175_),
    .Y(_0176_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit11.Q ),
    .A2(_0174_));
 sg13g2_mux2_1 _1512_ (.A0(net958),
    .A1(net954),
    .S(net988),
    .X(_0177_));
 sg13g2_nand2b_1 _1513_ (.Y(_0178_),
    .B(net989),
    .A_N(net928));
 sg13g2_o21ai_1 _1514_ (.B1(_0178_),
    .Y(_0179_),
    .A1(net989),
    .A2(net936));
 sg13g2_o21ai_1 _1515_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit12.Q ),
    .Y(_0180_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit11.Q ),
    .A2(_0177_));
 sg13g2_a21oi_1 _1516_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit11.Q ),
    .A2(_0179_),
    .Y(_0181_),
    .B1(_0180_));
 sg13g2_nor2_1 _1517_ (.A(_1035_),
    .B(_0181_),
    .Y(_0182_));
 sg13g2_nand2b_1 _1518_ (.Y(_0183_),
    .B(net988),
    .A_N(net68));
 sg13g2_o21ai_1 _1519_ (.B1(_0183_),
    .Y(_0184_),
    .A1(net60),
    .A2(net988));
 sg13g2_nand2b_1 _1520_ (.Y(_0185_),
    .B(net988),
    .A_N(net89));
 sg13g2_o21ai_1 _1521_ (.B1(_0185_),
    .Y(_0186_),
    .A1(net1006),
    .A2(net989));
 sg13g2_nand2b_1 _1522_ (.Y(_0187_),
    .B(net988),
    .A_N(net11));
 sg13g2_o21ai_1 _1523_ (.B1(_0187_),
    .Y(_0188_),
    .A1(net1216),
    .A2(net988));
 sg13g2_nand2b_1 _1524_ (.Y(_0189_),
    .B(net988),
    .A_N(net40));
 sg13g2_o21ai_1 _1525_ (.B1(_0189_),
    .Y(_0190_),
    .A1(net1009),
    .A2(net988));
 sg13g2_mux4_1 _1526_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit11.Q ),
    .A0(_0190_),
    .A1(_0188_),
    .A2(_0184_),
    .A3(_0186_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit12.Q ),
    .X(_0191_));
 sg13g2_a22oi_1 _1527_ (.Y(\Inst_LUT4AB_switch_matrix.JS2BEG4 ),
    .B1(_0191_),
    .B2(_1035_),
    .A2(_0176_),
    .A1(_0182_));
 sg13g2_o21ai_1 _1528_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit7.Q ),
    .Y(_0192_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit6.Q ),
    .A2(_1034_));
 sg13g2_a21o_1 _1529_ (.A2(net380),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit6.Q ),
    .B1(_0192_),
    .X(_0193_));
 sg13g2_nand2_1 _1530_ (.Y(_0194_),
    .A(net18),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit6.Q ));
 sg13g2_o21ai_1 _1531_ (.B1(_0194_),
    .Y(_0195_),
    .A1(_1021_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit6.Q ));
 sg13g2_o21ai_1 _1532_ (.B1(_0193_),
    .Y(_0196_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit7.Q ),
    .A2(_0195_));
 sg13g2_mux4_1 _1533_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit6.Q ),
    .A0(net47),
    .A1(net18),
    .A2(net75),
    .A3(net380),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit7.Q ),
    .X(_0197_));
 sg13g2_mux4_1 _1534_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit6.Q ),
    .A0(net48),
    .A1(net19),
    .A2(net76),
    .A3(net103),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit7.Q ),
    .X(_0198_));
 sg13g2_mux4_1 _1535_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit5.Q ),
    .A0(_0197_),
    .A1(_0198_),
    .A2(_0170_),
    .A3(_0169_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit6.Q ),
    .X(_0199_));
 sg13g2_nor2_1 _1536_ (.A(_0149_),
    .B(_0199_),
    .Y(_0200_));
 sg13g2_nand2_1 _1537_ (.Y(_0201_),
    .A(_0149_),
    .B(_0199_));
 sg13g2_mux4_1 _1538_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit25.Q ),
    .A0(_0147_),
    .A1(_0148_),
    .A2(_0130_),
    .A3(_0129_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit26.Q ),
    .X(_0202_));
 sg13g2_mux4_1 _1539_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit27.Q ),
    .A0(_0197_),
    .A1(_0198_),
    .A2(_0170_),
    .A3(_0169_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit28.Q ),
    .X(_0203_));
 sg13g2_or2_1 _1540_ (.X(_0204_),
    .B(_0203_),
    .A(_0202_));
 sg13g2_nand2_1 _1541_ (.Y(_0205_),
    .A(_0202_),
    .B(_0203_));
 sg13g2_inv_1 _1542_ (.Y(_0206_),
    .A(_0205_));
 sg13g2_a21o_1 _1543_ (.A2(_0083_),
    .A1(_0089_),
    .B1(_0080_),
    .X(_0207_));
 sg13g2_a21oi_2 _1544_ (.B1(_0206_),
    .Y(_0208_),
    .A2(_0204_),
    .A1(_0207_));
 sg13g2_o21ai_1 _1545_ (.B1(_0201_),
    .Y(_0209_),
    .A1(_0208_),
    .A2(_0200_));
 sg13g2_o21ai_1 _1546_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit15.Q ),
    .Y(_0210_),
    .A1(net998),
    .A2(net933));
 sg13g2_a21oi_1 _1547_ (.A1(net997),
    .A2(\Inst_LUT4AB_switch_matrix.M_AD ),
    .Y(_0211_),
    .B1(_0210_));
 sg13g2_nor2_1 _1548_ (.A(net997),
    .B(net965),
    .Y(_0212_));
 sg13g2_a21oi_1 _1549_ (.A1(net997),
    .A2(_1051_),
    .Y(_0213_),
    .B1(_0212_));
 sg13g2_o21ai_1 _1550_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit16.Q ),
    .Y(_0214_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit15.Q ),
    .A2(_0213_));
 sg13g2_nor2_1 _1551_ (.A(_0211_),
    .B(_0214_),
    .Y(_0215_));
 sg13g2_nand2b_1 _1552_ (.Y(_0216_),
    .B(net997),
    .A_N(net946));
 sg13g2_o21ai_1 _1553_ (.B1(_0216_),
    .Y(_0217_),
    .A1(net997),
    .A2(net941));
 sg13g2_mux2_1 _1554_ (.A0(net976),
    .A1(net971),
    .S(net998),
    .X(_0218_));
 sg13g2_a21oi_2 _1555_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit16.Q ),
    .Y(_0219_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit15.Q ),
    .A1(_0217_));
 sg13g2_o21ai_1 _1556_ (.B1(_0219_),
    .Y(_0220_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit15.Q ),
    .A2(_0218_));
 sg13g2_nand2_2 _1557_ (.Y(_0221_),
    .A(_0220_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit17.Q ));
 sg13g2_mux4_1 _1558_ (.S0(net998),
    .A0(net33),
    .A1(net41),
    .A2(net4),
    .A3(net12),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit15.Q ),
    .X(_0222_));
 sg13g2_nor2b_1 _1559_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit16.Q ),
    .B_N(_0222_),
    .Y(_0223_));
 sg13g2_nand2b_1 _1560_ (.Y(_0224_),
    .B(net997),
    .A_N(net1004));
 sg13g2_o21ai_1 _1561_ (.B1(_0224_),
    .Y(_0225_),
    .A1(net997),
    .A2(net87));
 sg13g2_mux2_1 _1562_ (.A0(net61),
    .A1(net69),
    .S(net997),
    .X(_0226_));
 sg13g2_o21ai_1 _1563_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit16.Q ),
    .Y(_0227_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit15.Q ),
    .A2(_0226_));
 sg13g2_a21oi_1 _1564_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit15.Q ),
    .A2(_0225_),
    .Y(_0228_),
    .B1(_0227_));
 sg13g2_or3_1 _1565_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit17.Q ),
    .B(_0223_),
    .C(_0228_),
    .X(_0229_));
 sg13g2_o21ai_1 _1566_ (.B1(_0229_),
    .Y(_0230_),
    .A1(_0221_),
    .A2(_0215_));
 sg13g2_inv_2 _1567_ (.Y(\Inst_LUT4AB_switch_matrix.JN2BEG5 ),
    .A(_0230_));
 sg13g2_o21ai_1 _1568_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit11.Q ),
    .Y(_0231_),
    .A1(net104),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit10.Q ));
 sg13g2_a21oi_1 _1569_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit10.Q ),
    .A2(_0230_),
    .Y(_0232_),
    .B1(_0231_));
 sg13g2_nor2b_1 _1570_ (.A(net20),
    .B_N(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit10.Q ),
    .Y(_0233_));
 sg13g2_nor2_1 _1571_ (.A(net49),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit10.Q ),
    .Y(_0234_));
 sg13g2_nor3_1 _1572_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit11.Q ),
    .B(_0233_),
    .C(_0234_),
    .Y(_0235_));
 sg13g2_nor2_1 _1573_ (.A(_0232_),
    .B(_0235_),
    .Y(_0236_));
 sg13g2_mux4_1 _1574_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit10.Q ),
    .A0(net50),
    .A1(net21),
    .A2(net78),
    .A3(net105),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit11.Q ),
    .X(_0237_));
 sg13g2_mux4_1 _1575_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit11.Q ),
    .A0(net54),
    .A1(net93),
    .A2(net9),
    .A3(\Inst_LUT4AB_switch_matrix.JN2BEG3 ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit10.Q ),
    .X(_0238_));
 sg13g2_mux4_1 _1576_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit11.Q ),
    .A0(net42),
    .A1(net70),
    .A2(net24),
    .A3(net97),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit10.Q ),
    .X(_0239_));
 sg13g2_nand2_1 _1577_ (.Y(_0240_),
    .A(\Inst_LE_LUT4c_frame_config_dffesr.c_I0mux ),
    .B(_0209_));
 sg13g2_nand2_1 _1578_ (.Y(_0241_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit11.Q ),
    .B(_0237_));
 sg13g2_o21ai_1 _1579_ (.B1(_0241_),
    .Y(_0242_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit11.Q ),
    .A2(_0236_));
 sg13g2_nor2b_1 _1580_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit11.Q ),
    .B_N(_0239_),
    .Y(_0243_));
 sg13g2_a21oi_2 _1581_ (.B1(_0243_),
    .Y(_0244_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit11.Q ),
    .A1(_0238_));
 sg13g2_a21oi_2 _1582_ (.B1(\Inst_LE_LUT4c_frame_config_dffesr.c_I0mux ),
    .Y(_0245_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit12.Q ),
    .A1(_0244_));
 sg13g2_o21ai_1 _1583_ (.B1(_0245_),
    .Y(_0246_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit12.Q ),
    .A2(_0242_));
 sg13g2_nand2_2 _1584_ (.Y(_0247_),
    .A(_0246_),
    .B(_0240_));
 sg13g2_mux4_1 _1585_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit14.Q ),
    .A0(net52),
    .A1(net84),
    .A2(net94),
    .A3(\Inst_LUT4AB_switch_matrix.JS2BEG3 ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit15.Q ),
    .X(_0248_));
 sg13g2_mux2_1 _1586_ (.A0(net40),
    .A1(net11),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit14.Q ),
    .X(_0249_));
 sg13g2_nand2b_1 _1587_ (.Y(_0250_),
    .B(net84),
    .A_N(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit14.Q ));
 sg13g2_nand2_1 _1588_ (.Y(_0251_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit14.Q ),
    .B(net95));
 sg13g2_nand3_1 _1589_ (.B(_0250_),
    .C(_0251_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit15.Q ),
    .Y(_0252_));
 sg13g2_o21ai_1 _1590_ (.B1(_0252_),
    .Y(_0253_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit15.Q ),
    .A2(_0249_));
 sg13g2_o21ai_1 _1591_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit16.Q ),
    .Y(_0254_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit15.Q ),
    .A2(_0253_));
 sg13g2_a21oi_1 _1592_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit15.Q ),
    .A2(_0248_),
    .Y(_0255_),
    .B1(_0254_));
 sg13g2_mux4_1 _1593_ (.S0(net987),
    .A0(net977),
    .A1(net971),
    .A2(net941),
    .A3(net946),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit15.Q ),
    .X(_0256_));
 sg13g2_and2_1 _1594_ (.A(_1042_),
    .B(_0256_),
    .X(_0257_));
 sg13g2_nor2_1 _1595_ (.A(net987),
    .B(net965),
    .Y(_0258_));
 sg13g2_a21oi_1 _1596_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit14.Q ),
    .A2(_1051_),
    .Y(_0259_),
    .B1(_0258_));
 sg13g2_mux2_1 _1597_ (.A0(net936),
    .A1(\Inst_LUT4AB_switch_matrix.M_EF ),
    .S(net987),
    .X(_0260_));
 sg13g2_nor2b_1 _1598_ (.A(_0260_),
    .B_N(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit15.Q ),
    .Y(_0261_));
 sg13g2_o21ai_1 _1599_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit16.Q ),
    .Y(_0262_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit15.Q ),
    .A2(_0259_));
 sg13g2_o21ai_1 _1600_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit17.Q ),
    .Y(_0263_),
    .A1(_0261_),
    .A2(_0262_));
 sg13g2_o21ai_1 _1601_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit15.Q ),
    .Y(_0264_),
    .A1(_1013_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit14.Q ));
 sg13g2_a21oi_1 _1602_ (.A1(net12),
    .A2(net987),
    .Y(_0265_),
    .B1(_0264_));
 sg13g2_mux2_1 _1603_ (.A0(net1008),
    .A1(net41),
    .S(net987),
    .X(_0266_));
 sg13g2_o21ai_1 _1604_ (.B1(_1042_),
    .Y(_0267_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit15.Q ),
    .A2(_0266_));
 sg13g2_nor2_1 _1605_ (.A(_0265_),
    .B(_0267_),
    .Y(_0268_));
 sg13g2_nand2b_1 _1606_ (.Y(_0269_),
    .B(net987),
    .A_N(net1004));
 sg13g2_o21ai_1 _1607_ (.B1(_0269_),
    .Y(_0270_),
    .A1(net87),
    .A2(net987));
 sg13g2_mux2_1 _1608_ (.A0(net61),
    .A1(net69),
    .S(net987),
    .X(_0271_));
 sg13g2_o21ai_1 _1609_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit16.Q ),
    .Y(_0272_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit15.Q ),
    .A2(_0271_));
 sg13g2_a21oi_1 _1610_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit15.Q ),
    .A2(_0270_),
    .Y(_0273_),
    .B1(_0272_));
 sg13g2_or3_1 _1611_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit17.Q ),
    .B(_0268_),
    .C(_0273_),
    .X(_0274_));
 sg13g2_o21ai_1 _1612_ (.B1(_0274_),
    .Y(_0275_),
    .A1(_0263_),
    .A2(_0257_));
 sg13g2_inv_1 _1613_ (.Y(\Inst_LUT4AB_switch_matrix.JS2BEG5 ),
    .A(_0275_));
 sg13g2_mux4_1 _1614_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit15.Q ),
    .A0(_1021_),
    .A1(_1026_),
    .A2(_1034_),
    .A3(_0275_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit14.Q ),
    .X(_0276_));
 sg13g2_mux4_1 _1615_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit14.Q ),
    .A0(net48),
    .A1(net19),
    .A2(net76),
    .A3(net103),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit15.Q ),
    .X(_0277_));
 sg13g2_a21oi_1 _1616_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit15.Q ),
    .A2(_0277_),
    .Y(_0278_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit16.Q ));
 sg13g2_o21ai_1 _1617_ (.B1(_0278_),
    .Y(_0279_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit15.Q ),
    .A2(_0276_));
 sg13g2_nor2b_1 _1618_ (.A(_0255_),
    .B_N(_0279_),
    .Y(_0280_));
 sg13g2_inv_1 _1619_ (.Y(_0281_),
    .A(_0280_));
 sg13g2_mux2_1 _1620_ (.A0(net57),
    .A1(net8),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit12.Q ),
    .X(_0282_));
 sg13g2_nor2b_1 _1621_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit12.Q ),
    .B_N(net81),
    .Y(_0283_));
 sg13g2_a21oi_2 _1622_ (.B1(_0283_),
    .Y(_0284_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit12.Q ),
    .A1(\Inst_LUT4AB_switch_matrix.E2BEG3 ));
 sg13g2_nand2_2 _1623_ (.Y(_0285_),
    .A(_0284_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit13.Q ));
 sg13g2_o21ai_1 _1624_ (.B1(_0285_),
    .Y(_0286_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit13.Q ),
    .A2(_0282_));
 sg13g2_o21ai_1 _1625_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit13.Q ),
    .Y(_0287_),
    .A1(net66),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit12.Q ));
 sg13g2_a21oi_1 _1626_ (.A1(_1030_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit12.Q ),
    .Y(_0288_),
    .B1(_0287_));
 sg13g2_mux2_1 _1627_ (.A0(net38),
    .A1(net9),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit12.Q ),
    .X(_0289_));
 sg13g2_a21oi_1 _1628_ (.A1(_1041_),
    .A2(_0289_),
    .Y(_0290_),
    .B1(_0288_));
 sg13g2_mux4_1 _1629_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit14.Q ),
    .A0(net979),
    .A1(net973),
    .A2(net943),
    .A3(net948),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit15.Q ),
    .X(_0291_));
 sg13g2_mux4_1 _1630_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit14.Q ),
    .A0(net967),
    .A1(net953),
    .A2(net937),
    .A3(net930),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit15.Q ),
    .X(_0292_));
 sg13g2_nand2b_1 _1631_ (.Y(_0293_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit16.Q ),
    .A_N(_0292_));
 sg13g2_o21ai_1 _1632_ (.B1(_0293_),
    .Y(_0294_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit16.Q ),
    .A2(_0291_));
 sg13g2_mux4_1 _1633_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit14.Q ),
    .A0(net1008),
    .A1(net41),
    .A2(net1215),
    .A3(net12),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit15.Q ),
    .X(_0295_));
 sg13g2_nand2b_1 _1634_ (.Y(_0296_),
    .B(_0295_),
    .A_N(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit16.Q ));
 sg13g2_mux2_1 _1635_ (.A0(net59),
    .A1(net61),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit14.Q ),
    .X(_0297_));
 sg13g2_nand2b_1 _1636_ (.Y(_0298_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit14.Q ),
    .A_N(net1005));
 sg13g2_o21ai_1 _1637_ (.B1(_0298_),
    .Y(_0299_),
    .A1(net69),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit14.Q ));
 sg13g2_o21ai_1 _1638_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit16.Q ),
    .Y(_0300_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit15.Q ),
    .A2(_0297_));
 sg13g2_a21oi_1 _1639_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit15.Q ),
    .A2(_0299_),
    .Y(_0301_),
    .B1(_0300_));
 sg13g2_nor2_1 _1640_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit17.Q ),
    .B(_0301_),
    .Y(_0302_));
 sg13g2_a22oi_1 _1641_ (.Y(\Inst_LUT4AB_switch_matrix.E2BEG5 ),
    .B1(_0296_),
    .B2(_0302_),
    .A2(_0294_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit17.Q ));
 sg13g2_mux2_1 _1642_ (.A0(net45),
    .A1(net16),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit12.Q ),
    .X(_0303_));
 sg13g2_nand2_1 _1643_ (.Y(_0304_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit12.Q ),
    .B(\Inst_LUT4AB_switch_matrix.E2BEG5 ));
 sg13g2_nand2b_1 _1644_ (.Y(_0305_),
    .B(net73),
    .A_N(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit12.Q ));
 sg13g2_nand3_1 _1645_ (.B(_0304_),
    .C(_0305_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit13.Q ),
    .Y(_0306_));
 sg13g2_o21ai_1 _1646_ (.B1(_0306_),
    .Y(_0307_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit13.Q ),
    .A2(_0303_));
 sg13g2_mux4_1 _1647_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit12.Q ),
    .A0(net46),
    .A1(net17),
    .A2(net74),
    .A3(net101),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit13.Q ),
    .X(_0308_));
 sg13g2_inv_1 _1648_ (.Y(_0309_),
    .A(_0308_));
 sg13g2_mux4_1 _1649_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit13.Q ),
    .A0(_0307_),
    .A1(_0309_),
    .A2(_0290_),
    .A3(_0286_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit14.Q ),
    .X(_0310_));
 sg13g2_nand2_1 _1650_ (.Y(_0311_),
    .A(_0281_),
    .B(_0310_));
 sg13g2_nor2_1 _1651_ (.A(_0281_),
    .B(_0310_),
    .Y(_0312_));
 sg13g2_mux4_1 _1652_ (.S0(_0280_),
    .A0(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ),
    .A1(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ),
    .A2(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ),
    .A3(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ),
    .S1(_0310_),
    .X(_0313_));
 sg13g2_nor2b_1 _1653_ (.A(_0313_),
    .B_N(_0247_),
    .Y(_0314_));
 sg13g2_mux4_1 _1654_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit17.Q ),
    .A0(_1040_),
    .A1(_1030_),
    .A2(_1022_),
    .A3(_0037_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit16.Q ),
    .X(_0315_));
 sg13g2_mux4_1 _1655_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit16.Q ),
    .A0(net57),
    .A1(net7),
    .A2(net64),
    .A3(net91),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit17.Q ),
    .X(_0316_));
 sg13g2_mux4_1 _1656_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit14.Q ),
    .A0(net977),
    .A1(net972),
    .A2(net942),
    .A3(net947),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit15.Q ),
    .X(_0317_));
 sg13g2_mux4_1 _1657_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit14.Q ),
    .A0(net966),
    .A1(net953),
    .A2(net937),
    .A3(net928),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit15.Q ),
    .X(_0318_));
 sg13g2_nand2b_1 _1658_ (.Y(_0319_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit16.Q ),
    .A_N(_0318_));
 sg13g2_o21ai_1 _1659_ (.B1(_0319_),
    .Y(_0320_),
    .A1(_0317_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit16.Q ));
 sg13g2_mux4_1 _1660_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit14.Q ),
    .A0(net1008),
    .A1(net41),
    .A2(net1215),
    .A3(net12),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit15.Q ),
    .X(_0321_));
 sg13g2_nand2b_1 _1661_ (.Y(_0322_),
    .B(_0321_),
    .A_N(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit16.Q ));
 sg13g2_nand2b_1 _1662_ (.Y(_0323_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit14.Q ),
    .A_N(net1004));
 sg13g2_o21ai_1 _1663_ (.B1(_0323_),
    .Y(_0324_),
    .A1(net69),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit14.Q ));
 sg13g2_mux2_1 _1664_ (.A0(net59),
    .A1(net61),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit14.Q ),
    .X(_0325_));
 sg13g2_o21ai_1 _1665_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit16.Q ),
    .Y(_0326_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit15.Q ),
    .A2(_0325_));
 sg13g2_a21oi_1 _1666_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit15.Q ),
    .A2(_0324_),
    .Y(_0327_),
    .B1(_0326_));
 sg13g2_nor2_1 _1667_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit17.Q ),
    .B(_0327_),
    .Y(_0328_));
 sg13g2_a22oi_1 _1668_ (.Y(\Inst_LUT4AB_switch_matrix.JW2BEG5 ),
    .B1(_0322_),
    .B2(_0328_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit17.Q ),
    .A1(_0320_));
 sg13g2_mux4_1 _1669_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit16.Q ),
    .A0(net14),
    .A1(net71),
    .A2(net98),
    .A3(net377),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit17.Q ),
    .X(_0329_));
 sg13g2_mux2_1 _1670_ (.A0(net44),
    .A1(net15),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit16.Q ),
    .X(_0330_));
 sg13g2_nand2b_1 _1671_ (.Y(_0331_),
    .B(net72),
    .A_N(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit16.Q ));
 sg13g2_nand2_1 _1672_ (.Y(_0332_),
    .A(net99),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit16.Q ));
 sg13g2_nand3_1 _1673_ (.B(_0331_),
    .C(_0332_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit17.Q ),
    .Y(_0333_));
 sg13g2_o21ai_1 _1674_ (.B1(_0333_),
    .Y(_0334_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit17.Q ),
    .A2(_0330_));
 sg13g2_a21oi_1 _1675_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit17.Q ),
    .A2(_0315_),
    .Y(_0335_),
    .B1(_1043_));
 sg13g2_o21ai_1 _1676_ (.B1(_0335_),
    .Y(_0336_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit17.Q ),
    .A2(_0316_));
 sg13g2_nand2_1 _1677_ (.Y(_0337_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit17.Q ),
    .B(_0334_));
 sg13g2_o21ai_1 _1678_ (.B1(_0337_),
    .Y(_0338_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit17.Q ),
    .A2(_0329_));
 sg13g2_o21ai_1 _1679_ (.B1(_0336_),
    .Y(_0339_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit18.Q ),
    .A2(_0338_));
 sg13g2_mux4_1 _1680_ (.S0(_0280_),
    .A0(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ),
    .A1(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ),
    .A2(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ),
    .A3(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ),
    .S1(_0310_),
    .X(_0340_));
 sg13g2_nor2_1 _1681_ (.A(_0247_),
    .B(_0340_),
    .Y(_0341_));
 sg13g2_nor3_2 _1682_ (.A(_0341_),
    .B(_0339_),
    .C(_0314_),
    .Y(_0342_));
 sg13g2_mux4_1 _1683_ (.S0(_0280_),
    .A0(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ),
    .A1(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ),
    .A2(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ),
    .A3(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ),
    .S1(_0310_),
    .X(_0343_));
 sg13g2_or2_1 _1684_ (.X(_0344_),
    .B(_0343_),
    .A(_0247_));
 sg13g2_mux4_1 _1685_ (.S0(_0280_),
    .A0(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ),
    .A1(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ),
    .A2(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ),
    .A3(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ),
    .S1(_0310_),
    .X(_0345_));
 sg13g2_nand2b_1 _1686_ (.Y(_0346_),
    .B(_0247_),
    .A_N(_0345_));
 sg13g2_nand3_1 _1687_ (.B(_0344_),
    .C(_0346_),
    .A(_0339_),
    .Y(_0347_));
 sg13g2_nand2b_1 _1688_ (.Y(_0348_),
    .B(_0347_),
    .A_N(_0342_));
 sg13g2_mux2_1 _1689_ (.A0(_0348_),
    .A1(\Inst_LE_LUT4c_frame_config_dffesr.LUT_flop ),
    .S(\Inst_LE_LUT4c_frame_config_dffesr.c_out_mux ),
    .X(E));
 sg13g2_mux4_1 _1690_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit2.Q ),
    .A0(net978),
    .A1(net973),
    .A2(net948),
    .A3(net967),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit3.Q ),
    .X(_0349_));
 sg13g2_mux4_1 _1691_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit2.Q ),
    .A0(net960),
    .A1(net954),
    .A2(net936),
    .A3(net928),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit3.Q ),
    .X(_0350_));
 sg13g2_nand2b_1 _1692_ (.Y(_0351_),
    .B(_1031_),
    .A_N(_0349_));
 sg13g2_o21ai_1 _1693_ (.B1(_0351_),
    .Y(_0352_),
    .A1(_1031_),
    .A2(_0350_));
 sg13g2_mux4_1 _1694_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit2.Q ),
    .A0(net38),
    .A1(net54),
    .A2(net3),
    .A3(net9),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit3.Q ),
    .X(_0353_));
 sg13g2_nand2_1 _1695_ (.Y(_0354_),
    .A(_1031_),
    .B(_0353_));
 sg13g2_mux2_1 _1696_ (.A0(net1211),
    .A1(net66),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit2.Q ),
    .X(_0355_));
 sg13g2_or2_1 _1697_ (.X(_0356_),
    .B(_0355_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit3.Q ));
 sg13g2_nand2_1 _1698_ (.Y(_0357_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit2.Q ),
    .B(_1030_));
 sg13g2_o21ai_1 _1699_ (.B1(_0357_),
    .Y(_0358_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit2.Q ),
    .A2(net93));
 sg13g2_a21oi_1 _1700_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit3.Q ),
    .A2(_0358_),
    .Y(_0359_),
    .B1(_1031_));
 sg13g2_a21oi_1 _1701_ (.A1(_0356_),
    .A2(_0359_),
    .Y(_0360_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit5.Q ));
 sg13g2_a22oi_1 _1702_ (.Y(\Inst_LUT4AB_switch_matrix.JN2BEG2 ),
    .B1(_0354_),
    .B2(_0360_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit5.Q ),
    .A1(_0352_));
 sg13g2_mux2_1 _1703_ (.A0(net9),
    .A1(net86),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit2.Q ),
    .X(_0361_));
 sg13g2_nor2_1 _1704_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit3.Q ),
    .B(_0361_),
    .Y(_0362_));
 sg13g2_o21ai_1 _1705_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit3.Q ),
    .Y(_0363_),
    .A1(_1023_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit2.Q ));
 sg13g2_a21oi_1 _1706_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit2.Q ),
    .A2(\Inst_LUT4AB_switch_matrix.JN2BEG2 ),
    .Y(_0364_),
    .B1(_0363_));
 sg13g2_or2_1 _1707_ (.X(_0365_),
    .B(_0364_),
    .A(_0362_));
 sg13g2_mux4_1 _1708_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit3.Q ),
    .A0(net58),
    .A1(net69),
    .A2(net12),
    .A3(net96),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit2.Q ),
    .X(_0366_));
 sg13g2_o21ai_1 _1709_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit24.Q ),
    .Y(_0367_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit23.Q ),
    .A2(_0366_));
 sg13g2_a21oi_1 _1710_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit23.Q ),
    .A2(_0365_),
    .Y(_0368_),
    .B1(_0367_));
 sg13g2_mux4_1 _1711_ (.S0(net999),
    .A0(net976),
    .A1(net971),
    .A2(net941),
    .A3(net946),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit11.Q ),
    .X(_0369_));
 sg13g2_nand2b_1 _1712_ (.Y(_0370_),
    .B(_0369_),
    .A_N(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit12.Q ));
 sg13g2_nor2_1 _1713_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit10.Q ),
    .B(net958),
    .Y(_0371_));
 sg13g2_a21oi_1 _1714_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit10.Q ),
    .A2(_1051_),
    .Y(_0372_),
    .B1(_0371_));
 sg13g2_nand2b_1 _1715_ (.Y(_0373_),
    .B(net999),
    .A_N(net930));
 sg13g2_o21ai_1 _1716_ (.B1(_0373_),
    .Y(_0374_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit10.Q ),
    .A2(net936));
 sg13g2_o21ai_1 _1717_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit12.Q ),
    .Y(_0375_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit11.Q ),
    .A2(_0372_));
 sg13g2_a21oi_1 _1718_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit11.Q ),
    .A2(_0374_),
    .Y(_0376_),
    .B1(_0375_));
 sg13g2_nor2b_1 _1719_ (.A(_0376_),
    .B_N(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit13.Q ),
    .Y(_0377_));
 sg13g2_nand2b_1 _1720_ (.Y(_0378_),
    .B(net999),
    .A_N(net11));
 sg13g2_o21ai_1 _1721_ (.B1(_0378_),
    .Y(_0379_),
    .A1(net999),
    .A2(net1216));
 sg13g2_mux2_1 _1722_ (.A0(net32),
    .A1(net40),
    .S(net999),
    .X(_0380_));
 sg13g2_a21oi_1 _1723_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit11.Q ),
    .A2(_0379_),
    .Y(_0381_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit12.Q ));
 sg13g2_o21ai_1 _1724_ (.B1(_0381_),
    .Y(_0382_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit11.Q ),
    .A2(_0380_));
 sg13g2_nand2b_1 _1725_ (.Y(_0383_),
    .B(net999),
    .A_N(net89));
 sg13g2_o21ai_1 _1726_ (.B1(_0383_),
    .Y(_0384_),
    .A1(net1006),
    .A2(net999));
 sg13g2_mux2_1 _1727_ (.A0(net60),
    .A1(net68),
    .S(net999),
    .X(_0385_));
 sg13g2_o21ai_1 _1728_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit12.Q ),
    .Y(_0386_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit11.Q ),
    .A2(_0385_));
 sg13g2_a21oi_1 _1729_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit11.Q ),
    .A2(_0384_),
    .Y(_0387_),
    .B1(_0386_));
 sg13g2_nor2_1 _1730_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit13.Q ),
    .B(_0387_),
    .Y(_0388_));
 sg13g2_a22oi_1 _1731_ (.Y(\Inst_LUT4AB_switch_matrix.JN2BEG4 ),
    .B1(_0382_),
    .B2(_0388_),
    .A2(_0370_),
    .A1(_0377_));
 sg13g2_mux4_1 _1732_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit3.Q ),
    .A0(net20),
    .A1(net104),
    .A2(net77),
    .A3(\Inst_LUT4AB_switch_matrix.JN2BEG4 ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit2.Q ),
    .X(_0389_));
 sg13g2_mux4_1 _1733_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit2.Q ),
    .A0(net50),
    .A1(net21),
    .A2(net78),
    .A3(net105),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit3.Q ),
    .X(_0390_));
 sg13g2_inv_1 _1734_ (.Y(_0391_),
    .A(_0390_));
 sg13g2_a21oi_1 _1735_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit23.Q ),
    .A2(_0391_),
    .Y(_0392_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit24.Q ));
 sg13g2_o21ai_1 _1736_ (.B1(_0392_),
    .Y(_0393_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit23.Q ),
    .A2(_0389_));
 sg13g2_nand2b_1 _1737_ (.Y(_0394_),
    .B(_0393_),
    .A_N(_0368_));
 sg13g2_mux2_1 _1738_ (.A0(_0394_),
    .A1(_0207_),
    .S(\Inst_LC_LUT4c_frame_config_dffesr.c_I0mux ),
    .X(_0395_));
 sg13g2_nand2_1 _1739_ (.Y(_0396_),
    .A(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ),
    .B(net926));
 sg13g2_nand2b_1 _1740_ (.Y(_0397_),
    .B(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ),
    .A_N(net926));
 sg13g2_nand3_1 _1741_ (.B(_0396_),
    .C(_0397_),
    .A(_0206_),
    .Y(_0398_));
 sg13g2_nand2b_1 _1742_ (.Y(_0399_),
    .B(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ),
    .A_N(net926));
 sg13g2_nand3b_1 _1743_ (.B(_0203_),
    .C(_0399_),
    .Y(_0400_),
    .A_N(_0202_));
 sg13g2_a21oi_1 _1744_ (.A1(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ),
    .A2(net926),
    .Y(_0401_),
    .B1(_0400_));
 sg13g2_mux4_1 _1745_ (.S0(net985),
    .A0(net975),
    .A1(net968),
    .A2(net944),
    .A3(net961),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit3.Q ),
    .X(_0402_));
 sg13g2_nand2b_1 _1746_ (.Y(_0403_),
    .B(_0402_),
    .A_N(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit4.Q ));
 sg13g2_nor2_2 _1747_ (.A(net985),
    .B(net955),
    .Y(_0404_));
 sg13g2_a21oi_2 _1748_ (.B1(_0404_),
    .Y(_0405_),
    .A2(_1051_),
    .A1(net985));
 sg13g2_nand2b_1 _1749_ (.Y(_0406_),
    .B(net985),
    .A_N(net929));
 sg13g2_o21ai_1 _1750_ (.B1(_0406_),
    .Y(_0407_),
    .A1(net985),
    .A2(net934));
 sg13g2_o21ai_1 _1751_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit4.Q ),
    .Y(_0408_),
    .A1(_0405_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit3.Q ));
 sg13g2_a21oi_2 _1752_ (.B1(_0408_),
    .Y(_0409_),
    .A2(_0407_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit3.Q ));
 sg13g2_nor2b_1 _1753_ (.A(_0409_),
    .B_N(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit5.Q ),
    .Y(_0410_));
 sg13g2_mux2_1 _1754_ (.A0(net82),
    .A1(net86),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit2.Q ),
    .X(_0411_));
 sg13g2_nand2_1 _1755_ (.Y(_0412_),
    .A(_1028_),
    .B(net985));
 sg13g2_o21ai_1 _1756_ (.B1(_0412_),
    .Y(_0413_),
    .A1(net93),
    .A2(net985));
 sg13g2_o21ai_1 _1757_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit4.Q ),
    .Y(_0414_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit3.Q ),
    .A2(_0411_));
 sg13g2_a21oi_1 _1758_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit3.Q ),
    .A2(_0413_),
    .Y(_0415_),
    .B1(_0414_));
 sg13g2_mux4_1 _1759_ (.S0(net985),
    .A0(net1009),
    .A1(net38),
    .A2(net25),
    .A3(net1210),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit3.Q ),
    .X(_0416_));
 sg13g2_nand2b_1 _1760_ (.Y(_0417_),
    .B(_0416_),
    .A_N(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit4.Q ));
 sg13g2_nor2_1 _1761_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit5.Q ),
    .B(_0415_),
    .Y(_0418_));
 sg13g2_a22oi_1 _1762_ (.Y(\Inst_LUT4AB_switch_matrix.JW2BEG2 ),
    .B1(_0417_),
    .B2(_0418_),
    .A2(_0403_),
    .A1(_0410_));
 sg13g2_nand2_1 _1763_ (.Y(_0419_),
    .A(net83),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit8.Q ));
 sg13g2_o21ai_1 _1764_ (.B1(_0419_),
    .Y(_0420_),
    .A1(_1012_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit8.Q ));
 sg13g2_nand2_2 _1765_ (.Y(_0421_),
    .A(\Inst_LUT4AB_switch_matrix.JW2BEG2 ),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit8.Q ));
 sg13g2_nand2b_1 _1766_ (.Y(_0422_),
    .B(net106),
    .A_N(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit8.Q ));
 sg13g2_nand3_1 _1767_ (.B(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit9.Q ),
    .C(_0422_),
    .A(_0421_),
    .Y(_0423_));
 sg13g2_o21ai_1 _1768_ (.B1(_0423_),
    .Y(_0424_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit9.Q ),
    .A2(_0420_));
 sg13g2_inv_2 _1769_ (.Y(_0425_),
    .A(_0424_));
 sg13g2_mux2_1 _1770_ (.A0(net35),
    .A1(net23),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit8.Q ),
    .X(_0426_));
 sg13g2_nand2b_1 _1771_ (.Y(_0427_),
    .B(net63),
    .A_N(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit8.Q ));
 sg13g2_nand2_1 _1772_ (.Y(_0428_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit8.Q ),
    .B(net90));
 sg13g2_nand3_1 _1773_ (.B(_0427_),
    .C(_0428_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit9.Q ),
    .Y(_0429_));
 sg13g2_o21ai_1 _1774_ (.B1(_0429_),
    .Y(_0430_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit9.Q ),
    .A2(_0426_));
 sg13g2_o21ai_1 _1775_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit30.Q ),
    .Y(_0431_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit29.Q ),
    .A2(_0430_));
 sg13g2_a21oi_2 _1776_ (.B1(_0431_),
    .Y(_0432_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit29.Q ),
    .A1(_0425_));
 sg13g2_mux4_1 _1777_ (.S0(net984),
    .A0(net976),
    .A1(net971),
    .A2(net941),
    .A3(net946),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit11.Q ),
    .X(_0433_));
 sg13g2_nor2_1 _1778_ (.A(net984),
    .B(net958),
    .Y(_0434_));
 sg13g2_a21oi_1 _1779_ (.A1(net984),
    .A2(_1051_),
    .Y(_0435_),
    .B1(_0434_));
 sg13g2_o21ai_1 _1780_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit11.Q ),
    .Y(_0436_),
    .A1(net984),
    .A2(net933));
 sg13g2_a21oi_2 _1781_ (.B1(_0436_),
    .Y(_0437_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit10.Q ),
    .A1(\Inst_LUT4AB_switch_matrix.M_AD ));
 sg13g2_o21ai_1 _1782_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit12.Q ),
    .Y(_0438_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit11.Q ),
    .A2(_0435_));
 sg13g2_o21ai_1 _1783_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit13.Q ),
    .Y(_0439_),
    .A1(_0438_),
    .A2(_0437_));
 sg13g2_a21oi_2 _1784_ (.B1(_0439_),
    .Y(_0440_),
    .A2(_0433_),
    .A1(_1039_));
 sg13g2_mux4_1 _1785_ (.S0(net984),
    .A0(net1009),
    .A1(net40),
    .A2(net1216),
    .A3(net11),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit11.Q ),
    .X(_0441_));
 sg13g2_nand2b_1 _1786_ (.Y(_0442_),
    .B(net984),
    .A_N(net1006));
 sg13g2_o21ai_1 _1787_ (.B1(_0442_),
    .Y(_0443_),
    .A1(net68),
    .A2(net984));
 sg13g2_mux2_1 _1788_ (.A0(net60),
    .A1(net62),
    .S(net984),
    .X(_0444_));
 sg13g2_or2_1 _1789_ (.X(_0445_),
    .B(_0444_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit11.Q ));
 sg13g2_a21oi_1 _1790_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit11.Q ),
    .A2(_0443_),
    .Y(_0446_),
    .B1(_1039_));
 sg13g2_a221oi_1 _1791_ (.B2(_0446_),
    .C1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit13.Q ),
    .B1(_0445_),
    .A1(_1039_),
    .Y(_0447_),
    .A2(_0441_));
 sg13g2_nor2_2 _1792_ (.A(_0447_),
    .B(_0440_),
    .Y(\Inst_LUT4AB_switch_matrix.JW2BEG4 ));
 sg13g2_nor2b_1 _1793_ (.A(\Inst_LUT4AB_switch_matrix.JW2BEG4 ),
    .B_N(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit8.Q ),
    .Y(_0448_));
 sg13g2_nor2_1 _1794_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit8.Q ),
    .B(net98),
    .Y(_0449_));
 sg13g2_o21ai_1 _1795_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit9.Q ),
    .Y(_0450_),
    .A1(_0449_),
    .A2(_0448_));
 sg13g2_mux2_1 _1796_ (.A0(net43),
    .A1(net71),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit8.Q ),
    .X(_0451_));
 sg13g2_o21ai_1 _1797_ (.B1(_0450_),
    .Y(_0452_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit9.Q ),
    .A2(_0451_));
 sg13g2_mux4_1 _1798_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit8.Q ),
    .A0(net44),
    .A1(net15),
    .A2(net72),
    .A3(net99),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit9.Q ),
    .X(_0453_));
 sg13g2_inv_1 _1799_ (.Y(_0454_),
    .A(_0453_));
 sg13g2_a21oi_1 _1800_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit29.Q ),
    .A2(_0453_),
    .Y(_0455_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit30.Q ));
 sg13g2_o21ai_1 _1801_ (.B1(_0455_),
    .Y(_0456_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit29.Q ),
    .A2(_0452_));
 sg13g2_nor2b_2 _1802_ (.A(_0432_),
    .B_N(_0456_),
    .Y(_0457_));
 sg13g2_nand2b_1 _1803_ (.Y(_0458_),
    .B(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ),
    .A_N(net926));
 sg13g2_nand3b_1 _1804_ (.B(_0458_),
    .C(_0202_),
    .Y(_0459_),
    .A_N(_0203_));
 sg13g2_a21oi_1 _1805_ (.A1(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ),
    .A2(net926),
    .Y(_0460_),
    .B1(_0459_));
 sg13g2_mux2_1 _1806_ (.A0(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ),
    .A1(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ),
    .S(net926),
    .X(_0461_));
 sg13g2_o21ai_1 _1807_ (.B1(_0398_),
    .Y(_0462_),
    .A1(_0204_),
    .A2(_0461_));
 sg13g2_nor4_2 _1808_ (.A(_0401_),
    .B(_0462_),
    .C(_0460_),
    .Y(_0463_),
    .D(_0457_));
 sg13g2_mux4_1 _1809_ (.S0(_0202_),
    .A0(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ),
    .A1(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ),
    .A2(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ),
    .A3(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ),
    .S1(net926),
    .X(_0464_));
 sg13g2_mux4_1 _1810_ (.S0(_0202_),
    .A0(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ),
    .A1(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ),
    .A2(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ),
    .A3(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ),
    .S1(_0395_),
    .X(_0465_));
 sg13g2_mux2_1 _1811_ (.A0(_0464_),
    .A1(_0465_),
    .S(_0203_),
    .X(_0466_));
 sg13g2_a21o_1 _1812_ (.A2(_0466_),
    .A1(_0457_),
    .B1(_0463_),
    .X(_0467_));
 sg13g2_mux2_1 _1813_ (.A0(_0467_),
    .A1(\Inst_LC_LUT4c_frame_config_dffesr.LUT_flop ),
    .S(\Inst_LC_LUT4c_frame_config_dffesr.c_out_mux ),
    .X(C));
 sg13g2_nor2_1 _1814_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit27.Q ),
    .B(_0316_),
    .Y(_0468_));
 sg13g2_a21oi_1 _1815_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit27.Q ),
    .A2(_0315_),
    .Y(_0469_),
    .B1(_0468_));
 sg13g2_nand2_1 _1816_ (.Y(_0470_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit27.Q ),
    .B(_0334_));
 sg13g2_nor2_1 _1817_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit27.Q ),
    .B(_0329_),
    .Y(_0471_));
 sg13g2_nor2_1 _1818_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit28.Q ),
    .B(_0471_),
    .Y(_0472_));
 sg13g2_a22oi_1 _1819_ (.Y(_0473_),
    .B1(_0470_),
    .B2(_0472_),
    .A2(_0469_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit28.Q ));
 sg13g2_nand2_1 _1820_ (.Y(_0474_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit21.Q ),
    .B(_0237_));
 sg13g2_o21ai_1 _1821_ (.B1(_0474_),
    .Y(_0475_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit21.Q ),
    .A2(_0236_));
 sg13g2_or2_1 _1822_ (.X(_0476_),
    .B(_0475_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit22.Q ));
 sg13g2_nor2b_1 _1823_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit21.Q ),
    .B_N(_0239_),
    .Y(_0477_));
 sg13g2_a21oi_1 _1824_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit21.Q ),
    .A2(_0238_),
    .Y(_0478_),
    .B1(_0477_));
 sg13g2_a21o_1 _1825_ (.A2(_0209_),
    .A1(_0311_),
    .B1(_0312_),
    .X(_0479_));
 sg13g2_a21oi_1 _1826_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit22.Q ),
    .A2(_0478_),
    .Y(_0480_),
    .B1(\Inst_LF_LUT4c_frame_config_dffesr.c_I0mux ));
 sg13g2_a22oi_1 _1827_ (.Y(_0481_),
    .B1(_0480_),
    .B2(_0476_),
    .A2(\Inst_LF_LUT4c_frame_config_dffesr.c_I0mux ),
    .A1(_0479_));
 sg13g2_o21ai_1 _1828_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit26.Q ),
    .Y(_0482_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit25.Q ),
    .A2(_0253_));
 sg13g2_a21oi_2 _1829_ (.B1(_0482_),
    .Y(_0483_),
    .A2(_0248_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit25.Q ));
 sg13g2_a21oi_1 _1830_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit25.Q ),
    .A2(_0277_),
    .Y(_0484_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit26.Q ));
 sg13g2_o21ai_1 _1831_ (.B1(_0484_),
    .Y(_0485_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit25.Q ),
    .A2(_0276_));
 sg13g2_nand2b_2 _1832_ (.Y(_0486_),
    .B(_0485_),
    .A_N(_0483_));
 sg13g2_mux4_1 _1833_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit23.Q ),
    .A0(_0307_),
    .A1(_0309_),
    .A2(_0290_),
    .A3(_0286_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit24.Q ),
    .X(_0487_));
 sg13g2_nor2_1 _1834_ (.A(_0486_),
    .B(_0487_),
    .Y(_0488_));
 sg13g2_mux4_1 _1835_ (.S0(_0481_),
    .A0(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ),
    .A1(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ),
    .A2(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ),
    .A3(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ),
    .S1(_0487_),
    .X(_0489_));
 sg13g2_nand2_1 _1836_ (.Y(_0490_),
    .A(_0486_),
    .B(_0487_));
 sg13g2_mux4_1 _1837_ (.S0(_0481_),
    .A0(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ),
    .A1(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ),
    .A2(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ),
    .A3(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ),
    .S1(_0487_),
    .X(_0491_));
 sg13g2_mux2_1 _1838_ (.A0(_0489_),
    .A1(_0491_),
    .S(_0486_),
    .X(_0492_));
 sg13g2_mux4_1 _1839_ (.S0(_0481_),
    .A0(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ),
    .A1(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ),
    .A2(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ),
    .A3(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ),
    .S1(_0487_),
    .X(_0493_));
 sg13g2_mux4_1 _1840_ (.S0(_0481_),
    .A0(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ),
    .A1(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ),
    .A2(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ),
    .A3(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ),
    .S1(_0487_),
    .X(_0494_));
 sg13g2_mux2_1 _1841_ (.A0(_0493_),
    .A1(_0494_),
    .S(_0486_),
    .X(_0495_));
 sg13g2_mux2_1 _1842_ (.A0(_0492_),
    .A1(_0495_),
    .S(_0473_),
    .X(_0496_));
 sg13g2_mux2_2 _1843_ (.A0(_0496_),
    .A1(\Inst_LF_LUT4c_frame_config_dffesr.LUT_flop ),
    .S(\Inst_LF_LUT4c_frame_config_dffesr.c_out_mux ),
    .X(F));
 sg13g2_o21ai_1 _1844_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit19.Q ),
    .Y(_0497_),
    .A1(net996),
    .A2(net933));
 sg13g2_a21oi_2 _1845_ (.B1(_0497_),
    .Y(_0498_),
    .A2(\Inst_LUT4AB_switch_matrix.M_AH ),
    .A1(net996));
 sg13g2_mux2_1 _1846_ (.A0(net965),
    .A1(net959),
    .S(net996),
    .X(_0499_));
 sg13g2_o21ai_1 _1847_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit20.Q ),
    .Y(_0500_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit19.Q ),
    .A2(_0499_));
 sg13g2_or2_1 _1848_ (.X(_0501_),
    .B(_0498_),
    .A(_0500_));
 sg13g2_nand2b_1 _1849_ (.Y(_0502_),
    .B(net996),
    .A_N(net947));
 sg13g2_o21ai_1 _1850_ (.B1(_0502_),
    .Y(_0503_),
    .A1(net996),
    .A2(net942));
 sg13g2_mux2_1 _1851_ (.A0(net976),
    .A1(net972),
    .S(net996),
    .X(_0504_));
 sg13g2_a21oi_1 _1852_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit19.Q ),
    .A2(_0503_),
    .Y(_0505_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit20.Q ));
 sg13g2_o21ai_1 _1853_ (.B1(_0505_),
    .Y(_0506_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit19.Q ),
    .A2(_0504_));
 sg13g2_and2_1 _1854_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit21.Q ),
    .B(_0506_),
    .X(_0507_));
 sg13g2_mux4_1 _1855_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit18.Q ),
    .A0(net34),
    .A1(net42),
    .A2(net5),
    .A3(net13),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit19.Q ),
    .X(_0508_));
 sg13g2_nand2b_1 _1856_ (.Y(_0509_),
    .B(_0508_),
    .A_N(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit20.Q ));
 sg13g2_nand2b_1 _1857_ (.Y(_0510_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit18.Q ),
    .A_N(net89));
 sg13g2_o21ai_1 _1858_ (.B1(_0510_),
    .Y(_0511_),
    .A1(net996),
    .A2(net1006));
 sg13g2_mux2_1 _1859_ (.A0(net62),
    .A1(net70),
    .S(net996),
    .X(_0512_));
 sg13g2_o21ai_1 _1860_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit20.Q ),
    .Y(_0513_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit19.Q ),
    .A2(_0512_));
 sg13g2_a21oi_1 _1861_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit19.Q ),
    .A2(_0511_),
    .Y(_0514_),
    .B1(_0513_));
 sg13g2_nor2_1 _1862_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit21.Q ),
    .B(_0514_),
    .Y(_0515_));
 sg13g2_a22oi_1 _1863_ (.Y(\Inst_LUT4AB_switch_matrix.JN2BEG6 ),
    .B1(_0509_),
    .B2(_0515_),
    .A2(_0507_),
    .A1(_0501_));
 sg13g2_nor2b_1 _1864_ (.A(\Inst_LUT4AB_switch_matrix.JN2BEG6 ),
    .B_N(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit18.Q ),
    .Y(_0516_));
 sg13g2_nor2_1 _1865_ (.A(net77),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit18.Q ),
    .Y(_0517_));
 sg13g2_o21ai_1 _1866_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit19.Q ),
    .Y(_0518_),
    .A1(_0517_),
    .A2(_0516_));
 sg13g2_mux2_1 _1867_ (.A0(net49),
    .A1(net20),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit18.Q ),
    .X(_0519_));
 sg13g2_o21ai_1 _1868_ (.B1(_0518_),
    .Y(_0520_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit19.Q ),
    .A2(_0519_));
 sg13g2_mux2_1 _1869_ (.A0(net50),
    .A1(net21),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit18.Q ),
    .X(_0521_));
 sg13g2_nand2b_1 _1870_ (.Y(_0522_),
    .B(net78),
    .A_N(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit18.Q ));
 sg13g2_nand2_1 _1871_ (.Y(_0523_),
    .A(net105),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit18.Q ));
 sg13g2_nand3_1 _1872_ (.B(_0522_),
    .C(_0523_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit19.Q ),
    .Y(_0524_));
 sg13g2_o21ai_1 _1873_ (.B1(_0524_),
    .Y(_0525_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit19.Q ),
    .A2(_0521_));
 sg13g2_mux4_1 _1874_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit18.Q ),
    .A0(net54),
    .A1(net22),
    .A2(net82),
    .A3(\Inst_LUT4AB_switch_matrix.JN2BEG4 ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit19.Q ),
    .X(_0526_));
 sg13g2_inv_1 _1875_ (.Y(_0527_),
    .A(_0526_));
 sg13g2_mux4_1 _1876_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit18.Q ),
    .A0(net42),
    .A1(net13),
    .A2(net70),
    .A3(net108),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit19.Q ),
    .X(_0528_));
 sg13g2_inv_1 _1877_ (.Y(_0529_),
    .A(_0528_));
 sg13g2_mux4_1 _1878_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit31.Q ),
    .A0(_0520_),
    .A1(_0525_),
    .A2(_0529_),
    .A3(_0527_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit0.Q ),
    .X(_0530_));
 sg13g2_a21oi_1 _1879_ (.A1(net386),
    .A2(_0490_),
    .Y(_0531_),
    .B1(_0488_));
 sg13g2_mux2_1 _1880_ (.A0(_0530_),
    .A1(_0531_),
    .S(\Inst_LG_LUT4c_frame_config_dffesr.c_I0mux ),
    .X(_0532_));
 sg13g2_mux2_1 _1881_ (.A0(net1211),
    .A1(net80),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit22.Q ),
    .X(_0533_));
 sg13g2_nand2_1 _1882_ (.Y(_0534_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit22.Q ),
    .B(net380));
 sg13g2_nand2b_1 _1883_ (.Y(_0535_),
    .B(net111),
    .A_N(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit22.Q ));
 sg13g2_nand3_1 _1884_ (.B(_0534_),
    .C(_0535_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit23.Q ),
    .Y(_0536_));
 sg13g2_o21ai_1 _1885_ (.B1(_0536_),
    .Y(_0537_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit23.Q ),
    .A2(_0533_));
 sg13g2_mux4_1 _1886_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit23.Q ),
    .A0(net56),
    .A1(net68),
    .A2(net11),
    .A3(net95),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit22.Q ),
    .X(_0538_));
 sg13g2_mux4_1 _1887_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit18.Q ),
    .A0(net976),
    .A1(net971),
    .A2(net941),
    .A3(net946),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit19.Q ),
    .X(_0539_));
 sg13g2_mux2_1 _1888_ (.A0(net965),
    .A1(net958),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit18.Q ),
    .X(_0540_));
 sg13g2_o21ai_1 _1889_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit19.Q ),
    .Y(_0541_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit18.Q ),
    .A2(net933));
 sg13g2_a21oi_1 _1890_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit18.Q ),
    .A2(\Inst_LUT4AB_switch_matrix.M_AB ),
    .Y(_0542_),
    .B1(_0541_));
 sg13g2_o21ai_1 _1891_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit20.Q ),
    .Y(_0543_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit19.Q ),
    .A2(_0540_));
 sg13g2_o21ai_1 _1892_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit21.Q ),
    .Y(_0544_),
    .A1(_0542_),
    .A2(_0543_));
 sg13g2_a21oi_1 _1893_ (.A1(_1044_),
    .A2(_0539_),
    .Y(_0545_),
    .B1(_0544_));
 sg13g2_mux4_1 _1894_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit18.Q ),
    .A0(net34),
    .A1(net42),
    .A2(net5),
    .A3(net13),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit19.Q ),
    .X(_0546_));
 sg13g2_nand2b_1 _1895_ (.Y(_0547_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit18.Q ),
    .A_N(net1003));
 sg13g2_o21ai_1 _1896_ (.B1(_0547_),
    .Y(_0548_),
    .A1(net1006),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit18.Q ));
 sg13g2_mux2_1 _1897_ (.A0(net62),
    .A1(net70),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit18.Q ),
    .X(_0549_));
 sg13g2_or2_1 _1898_ (.X(_0550_),
    .B(_0549_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit19.Q ));
 sg13g2_a21oi_1 _1899_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit19.Q ),
    .A2(_0548_),
    .Y(_0551_),
    .B1(_1044_));
 sg13g2_a221oi_1 _1900_ (.B2(_0551_),
    .C1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit21.Q ),
    .B1(_0550_),
    .A1(_1044_),
    .Y(_0552_),
    .A2(_0546_));
 sg13g2_nor2_2 _1901_ (.A(_0545_),
    .B(_0552_),
    .Y(\Inst_LUT4AB_switch_matrix.JS2BEG6 ));
 sg13g2_o21ai_1 _1902_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit23.Q ),
    .Y(_0553_),
    .A1(_1026_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit22.Q ));
 sg13g2_a21o_1 _1903_ (.A2(\Inst_LUT4AB_switch_matrix.JS2BEG6 ),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit22.Q ),
    .B1(_0553_),
    .X(_0554_));
 sg13g2_mux2_1 _1904_ (.A0(net18),
    .A1(net75),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit22.Q ),
    .X(_0555_));
 sg13g2_o21ai_1 _1905_ (.B1(_0554_),
    .Y(_0556_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit23.Q ),
    .A2(_0555_));
 sg13g2_mux2_1 _1906_ (.A0(net48),
    .A1(net19),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit22.Q ),
    .X(_0557_));
 sg13g2_nand2b_1 _1907_ (.Y(_0558_),
    .B(net76),
    .A_N(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit22.Q ));
 sg13g2_nand2_1 _1908_ (.Y(_0559_),
    .A(net103),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit22.Q ));
 sg13g2_nand3_1 _1909_ (.B(_0558_),
    .C(_0559_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit23.Q ),
    .Y(_0560_));
 sg13g2_o21ai_1 _1910_ (.B1(_0560_),
    .Y(_0561_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit23.Q ),
    .A2(_0557_));
 sg13g2_mux2_1 _1911_ (.A0(_0556_),
    .A1(_0561_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit3.Q ),
    .X(_0562_));
 sg13g2_o21ai_1 _1912_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit4.Q ),
    .Y(_0563_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit3.Q ),
    .A2(_0538_));
 sg13g2_a21o_1 _1913_ (.A2(_0537_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit3.Q ),
    .B1(_0563_),
    .X(_0564_));
 sg13g2_o21ai_1 _1914_ (.B1(_0564_),
    .Y(_0565_),
    .A1(_0562_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit4.Q ));
 sg13g2_mux4_1 _1915_ (.S0(net992),
    .A0(net978),
    .A1(net973),
    .A2(net943),
    .A3(D),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit19.Q ),
    .X(_0566_));
 sg13g2_nand2b_1 _1916_ (.Y(_0567_),
    .B(_0566_),
    .A_N(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit20.Q ));
 sg13g2_mux2_1 _1917_ (.A0(net966),
    .A1(net960),
    .S(net992),
    .X(_0568_));
 sg13g2_nand2b_1 _1918_ (.Y(_0569_),
    .B(net992),
    .A_N(net931));
 sg13g2_o21ai_1 _1919_ (.B1(_0569_),
    .Y(_0570_),
    .A1(net992),
    .A2(net936));
 sg13g2_o21ai_1 _1920_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit20.Q ),
    .Y(_0571_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit19.Q ),
    .A2(_0568_));
 sg13g2_a21oi_1 _1921_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit19.Q ),
    .A2(_0570_),
    .Y(_0572_),
    .B1(_0571_));
 sg13g2_nor2b_1 _1922_ (.A(_0572_),
    .B_N(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit21.Q ),
    .Y(_0573_));
 sg13g2_nand2b_1 _1923_ (.Y(_0574_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit18.Q ),
    .A_N(net13));
 sg13g2_o21ai_1 _1924_ (.B1(_0574_),
    .Y(_0575_),
    .A1(net5),
    .A2(net992));
 sg13g2_mux2_1 _1925_ (.A0(net1007),
    .A1(net42),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit18.Q ),
    .X(_0576_));
 sg13g2_a21oi_1 _1926_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit19.Q ),
    .A2(_0575_),
    .Y(_0577_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit20.Q ));
 sg13g2_o21ai_1 _1927_ (.B1(_0577_),
    .Y(_0578_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit19.Q ),
    .A2(_0576_));
 sg13g2_nand2b_1 _1928_ (.Y(_0579_),
    .B(net992),
    .A_N(net1003));
 sg13g2_o21ai_1 _1929_ (.B1(_0579_),
    .Y(_0580_),
    .A1(net70),
    .A2(net992));
 sg13g2_mux2_1 _1930_ (.A0(net60),
    .A1(net62),
    .S(net992),
    .X(_0581_));
 sg13g2_o21ai_1 _1931_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit20.Q ),
    .Y(_0582_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit19.Q ),
    .A2(_0581_));
 sg13g2_a21oi_1 _1932_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit19.Q ),
    .A2(_0580_),
    .Y(_0583_),
    .B1(_0582_));
 sg13g2_nor2_1 _1933_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit21.Q ),
    .B(_0583_),
    .Y(_0584_));
 sg13g2_a22oi_1 _1934_ (.Y(\Inst_LUT4AB_switch_matrix.E2BEG6 ),
    .B1(_0578_),
    .B2(_0584_),
    .A2(_0573_),
    .A1(_0567_));
 sg13g2_mux4_1 _1935_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit21.Q ),
    .A0(net45),
    .A1(net100),
    .A2(net73),
    .A3(\Inst_LUT4AB_switch_matrix.E2BEG6 ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit20.Q ),
    .X(_0585_));
 sg13g2_mux4_1 _1936_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit20.Q ),
    .A0(net46),
    .A1(net17),
    .A2(net74),
    .A3(net101),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit21.Q ),
    .X(_0586_));
 sg13g2_mux4_1 _1937_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit21.Q ),
    .A0(net53),
    .A1(net92),
    .A2(net85),
    .A3(\Inst_LUT4AB_switch_matrix.E2BEG4 ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit20.Q ),
    .X(_0587_));
 sg13g2_mux4_1 _1938_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit21.Q ),
    .A0(net38),
    .A1(net83),
    .A2(net9),
    .A3(net93),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit20.Q ),
    .X(_0588_));
 sg13g2_inv_1 _1939_ (.Y(_0589_),
    .A(_0588_));
 sg13g2_mux4_1 _1940_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit1.Q ),
    .A0(_0585_),
    .A1(net981),
    .A2(_0588_),
    .A3(_0587_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit2.Q ),
    .X(_0590_));
 sg13g2_nor2_2 _1941_ (.A(_0590_),
    .B(_0565_),
    .Y(_0591_));
 sg13g2_mux4_1 _1942_ (.S0(net378),
    .A0(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ),
    .A1(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ),
    .A2(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ),
    .A3(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ),
    .S1(net374),
    .X(_0592_));
 sg13g2_inv_1 _1943_ (.Y(_0593_),
    .A(_0592_));
 sg13g2_o21ai_1 _1944_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit19.Q ),
    .Y(_0594_),
    .A1(net983),
    .A2(net933));
 sg13g2_a21oi_2 _1945_ (.B1(_0594_),
    .Y(_0595_),
    .A2(\Inst_LUT4AB_switch_matrix.M_EF ),
    .A1(net983));
 sg13g2_mux2_1 _1946_ (.A0(net965),
    .A1(net958),
    .S(net983),
    .X(_0596_));
 sg13g2_o21ai_1 _1947_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit20.Q ),
    .Y(_0597_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit19.Q ),
    .A2(_0596_));
 sg13g2_or2_1 _1948_ (.X(_0598_),
    .B(_0595_),
    .A(_0597_));
 sg13g2_nand2b_1 _1949_ (.Y(_0599_),
    .B(net983),
    .A_N(net946));
 sg13g2_o21ai_1 _1950_ (.B1(_0599_),
    .Y(_0600_),
    .A1(net983),
    .A2(net941));
 sg13g2_mux2_1 _1951_ (.A0(net976),
    .A1(net971),
    .S(net983),
    .X(_0601_));
 sg13g2_a21oi_1 _1952_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit19.Q ),
    .A2(_0600_),
    .Y(_0602_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit20.Q ));
 sg13g2_o21ai_1 _1953_ (.B1(_0602_),
    .Y(_0603_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit19.Q ),
    .A2(_0601_));
 sg13g2_and2_1 _1954_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit21.Q ),
    .B(_0603_),
    .X(_0604_));
 sg13g2_mux2_1 _1955_ (.A0(net60),
    .A1(net62),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit18.Q ),
    .X(_0605_));
 sg13g2_nand2b_1 _1956_ (.Y(_0606_),
    .B(net983),
    .A_N(net1003));
 sg13g2_o21ai_1 _1957_ (.B1(_0606_),
    .Y(_0607_),
    .A1(net70),
    .A2(net983));
 sg13g2_o21ai_1 _1958_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit20.Q ),
    .Y(_0608_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit19.Q ),
    .A2(_0605_));
 sg13g2_a21oi_1 _1959_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit19.Q ),
    .A2(_0607_),
    .Y(_0609_),
    .B1(_0608_));
 sg13g2_mux4_1 _1960_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit18.Q ),
    .A0(net1007),
    .A1(net42),
    .A2(net1214),
    .A3(net13),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit19.Q ),
    .X(_0610_));
 sg13g2_nand2b_1 _1961_ (.Y(_0611_),
    .B(_0610_),
    .A_N(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit20.Q ));
 sg13g2_nor2_1 _1962_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit21.Q ),
    .B(_0609_),
    .Y(_0612_));
 sg13g2_a22oi_1 _1963_ (.Y(\Inst_LUT4AB_switch_matrix.JW2BEG6 ),
    .B1(_0611_),
    .B2(_0612_),
    .A2(_0604_),
    .A1(_0598_));
 sg13g2_nor2b_1 _1964_ (.A(\Inst_LUT4AB_switch_matrix.JW2BEG6 ),
    .B_N(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit24.Q ),
    .Y(_0613_));
 sg13g2_nor2_1 _1965_ (.A(net98),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit24.Q ),
    .Y(_0614_));
 sg13g2_o21ai_1 _1966_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit25.Q ),
    .Y(_0615_),
    .A1(_0614_),
    .A2(_0613_));
 sg13g2_mux2_1 _1967_ (.A0(net43),
    .A1(net14),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit24.Q ),
    .X(_0616_));
 sg13g2_o21ai_1 _1968_ (.B1(_0615_),
    .Y(_0617_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit25.Q ),
    .A2(_0616_));
 sg13g2_mux2_1 _1969_ (.A0(net44),
    .A1(net15),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit24.Q ),
    .X(_0618_));
 sg13g2_nand2b_1 _1970_ (.Y(_0619_),
    .B(net72),
    .A_N(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit24.Q ));
 sg13g2_nand2_1 _1971_ (.Y(_0620_),
    .A(net99),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit24.Q ));
 sg13g2_nand3_1 _1972_ (.B(_0619_),
    .C(_0620_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit25.Q ),
    .Y(_0621_));
 sg13g2_o21ai_1 _1973_ (.B1(_0621_),
    .Y(_0622_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit25.Q ),
    .A2(_0618_));
 sg13g2_mux4_1 _1974_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit25.Q ),
    .A0(net55),
    .A1(net90),
    .A2(net1213),
    .A3(\Inst_LUT4AB_switch_matrix.JW2BEG4 ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit24.Q ),
    .X(_0623_));
 sg13g2_inv_1 _1975_ (.Y(_0624_),
    .A(_0623_));
 sg13g2_mux4_1 _1976_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit25.Q ),
    .A0(net36),
    .A1(net64),
    .A2(net25),
    .A3(net91),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit24.Q ),
    .X(_0625_));
 sg13g2_inv_1 _1977_ (.Y(_0626_),
    .A(_0625_));
 sg13g2_mux4_1 _1978_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit5.Q ),
    .A0(_0617_),
    .A1(_0622_),
    .A2(_0626_),
    .A3(_0624_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit6.Q ),
    .X(_0627_));
 sg13g2_mux4_1 _1979_ (.S0(net378),
    .A0(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ),
    .A1(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ),
    .A2(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ),
    .A3(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ),
    .S1(_0565_),
    .X(_0628_));
 sg13g2_o21ai_1 _1980_ (.B1(_0627_),
    .Y(_0629_),
    .A1(_0628_),
    .A2(_0532_));
 sg13g2_a21oi_2 _1981_ (.B1(_0629_),
    .Y(_0630_),
    .A2(_0593_),
    .A1(_0532_));
 sg13g2_mux4_1 _1982_ (.S0(net378),
    .A0(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ),
    .A1(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ),
    .A2(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ),
    .A3(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ),
    .S1(net374),
    .X(_0631_));
 sg13g2_nand2b_1 _1983_ (.Y(_0632_),
    .B(_0532_),
    .A_N(_0631_));
 sg13g2_mux4_1 _1984_ (.S0(net378),
    .A0(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ),
    .A1(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ),
    .A2(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ),
    .A3(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ),
    .S1(net374),
    .X(_0633_));
 sg13g2_nor2_1 _1985_ (.A(_0532_),
    .B(_0633_),
    .Y(_0634_));
 sg13g2_nor2_1 _1986_ (.A(_0627_),
    .B(_0634_),
    .Y(_0635_));
 sg13g2_a21oi_2 _1987_ (.B1(_0630_),
    .Y(_0636_),
    .A2(_0635_),
    .A1(_0632_));
 sg13g2_nand2_1 _1988_ (.Y(_0637_),
    .A(\Inst_LG_LUT4c_frame_config_dffesr.LUT_flop ),
    .B(\Inst_LG_LUT4c_frame_config_dffesr.c_out_mux ));
 sg13g2_o21ai_1 _1989_ (.B1(_0637_),
    .Y(G),
    .A1(_0636_),
    .A2(\Inst_LG_LUT4c_frame_config_dffesr.c_out_mux ));
 sg13g2_a221oi_1 _1990_ (.B2(net378),
    .C1(_0488_),
    .B1(net374),
    .A1(net386),
    .Y(_0638_),
    .A2(_0490_));
 sg13g2_or2_1 _1991_ (.X(_0639_),
    .B(net387),
    .A(_0591_));
 sg13g2_o21ai_1 _1992_ (.B1(\Inst_LH_LUT4c_frame_config_dffesr.c_I0mux ),
    .Y(_0640_),
    .A1(_0638_),
    .A2(_0591_));
 sg13g2_o21ai_1 _1993_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit10.Q ),
    .Y(_0641_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit9.Q ),
    .A2(_0528_));
 sg13g2_a21oi_1 _1994_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit9.Q ),
    .A2(_0527_),
    .Y(_0642_),
    .B1(_0641_));
 sg13g2_mux2_1 _1995_ (.A0(_0520_),
    .A1(_0525_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit9.Q ),
    .X(_0643_));
 sg13g2_nor2_1 _1996_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit10.Q ),
    .B(_0643_),
    .Y(_0644_));
 sg13g2_or3_1 _1997_ (.A(\Inst_LH_LUT4c_frame_config_dffesr.c_I0mux ),
    .B(_0642_),
    .C(_0644_),
    .X(_0645_));
 sg13g2_mux2_1 _1998_ (.A0(_0556_),
    .A1(_0561_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit13.Q ),
    .X(_0646_));
 sg13g2_o21ai_1 _1999_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit14.Q ),
    .Y(_0647_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit13.Q ),
    .A2(_0538_));
 sg13g2_a21o_1 _2000_ (.A2(_0537_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit13.Q ),
    .B1(_0647_),
    .X(_0648_));
 sg13g2_o21ai_1 _2001_ (.B1(_0648_),
    .Y(_0649_),
    .A1(_0646_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit14.Q ));
 sg13g2_mux4_1 _2002_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit11.Q ),
    .A0(_0585_),
    .A1(net981),
    .A2(_0588_),
    .A3(_0587_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit12.Q ),
    .X(_0650_));
 sg13g2_nand2_1 _2003_ (.Y(_0651_),
    .A(_0649_),
    .B(_0650_));
 sg13g2_nor2_2 _2004_ (.A(_0649_),
    .B(_0650_),
    .Y(_0652_));
 sg13g2_mux4_1 _2005_ (.S0(_0650_),
    .A0(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ),
    .A1(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ),
    .A2(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ),
    .A3(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ),
    .S1(net379),
    .X(_0653_));
 sg13g2_a21o_1 _2006_ (.A2(_0645_),
    .A1(net388),
    .B1(_0653_),
    .X(_0654_));
 sg13g2_mux4_1 _2007_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit15.Q ),
    .A0(_0617_),
    .A1(_0622_),
    .A2(_0626_),
    .A3(_0624_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit16.Q ),
    .X(_0655_));
 sg13g2_mux4_1 _2008_ (.S0(_0650_),
    .A0(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ),
    .A1(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ),
    .A2(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ),
    .A3(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ),
    .S1(_0649_),
    .X(_0656_));
 sg13g2_inv_1 _2009_ (.Y(_0657_),
    .A(_0656_));
 sg13g2_nand3_1 _2010_ (.B(_0645_),
    .C(_0657_),
    .A(net381),
    .Y(_0658_));
 sg13g2_and3_1 _2011_ (.X(_0659_),
    .A(_0654_),
    .B(_0655_),
    .C(_0658_));
 sg13g2_mux4_1 _2012_ (.S0(_0650_),
    .A0(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ),
    .A1(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ),
    .A2(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ),
    .A3(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ),
    .S1(_0649_),
    .X(_0660_));
 sg13g2_a21o_1 _2013_ (.A2(_0645_),
    .A1(net381),
    .B1(_0660_),
    .X(_0661_));
 sg13g2_mux4_1 _2014_ (.S0(_0650_),
    .A0(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ),
    .A1(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ),
    .A2(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ),
    .A3(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ),
    .S1(net379),
    .X(_0662_));
 sg13g2_inv_1 _2015_ (.Y(_0663_),
    .A(_0662_));
 sg13g2_nand3_1 _2016_ (.B(_0645_),
    .C(_0663_),
    .A(net381),
    .Y(_0664_));
 sg13g2_nor2b_1 _2017_ (.A(_0655_),
    .B_N(_0664_),
    .Y(_0665_));
 sg13g2_a21oi_2 _2018_ (.B1(_0659_),
    .Y(_0666_),
    .A2(_0665_),
    .A1(_0661_));
 sg13g2_nand2_1 _2019_ (.Y(_0667_),
    .A(\Inst_LH_LUT4c_frame_config_dffesr.LUT_flop ),
    .B(\Inst_LH_LUT4c_frame_config_dffesr.c_out_mux ));
 sg13g2_o21ai_1 _2020_ (.B1(_0667_),
    .Y(H),
    .A1(_0666_),
    .A2(\Inst_LH_LUT4c_frame_config_dffesr.c_out_mux ));
 sg13g2_mux4_1 _2021_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit23.Q ),
    .A0(\Inst_LUT4AB_switch_matrix.JN2BEG6 ),
    .A1(\Inst_LUT4AB_switch_matrix.JS2BEG6 ),
    .A2(\Inst_LUT4AB_switch_matrix.E2BEG6 ),
    .A3(\Inst_LUT4AB_switch_matrix.JW2BEG6 ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit22.Q ),
    .X(_0668_));
 sg13g2_mux4_1 _2022_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit19.Q ),
    .A0(\Inst_LUT4AB_switch_matrix.JN2BEG4 ),
    .A1(\Inst_LUT4AB_switch_matrix.JS2BEG4 ),
    .A2(\Inst_LUT4AB_switch_matrix.E2BEG4 ),
    .A3(\Inst_LUT4AB_switch_matrix.JW2BEG4 ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit18.Q ),
    .X(_0669_));
 sg13g2_mux2_1 _2023_ (.A0(_0668_),
    .A1(_0669_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit17.Q ),
    .X(_0670_));
 sg13g2_mux2_2 _2024_ (.A0(net965),
    .A1(net958),
    .S(_0670_),
    .X(\Inst_LUT4AB_switch_matrix.M_EF ));
 sg13g2_o21ai_1 _2025_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit2.Q ),
    .Y(_0671_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit1.Q ),
    .A2(_0366_));
 sg13g2_a21o_1 _2026_ (.A2(_0365_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit1.Q ),
    .B1(_0671_),
    .X(_0672_));
 sg13g2_a21oi_1 _2027_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit1.Q ),
    .A2(_0391_),
    .Y(_0673_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit2.Q ));
 sg13g2_o21ai_1 _2028_ (.B1(_0673_),
    .Y(_0674_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit1.Q ),
    .A2(_0389_));
 sg13g2_nor2b_1 _2029_ (.A(\Inst_LD_LUT4c_frame_config_dffesr.c_I0mux ),
    .B_N(_0674_),
    .Y(_0675_));
 sg13g2_a22oi_1 _2030_ (.Y(_0676_),
    .B1(_0672_),
    .B2(_0675_),
    .A2(_0208_),
    .A1(\Inst_LD_LUT4c_frame_config_dffesr.c_I0mux ));
 sg13g2_mux4_1 _2031_ (.S0(_0149_),
    .A0(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ),
    .A1(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ),
    .A2(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ),
    .A3(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ),
    .S1(_0199_),
    .X(_0677_));
 sg13g2_nor2_1 _2032_ (.A(_0676_),
    .B(_0677_),
    .Y(_0678_));
 sg13g2_mux4_1 _2033_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit7.Q ),
    .A0(_0452_),
    .A1(_0454_),
    .A2(_0430_),
    .A3(_0424_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit8.Q ),
    .X(_0679_));
 sg13g2_mux4_1 _2034_ (.S0(_0149_),
    .A0(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ),
    .A1(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ),
    .A2(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ),
    .A3(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ),
    .S1(_0199_),
    .X(_0680_));
 sg13g2_nor2b_1 _2035_ (.A(_0680_),
    .B_N(_0676_),
    .Y(_0681_));
 sg13g2_nor3_2 _2036_ (.A(_0678_),
    .B(_0681_),
    .C(_0679_),
    .Y(_0682_));
 sg13g2_mux4_1 _2037_ (.S0(_0149_),
    .A0(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ),
    .A1(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ),
    .A2(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ),
    .A3(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ),
    .S1(_0199_),
    .X(_0683_));
 sg13g2_or2_1 _2038_ (.X(_0684_),
    .B(_0683_),
    .A(_0676_));
 sg13g2_mux4_1 _2039_ (.S0(_0149_),
    .A0(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ),
    .A1(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ),
    .A2(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ),
    .A3(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ),
    .S1(_0199_),
    .X(_0685_));
 sg13g2_nand2b_1 _2040_ (.Y(_0686_),
    .B(_0676_),
    .A_N(_0685_));
 sg13g2_and2_1 _2041_ (.A(_0679_),
    .B(_0686_),
    .X(_0687_));
 sg13g2_a21o_1 _2042_ (.A2(_0687_),
    .A1(_0684_),
    .B1(_0682_),
    .X(_0688_));
 sg13g2_mux2_2 _2043_ (.A0(_0688_),
    .A1(\Inst_LD_LUT4c_frame_config_dffesr.LUT_flop ),
    .S(\Inst_LD_LUT4c_frame_config_dffesr.c_out_mux ),
    .X(D));
 sg13g2_a21oi_1 _2044_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit20.Q ),
    .A2(\Inst_LUT4AB_switch_matrix.E2BEG5 ),
    .Y(_0689_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit21.Q ));
 sg13g2_o21ai_1 _2045_ (.B1(_0689_),
    .Y(_0690_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit20.Q ),
    .A2(_0230_));
 sg13g2_a21oi_2 _2046_ (.B1(_1047_),
    .Y(_0691_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit20.Q ),
    .A1(\Inst_LUT4AB_switch_matrix.JW2BEG5 ));
 sg13g2_o21ai_1 _2047_ (.B1(_0691_),
    .Y(_0692_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit20.Q ),
    .A2(_0275_));
 sg13g2_nand2_2 _2048_ (.Y(_0693_),
    .A(_0692_),
    .B(_0690_));
 sg13g2_nand2_1 _2049_ (.Y(_0694_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit16.Q ),
    .B(_0669_));
 sg13g2_o21ai_1 _2050_ (.B1(_0694_),
    .Y(_0695_),
    .A1(_0693_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit16.Q ));
 sg13g2_mux2_1 _2051_ (.A0(net942),
    .A1(net948),
    .S(_0695_),
    .X(_0696_));
 sg13g2_mux2_1 _2052_ (.A0(_0696_),
    .A1(net930),
    .S(_0693_),
    .X(_0697_));
 sg13g2_mux2_1 _2053_ (.A0(_0696_),
    .A1(_0697_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit16.Q ),
    .X(\Inst_LUT4AB_switch_matrix.M_AD ));
 sg13g2_o21ai_1 _2054_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit23.Q ),
    .Y(_0698_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit22.Q ),
    .A2(_1051_));
 sg13g2_a21oi_1 _2055_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit22.Q ),
    .A2(net931),
    .Y(_0699_),
    .B1(_0698_));
 sg13g2_mux2_1 _2056_ (.A0(net963),
    .A1(net956),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit22.Q ),
    .X(_0700_));
 sg13g2_o21ai_1 _2057_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit24.Q ),
    .Y(_0701_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit23.Q ),
    .A2(_0700_));
 sg13g2_mux4_1 _2058_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit22.Q ),
    .A0(net974),
    .A1(net969),
    .A2(net939),
    .A3(net945),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit23.Q ),
    .X(_0702_));
 sg13g2_o21ai_1 _2059_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit25.Q ),
    .Y(_0703_),
    .A1(_0699_),
    .A2(_0701_));
 sg13g2_a21oi_1 _2060_ (.A1(_1045_),
    .A2(_0702_),
    .Y(_0704_),
    .B1(_0703_));
 sg13g2_mux4_1 _2061_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit22.Q ),
    .A0(net1010),
    .A1(net35),
    .A2(net1217),
    .A3(net6),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit23.Q ),
    .X(_0705_));
 sg13g2_nand2b_1 _2062_ (.Y(_0706_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit22.Q ),
    .A_N(net1004));
 sg13g2_o21ai_1 _2063_ (.B1(_0706_),
    .Y(_0707_),
    .A1(net87),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit22.Q ));
 sg13g2_mux2_1 _2064_ (.A0(net59),
    .A1(net63),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit22.Q ),
    .X(_0708_));
 sg13g2_o21ai_1 _2065_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit24.Q ),
    .Y(_0709_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit23.Q ),
    .A2(_0708_));
 sg13g2_a21oi_1 _2066_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit23.Q ),
    .A2(_0707_),
    .Y(_0710_),
    .B1(_0709_));
 sg13g2_a21oi_1 _2067_ (.A1(_1045_),
    .A2(_0705_),
    .Y(_0711_),
    .B1(_0710_));
 sg13g2_a21oi_1 _2068_ (.A1(_1046_),
    .A2(_0711_),
    .Y(\Inst_LUT4AB_switch_matrix.JS2BEG7 ),
    .B1(_0704_));
 sg13g2_mux4_1 _2069_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit23.Q ),
    .A0(net963),
    .A1(net951),
    .A2(net956),
    .A3(net930),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit22.Q ),
    .X(_0712_));
 sg13g2_mux4_1 _2070_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit22.Q ),
    .A0(net974),
    .A1(net969),
    .A2(net939),
    .A3(net945),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit23.Q ),
    .X(_0713_));
 sg13g2_nand2b_1 _2071_ (.Y(_0714_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit24.Q ),
    .A_N(_0712_));
 sg13g2_o21ai_1 _2072_ (.B1(_0714_),
    .Y(_0715_),
    .A1(_0713_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit24.Q ));
 sg13g2_mux4_1 _2073_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit22.Q ),
    .A0(net1010),
    .A1(net55),
    .A2(net1217),
    .A3(net6),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit23.Q ),
    .X(_0716_));
 sg13g2_nand2b_1 _2074_ (.Y(_0717_),
    .B(_0716_),
    .A_N(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit24.Q ));
 sg13g2_mux2_1 _2075_ (.A0(net59),
    .A1(net61),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit22.Q ),
    .X(_0718_));
 sg13g2_nand2b_1 _2076_ (.Y(_0719_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit22.Q ),
    .A_N(net87));
 sg13g2_o21ai_1 _2077_ (.B1(_0719_),
    .Y(_0720_),
    .A1(net63),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit22.Q ));
 sg13g2_o21ai_1 _2078_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit24.Q ),
    .Y(_0721_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit23.Q ),
    .A2(_0718_));
 sg13g2_a21oi_1 _2079_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit23.Q ),
    .A2(_0720_),
    .Y(_0722_),
    .B1(_0721_));
 sg13g2_nor2_1 _2080_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit25.Q ),
    .B(_0722_),
    .Y(_0723_));
 sg13g2_a22oi_1 _2081_ (.Y(\Inst_LUT4AB_switch_matrix.JW2BEG7 ),
    .B1(_0717_),
    .B2(_0723_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit25.Q ),
    .A1(_0715_));
 sg13g2_mux4_1 _2082_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit22.Q ),
    .A0(net977),
    .A1(net972),
    .A2(net942),
    .A3(net947),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit23.Q ),
    .X(_0724_));
 sg13g2_mux4_1 _2083_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit23.Q ),
    .A0(net966),
    .A1(net953),
    .A2(net959),
    .A3(net929),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit22.Q ),
    .X(_0725_));
 sg13g2_nand2b_1 _2084_ (.Y(_0726_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit24.Q ),
    .A_N(_0725_));
 sg13g2_o21ai_1 _2085_ (.B1(_0726_),
    .Y(_0727_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit24.Q ),
    .A2(_0724_));
 sg13g2_nand2b_1 _2086_ (.Y(_0728_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit22.Q ),
    .A_N(net1004));
 sg13g2_o21ai_1 _2087_ (.B1(_0728_),
    .Y(_0729_),
    .A1(net87),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit22.Q ));
 sg13g2_mux2_1 _2088_ (.A0(net59),
    .A1(net63),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit22.Q ),
    .X(_0730_));
 sg13g2_o21ai_1 _2089_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit24.Q ),
    .Y(_0731_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit23.Q ),
    .A2(_0730_));
 sg13g2_a21oi_1 _2090_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit23.Q ),
    .A2(_0729_),
    .Y(_0732_),
    .B1(_0731_));
 sg13g2_mux4_1 _2091_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit22.Q ),
    .A0(net1010),
    .A1(net35),
    .A2(net1217),
    .A3(net22),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit23.Q ),
    .X(_0733_));
 sg13g2_nand2b_1 _2092_ (.Y(_0734_),
    .B(_0733_),
    .A_N(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit24.Q ));
 sg13g2_nor2_1 _2093_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit25.Q ),
    .B(_0732_),
    .Y(_0735_));
 sg13g2_a22oi_1 _2094_ (.Y(\Inst_LUT4AB_switch_matrix.JN2BEG7 ),
    .B1(_0734_),
    .B2(_0735_),
    .A2(_0727_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit25.Q ));
 sg13g2_mux4_1 _2095_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit22.Q ),
    .A0(net978),
    .A1(net973),
    .A2(net943),
    .A3(net948),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit23.Q ),
    .X(_0736_));
 sg13g2_mux4_1 _2096_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit23.Q ),
    .A0(net966),
    .A1(net954),
    .A2(net960),
    .A3(net928),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit22.Q ),
    .X(_0737_));
 sg13g2_nand2b_1 _2097_ (.Y(_0738_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit24.Q ),
    .A_N(_0737_));
 sg13g2_o21ai_1 _2098_ (.B1(_0738_),
    .Y(_0739_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit24.Q ),
    .A2(_0736_));
 sg13g2_mux4_1 _2099_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit22.Q ),
    .A0(net1010),
    .A1(net35),
    .A2(net1217),
    .A3(net6),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit23.Q ),
    .X(_0740_));
 sg13g2_nand2b_1 _2100_ (.Y(_0741_),
    .B(_0740_),
    .A_N(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit24.Q ));
 sg13g2_nand2b_1 _2101_ (.Y(_0742_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit22.Q ),
    .A_N(net108));
 sg13g2_o21ai_1 _2102_ (.B1(_0742_),
    .Y(_0743_),
    .A1(net83),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit22.Q ));
 sg13g2_mux2_1 _2103_ (.A0(net59),
    .A1(net61),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit22.Q ),
    .X(_0744_));
 sg13g2_o21ai_1 _2104_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit24.Q ),
    .Y(_0745_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit23.Q ),
    .A2(_0744_));
 sg13g2_a21oi_1 _2105_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit23.Q ),
    .A2(_0743_),
    .Y(_0746_),
    .B1(_0745_));
 sg13g2_nor2_1 _2106_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit25.Q ),
    .B(_0746_),
    .Y(_0747_));
 sg13g2_a22oi_1 _2107_ (.Y(\Inst_LUT4AB_switch_matrix.E2BEG7 ),
    .B1(_0741_),
    .B2(_0747_),
    .A2(_0739_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit25.Q ));
 sg13g2_mux2_1 _2108_ (.A0(\Inst_LUT4AB_switch_matrix.JN2BEG7 ),
    .A1(\Inst_LUT4AB_switch_matrix.E2BEG7 ),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit24.Q ),
    .X(_0748_));
 sg13g2_nand2_2 _2109_ (.Y(_0749_),
    .A(\Inst_LUT4AB_switch_matrix.JW2BEG7 ),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit24.Q ));
 sg13g2_nand2b_1 _2110_ (.Y(_0750_),
    .B(\Inst_LUT4AB_switch_matrix.JS2BEG7 ),
    .A_N(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit24.Q ));
 sg13g2_nand3_1 _2111_ (.B(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit25.Q ),
    .C(_0750_),
    .A(_0749_),
    .Y(_0751_));
 sg13g2_o21ai_1 _2112_ (.B1(_0751_),
    .Y(_0752_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit25.Q ),
    .A2(_0748_));
 sg13g2_mux2_1 _2113_ (.A0(_0752_),
    .A1(_0693_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit17.Q ),
    .X(_0753_));
 sg13g2_nand2_1 _2114_ (.Y(_0754_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit16.Q ),
    .B(_0670_));
 sg13g2_o21ai_1 _2115_ (.B1(_0754_),
    .Y(_0755_),
    .A1(_0753_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit16.Q ));
 sg13g2_nor2_2 _2116_ (.A(net954),
    .B(_0755_),
    .Y(_0756_));
 sg13g2_a21oi_2 _2117_ (.B1(_0756_),
    .Y(_0757_),
    .A2(_0755_),
    .A1(net932));
 sg13g2_mux2_1 _2118_ (.A0(_0757_),
    .A1(net929),
    .S(_0753_),
    .X(_0758_));
 sg13g2_nor2b_1 _2119_ (.A(_0758_),
    .B_N(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit16.Q ),
    .Y(_0759_));
 sg13g2_nor2_1 _2120_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit16.Q ),
    .B(_0757_),
    .Y(_0760_));
 sg13g2_nor3_2 _2121_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit17.Q ),
    .B(_0760_),
    .C(_0759_),
    .Y(_0761_));
 sg13g2_mux2_1 _2122_ (.A0(_0758_),
    .A1(_0697_),
    .S(_0752_),
    .X(_0762_));
 sg13g2_a21o_1 _2123_ (.A2(_0762_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit17.Q ),
    .B1(_0761_),
    .X(\Inst_LUT4AB_switch_matrix.M_AH ));
 sg13g2_mux2_2 _2124_ (.A0(net979),
    .A1(net972),
    .S(_0669_),
    .X(\Inst_LUT4AB_switch_matrix.M_AB ));
 sg13g2_mux4_1 _2125_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit27.Q ),
    .A0(net968),
    .A1(net944),
    .A2(net938),
    .A3(net961),
    .S1(net986),
    .X(_0763_));
 sg13g2_nor2b_1 _2126_ (.A(net986),
    .B_N(net955),
    .Y(_0764_));
 sg13g2_a21oi_1 _2127_ (.A1(net986),
    .A2(net950),
    .Y(_0765_),
    .B1(_0764_));
 sg13g2_nand2_1 _2128_ (.Y(_0766_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit26.Q ),
    .B(net931));
 sg13g2_o21ai_1 _2129_ (.B1(_0766_),
    .Y(_0767_),
    .A1(net986),
    .A2(net932));
 sg13g2_o21ai_1 _2130_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit28.Q ),
    .Y(_0768_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit27.Q ),
    .A2(_0765_));
 sg13g2_a21oi_1 _2131_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit27.Q ),
    .A2(_0767_),
    .Y(_0769_),
    .B1(_0768_));
 sg13g2_nor2b_1 _2132_ (.A(_0769_),
    .B_N(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit29.Q ),
    .Y(_0770_));
 sg13g2_o21ai_1 _2133_ (.B1(_0770_),
    .Y(_0771_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit28.Q ),
    .A2(_0763_));
 sg13g2_mux4_1 _2134_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit27.Q ),
    .A0(net1007),
    .A1(net7),
    .A2(net36),
    .A3(net1210),
    .S1(net986),
    .X(_0772_));
 sg13g2_mux2_1 _2135_ (.A0(net91),
    .A1(net107),
    .S(net986),
    .X(_0773_));
 sg13g2_nor2b_1 _2136_ (.A(net986),
    .B_N(net64),
    .Y(_0774_));
 sg13g2_a21oi_1 _2137_ (.A1(net80),
    .A2(net986),
    .Y(_0775_),
    .B1(_0774_));
 sg13g2_o21ai_1 _2138_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit28.Q ),
    .Y(_0776_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit27.Q ),
    .A2(_0775_));
 sg13g2_a21o_1 _2139_ (.A2(_0773_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit27.Q ),
    .B1(_0776_),
    .X(_0777_));
 sg13g2_o21ai_1 _2140_ (.B1(_0777_),
    .Y(_0778_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit28.Q ),
    .A2(_0772_));
 sg13g2_o21ai_1 _2141_ (.B1(_0771_),
    .Y(\Inst_LUT4AB_switch_matrix.JW2BEG0 ),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit29.Q ),
    .A2(_0778_));
 sg13g2_mux4_1 _2142_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit27.Q ),
    .A0(net969),
    .A1(net944),
    .A2(net938),
    .A3(net964),
    .S1(net991),
    .X(_0779_));
 sg13g2_nand2_1 _2143_ (.Y(_0780_),
    .A(net991),
    .B(net928));
 sg13g2_o21ai_1 _2144_ (.B1(_0780_),
    .Y(_0781_),
    .A1(net991),
    .A2(net932));
 sg13g2_nor2b_1 _2145_ (.A(net991),
    .B_N(net956),
    .Y(_0782_));
 sg13g2_a21oi_1 _2146_ (.A1(net991),
    .A2(net951),
    .Y(_0783_),
    .B1(_0782_));
 sg13g2_o21ai_1 _2147_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit28.Q ),
    .Y(_0784_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit27.Q ),
    .A2(_0783_));
 sg13g2_a21oi_1 _2148_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit27.Q ),
    .A2(_0781_),
    .Y(_0785_),
    .B1(_0784_));
 sg13g2_o21ai_1 _2149_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit29.Q ),
    .Y(_0786_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit28.Q ),
    .A2(_0779_));
 sg13g2_mux4_1 _2150_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit27.Q ),
    .A0(net56),
    .A1(net7),
    .A2(net1214),
    .A3(net1210),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit26.Q ),
    .X(_0787_));
 sg13g2_a21oi_1 _2151_ (.A1(_1036_),
    .A2(net991),
    .Y(_0788_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit27.Q ));
 sg13g2_o21ai_1 _2152_ (.B1(_0788_),
    .Y(_0789_),
    .A1(net64),
    .A2(net991));
 sg13g2_o21ai_1 _2153_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit27.Q ),
    .Y(_0790_),
    .A1(net91),
    .A2(net991));
 sg13g2_a21oi_1 _2154_ (.A1(_1028_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit26.Q ),
    .Y(_0791_),
    .B1(_0790_));
 sg13g2_nor2b_1 _2155_ (.A(_0791_),
    .B_N(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit28.Q ),
    .Y(_0792_));
 sg13g2_a21oi_1 _2156_ (.A1(_0789_),
    .A2(_0792_),
    .Y(_0793_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit29.Q ));
 sg13g2_o21ai_1 _2157_ (.B1(_0793_),
    .Y(_0794_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit28.Q ),
    .A2(_0787_));
 sg13g2_o21ai_1 _2158_ (.B1(_0794_),
    .Y(\Inst_LUT4AB_switch_matrix.JS2BEG0 ),
    .A1(_0785_),
    .A2(_0786_));
 sg13g2_nor2b_1 _2159_ (.A(net994),
    .B_N(net955),
    .Y(_0795_));
 sg13g2_a21oi_1 _2160_ (.A1(net994),
    .A2(net950),
    .Y(_0796_),
    .B1(_0795_));
 sg13g2_nand2_1 _2161_ (.Y(_0797_),
    .A(net995),
    .B(net929));
 sg13g2_o21ai_1 _2162_ (.B1(_0797_),
    .Y(_0798_),
    .A1(net995),
    .A2(net932));
 sg13g2_o21ai_1 _2163_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit28.Q ),
    .Y(_0799_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit27.Q ),
    .A2(_0796_));
 sg13g2_a21o_1 _2164_ (.A2(_0798_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit27.Q ),
    .B1(_0799_),
    .X(_0800_));
 sg13g2_mux2_1 _2165_ (.A0(net944),
    .A1(net961),
    .S(net994),
    .X(_0801_));
 sg13g2_nor2b_1 _2166_ (.A(net994),
    .B_N(net968),
    .Y(_0802_));
 sg13g2_a21oi_1 _2167_ (.A1(net994),
    .A2(net938),
    .Y(_0803_),
    .B1(_0802_));
 sg13g2_a21oi_1 _2168_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit27.Q ),
    .A2(_0801_),
    .Y(_0804_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit28.Q ));
 sg13g2_o21ai_1 _2169_ (.B1(_0804_),
    .Y(_0805_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit27.Q ),
    .A2(_0803_));
 sg13g2_nand3_1 _2170_ (.B(_0800_),
    .C(_0805_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit29.Q ),
    .Y(_0806_));
 sg13g2_mux2_1 _2171_ (.A0(net52),
    .A1(net23),
    .S(net995),
    .X(_0807_));
 sg13g2_nor2b_1 _2172_ (.A(net994),
    .B_N(net1007),
    .Y(_0808_));
 sg13g2_a21oi_1 _2173_ (.A1(net36),
    .A2(net994),
    .Y(_0809_),
    .B1(_0808_));
 sg13g2_a21oi_1 _2174_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit27.Q ),
    .A2(_0807_),
    .Y(_0810_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit28.Q ));
 sg13g2_o21ai_1 _2175_ (.B1(_0810_),
    .Y(_0811_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit27.Q ),
    .A2(_0809_));
 sg13g2_nor2b_1 _2176_ (.A(net995),
    .B_N(net1210),
    .Y(_0812_));
 sg13g2_a21oi_1 _2177_ (.A1(net64),
    .A2(net994),
    .Y(_0813_),
    .B1(_0812_));
 sg13g2_mux2_1 _2178_ (.A0(net91),
    .A1(net107),
    .S(net995),
    .X(_0814_));
 sg13g2_o21ai_1 _2179_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit28.Q ),
    .Y(_0815_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit27.Q ),
    .A2(_0813_));
 sg13g2_a21oi_1 _2180_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit27.Q ),
    .A2(_0814_),
    .Y(_0816_),
    .B1(_0815_));
 sg13g2_nand2b_1 _2181_ (.Y(_0817_),
    .B(_0811_),
    .A_N(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit29.Q ));
 sg13g2_o21ai_1 _2182_ (.B1(_0806_),
    .Y(\Inst_LUT4AB_switch_matrix.E2BEG0 ),
    .A1(_0816_),
    .A2(_0817_));
 sg13g2_mux4_1 _2183_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit27.Q ),
    .A0(net968),
    .A1(net944),
    .A2(net938),
    .A3(net961),
    .S1(net1001),
    .X(_0818_));
 sg13g2_nor2b_1 _2184_ (.A(net1001),
    .B_N(net956),
    .Y(_0819_));
 sg13g2_a21oi_1 _2185_ (.A1(net1001),
    .A2(net951),
    .Y(_0820_),
    .B1(_0819_));
 sg13g2_nand2_1 _2186_ (.Y(_0821_),
    .A(net1001),
    .B(net930));
 sg13g2_o21ai_1 _2187_ (.B1(_0821_),
    .Y(_0822_),
    .A1(net1001),
    .A2(net932));
 sg13g2_o21ai_1 _2188_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit28.Q ),
    .Y(_0823_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit27.Q ),
    .A2(_0820_));
 sg13g2_a21oi_1 _2189_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit27.Q ),
    .A2(_0822_),
    .Y(_0824_),
    .B1(_0823_));
 sg13g2_nor2b_1 _2190_ (.A(_0824_),
    .B_N(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit29.Q ),
    .Y(_0825_));
 sg13g2_o21ai_1 _2191_ (.B1(_0825_),
    .Y(_0826_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit28.Q ),
    .A2(_0818_));
 sg13g2_mux2_1 _2192_ (.A0(net1214),
    .A1(net7),
    .S(net1002),
    .X(_0827_));
 sg13g2_nor2b_1 _2193_ (.A(net1001),
    .B_N(net36),
    .Y(_0828_));
 sg13g2_a21oi_1 _2194_ (.A1(net52),
    .A2(net1001),
    .Y(_0829_),
    .B1(_0828_));
 sg13g2_a21oi_1 _2195_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit27.Q ),
    .A2(_0827_),
    .Y(_0830_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit28.Q ));
 sg13g2_o21ai_1 _2196_ (.B1(_0830_),
    .Y(_0831_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit27.Q ),
    .A2(_0829_));
 sg13g2_o21ai_1 _2197_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit27.Q ),
    .Y(_0832_),
    .A1(net91),
    .A2(net1001));
 sg13g2_a21oi_1 _2198_ (.A1(_1028_),
    .A2(net1002),
    .Y(_0833_),
    .B1(_0832_));
 sg13g2_nor2b_1 _2199_ (.A(net1002),
    .B_N(net1210),
    .Y(_0834_));
 sg13g2_a21oi_1 _2200_ (.A1(net84),
    .A2(net1002),
    .Y(_0835_),
    .B1(_0834_));
 sg13g2_o21ai_1 _2201_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit28.Q ),
    .Y(_0836_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit27.Q ),
    .A2(_0835_));
 sg13g2_o21ai_1 _2202_ (.B1(_0831_),
    .Y(_0837_),
    .A1(_0833_),
    .A2(_0836_));
 sg13g2_o21ai_1 _2203_ (.B1(_0826_),
    .Y(\Inst_LUT4AB_switch_matrix.JN2BEG0 ),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit29.Q ),
    .A2(_0837_));
 sg13g2_mux4_1 _2204_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit30.Q ),
    .A0(_1158_),
    .A1(_0196_),
    .A2(_0276_),
    .A3(_0556_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit31.Q ),
    .X(_0838_));
 sg13g2_mux4_1 _2205_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit30.Q ),
    .A0(net953),
    .A1(net935),
    .A2(net931),
    .A3(net929),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit31.Q ),
    .X(_0839_));
 sg13g2_o21ai_1 _2206_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit1.Q ),
    .Y(_0840_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit0.Q ),
    .A2(_0839_));
 sg13g2_a21oi_2 _2207_ (.B1(_0840_),
    .Y(_0841_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit0.Q ),
    .A1(_0838_));
 sg13g2_mux4_1 _2208_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit30.Q ),
    .A0(net1215),
    .A1(net1004),
    .A2(net974),
    .A3(net969),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit31.Q ),
    .X(_0842_));
 sg13g2_mux4_1 _2209_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit30.Q ),
    .A0(net939),
    .A1(net944),
    .A2(net963),
    .A3(net956),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit31.Q ),
    .X(_0843_));
 sg13g2_inv_1 _2210_ (.Y(_0844_),
    .A(_0843_));
 sg13g2_a21oi_1 _2211_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit0.Q ),
    .A2(_0844_),
    .Y(_0845_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit1.Q ));
 sg13g2_o21ai_1 _2212_ (.B1(_0845_),
    .Y(_0846_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit0.Q ),
    .A2(_0842_));
 sg13g2_nand2b_1 _2213_ (.Y(\Inst_LUT4AB_switch_matrix.W6BEG1 ),
    .B(_0846_),
    .A_N(_0841_));
 sg13g2_mux4_1 _2214_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit26.Q ),
    .A0(net1214),
    .A1(net1003),
    .A2(net977),
    .A3(net972),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit27.Q ),
    .X(_0847_));
 sg13g2_mux4_1 _2215_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit26.Q ),
    .A0(net942),
    .A1(net947),
    .A2(net966),
    .A3(net959),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit27.Q ),
    .X(_0848_));
 sg13g2_mux4_1 _2216_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit26.Q ),
    .A0(net953),
    .A1(net937),
    .A2(\Inst_LUT4AB_switch_matrix.M_AB ),
    .A3(\Inst_LUT4AB_switch_matrix.M_AH ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit27.Q ),
    .X(_0849_));
 sg13g2_mux4_1 _2217_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit26.Q ),
    .A0(_1084_),
    .A1(_0148_),
    .A2(_0308_),
    .A3(net981),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit27.Q ),
    .X(_0850_));
 sg13g2_mux4_1 _2218_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit28.Q ),
    .A0(_0847_),
    .A1(_0848_),
    .A2(_0849_),
    .A3(_0850_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit29.Q ),
    .X(\Inst_LUT4AB_switch_matrix.W6BEG0 ));
 sg13g2_mux2_1 _2219_ (.A0(net1009),
    .A1(net60),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit23.Q ),
    .X(_0851_));
 sg13g2_mux2_1 _2220_ (.A0(net1006),
    .A1(net945),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit23.Q ),
    .X(_0852_));
 sg13g2_nor2_1 _2221_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit23.Q ),
    .B(net966),
    .Y(_0853_));
 sg13g2_a21oi_2 _2222_ (.B1(_0853_),
    .Y(_0854_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit23.Q ),
    .A1(_0276_));
 sg13g2_nand2_1 _2223_ (.Y(_0855_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit23.Q ),
    .B(_1141_));
 sg13g2_o21ai_1 _2224_ (.B1(_0855_),
    .Y(_0856_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit23.Q ),
    .A2(_0556_));
 sg13g2_mux4_1 _2225_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit24.Q ),
    .A0(_0851_),
    .A1(_0852_),
    .A2(_0854_),
    .A3(_0856_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit25.Q ),
    .X(\Inst_LUT4AB_switch_matrix.WW4BEG3 ));
 sg13g2_o21ai_1 _2226_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit21.Q ),
    .Y(_0857_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit20.Q ),
    .A2(net980));
 sg13g2_a21oi_1 _2227_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit20.Q ),
    .A2(_0171_),
    .Y(_0858_),
    .B1(_0857_));
 sg13g2_nor2b_1 _2228_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit20.Q ),
    .B_N(net939),
    .Y(_0859_));
 sg13g2_a21oi_1 _2229_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit20.Q ),
    .A2(_0308_),
    .Y(_0860_),
    .B1(_0859_));
 sg13g2_o21ai_1 _2230_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit22.Q ),
    .Y(_0861_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit21.Q ),
    .A2(_0860_));
 sg13g2_nor2_1 _2231_ (.A(_0858_),
    .B(_0861_),
    .Y(_0862_));
 sg13g2_mux4_1 _2232_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit21.Q ),
    .A0(net1010),
    .A1(net87),
    .A2(net59),
    .A3(net969),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit20.Q ),
    .X(_0863_));
 sg13g2_nor2_1 _2233_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit22.Q ),
    .B(_0863_),
    .Y(_0864_));
 sg13g2_nor2_1 _2234_ (.A(_0862_),
    .B(_0864_),
    .Y(\Inst_LUT4AB_switch_matrix.WW4BEG2 ));
 sg13g2_mux4_1 _2235_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit17.Q ),
    .A0(net932),
    .A1(_1158_),
    .A2(_0196_),
    .A3(_0253_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit18.Q ),
    .X(_0865_));
 sg13g2_mux4_1 _2236_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit17.Q ),
    .A0(net1007),
    .A1(net62),
    .A2(net1003),
    .A3(net977),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit18.Q ),
    .X(_0866_));
 sg13g2_nand2_1 _2237_ (.Y(_0867_),
    .A(_1048_),
    .B(_0866_));
 sg13g2_o21ai_1 _2238_ (.B1(_0867_),
    .Y(\Inst_LUT4AB_switch_matrix.WW4BEG1 ),
    .A1(_1048_),
    .A2(_0865_));
 sg13g2_mux4_1 _2239_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit14.Q ),
    .A0(net33),
    .A1(net61),
    .A2(net1004),
    .A3(net959),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit15.Q ),
    .X(_0868_));
 sg13g2_mux4_1 _2240_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit14.Q ),
    .A0(net953),
    .A1(_1084_),
    .A2(_0148_),
    .A3(_0538_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit15.Q ),
    .X(_0869_));
 sg13g2_mux2_1 _2241_ (.A0(_0868_),
    .A1(_0869_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit16.Q ),
    .X(\Inst_LUT4AB_switch_matrix.WW4BEG0 ));
 sg13g2_mux4_1 _2242_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit3.Q ),
    .A0(net1009),
    .A1(net1216),
    .A2(net88),
    .A3(D),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit4.Q ),
    .X(_0870_));
 sg13g2_nor2_1 _2243_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit5.Q ),
    .B(_0870_),
    .Y(_0871_));
 sg13g2_nand2_2 _2244_ (.Y(_0872_),
    .A(_0276_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit3.Q ));
 sg13g2_o21ai_1 _2245_ (.B1(_0872_),
    .Y(_0873_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit3.Q ),
    .A2(net967));
 sg13g2_nand2_1 _2246_ (.Y(_0874_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit3.Q ),
    .B(_0023_));
 sg13g2_o21ai_1 _2247_ (.B1(_0874_),
    .Y(_0875_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit3.Q ),
    .A2(_0556_));
 sg13g2_o21ai_1 _2248_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit5.Q ),
    .Y(_0876_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit4.Q ),
    .A2(_0873_));
 sg13g2_a21oi_2 _2249_ (.B1(_0876_),
    .Y(_0877_),
    .A2(_0875_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit4.Q ));
 sg13g2_nor2_2 _2250_ (.A(_0871_),
    .B(_0877_),
    .Y(\Inst_LUT4AB_switch_matrix.SS4BEG3 ));
 sg13g2_o21ai_1 _2251_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit1.Q ),
    .Y(_0878_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit0.Q ),
    .A2(net980));
 sg13g2_a21oi_1 _2252_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit0.Q ),
    .A2(_0430_),
    .Y(_0879_),
    .B1(_0878_));
 sg13g2_nor2b_1 _2253_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit0.Q ),
    .B_N(net940),
    .Y(_0880_));
 sg13g2_a21oi_1 _2254_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit0.Q ),
    .A2(_0308_),
    .Y(_0881_),
    .B1(_0880_));
 sg13g2_o21ai_1 _2255_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit2.Q ),
    .Y(_0882_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit1.Q ),
    .A2(_0881_));
 sg13g2_nor2_1 _2256_ (.A(_0879_),
    .B(_0882_),
    .Y(_0883_));
 sg13g2_mux4_1 _2257_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit1.Q ),
    .A0(net31),
    .A1(net87),
    .A2(net1217),
    .A3(net970),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit0.Q ),
    .X(_0884_));
 sg13g2_nor2_1 _2258_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit2.Q ),
    .B(_0884_),
    .Y(_0885_));
 sg13g2_nor2_1 _2259_ (.A(_0883_),
    .B(_0885_),
    .Y(\Inst_LUT4AB_switch_matrix.SS4BEG2 ));
 sg13g2_mux4_1 _2260_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit29.Q ),
    .A0(net1007),
    .A1(net1214),
    .A2(net1003),
    .A3(net975),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit30.Q ),
    .X(_0886_));
 sg13g2_nor2_1 _2261_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit31.Q ),
    .B(_0886_),
    .Y(_0887_));
 sg13g2_mux2_1 _2262_ (.A0(_0197_),
    .A1(_0316_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit29.Q ),
    .X(_0888_));
 sg13g2_nor2_1 _2263_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit29.Q ),
    .B(net932),
    .Y(_0889_));
 sg13g2_a21oi_1 _2264_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit29.Q ),
    .A2(_1157_),
    .Y(_0890_),
    .B1(_0889_));
 sg13g2_o21ai_1 _2265_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit31.Q ),
    .Y(_0891_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit30.Q ),
    .A2(_0890_));
 sg13g2_a21oi_1 _2266_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit30.Q ),
    .A2(_0888_),
    .Y(_0892_),
    .B1(_0891_));
 sg13g2_nor2_1 _2267_ (.A(_0887_),
    .B(_0892_),
    .Y(\Inst_LUT4AB_switch_matrix.SS4BEG1 ));
 sg13g2_o21ai_1 _2268_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit27.Q ),
    .Y(_0893_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit26.Q ),
    .A2(_0148_));
 sg13g2_a21oi_1 _2269_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit26.Q ),
    .A2(_0626_),
    .Y(_0894_),
    .B1(_0893_));
 sg13g2_nor2b_1 _2270_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit26.Q ),
    .B_N(net952),
    .Y(_0895_));
 sg13g2_a21oi_1 _2271_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit26.Q ),
    .A2(_1084_),
    .Y(_0896_),
    .B1(_0895_));
 sg13g2_o21ai_1 _2272_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit28.Q ),
    .Y(_0897_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit27.Q ),
    .A2(_0896_));
 sg13g2_nor2_1 _2273_ (.A(_0894_),
    .B(_0897_),
    .Y(_0898_));
 sg13g2_mux4_1 _2274_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit27.Q ),
    .A0(net1008),
    .A1(net1005),
    .A2(net1215),
    .A3(net957),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit26.Q ),
    .X(_0899_));
 sg13g2_nor2_2 _2275_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit28.Q ),
    .B(_0899_),
    .Y(_0900_));
 sg13g2_nor2_2 _2276_ (.A(_0898_),
    .B(_0900_),
    .Y(\Inst_LUT4AB_switch_matrix.SS4BEG0 ));
 sg13g2_a21oi_1 _2277_ (.A1(net1004),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit6.Q ),
    .Y(_0901_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit7.Q ));
 sg13g2_o21ai_1 _2278_ (.B1(_0901_),
    .Y(_0902_),
    .A1(_1013_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit6.Q ));
 sg13g2_nor2b_1 _2279_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit6.Q ),
    .B_N(net978),
    .Y(_0903_));
 sg13g2_a21oi_1 _2280_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit6.Q ),
    .A2(net971),
    .Y(_0904_),
    .B1(_0903_));
 sg13g2_a21oi_1 _2281_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit7.Q ),
    .A2(_0904_),
    .Y(_0905_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit8.Q ));
 sg13g2_mux4_1 _2282_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit6.Q ),
    .A0(net941),
    .A1(net946),
    .A2(net965),
    .A3(net958),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit7.Q ),
    .X(_0906_));
 sg13g2_a221oi_1 _2283_ (.B2(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit8.Q ),
    .C1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit9.Q ),
    .B1(_0906_),
    .A1(_0902_),
    .Y(_0907_),
    .A2(_0905_));
 sg13g2_mux4_1 _2284_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit6.Q ),
    .A0(_1158_),
    .A1(_0196_),
    .A2(_0276_),
    .A3(_0556_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit7.Q ),
    .X(_0908_));
 sg13g2_mux4_1 _2285_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit6.Q ),
    .A0(net953),
    .A1(net936),
    .A2(net931),
    .A3(net929),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit7.Q ),
    .X(_0909_));
 sg13g2_o21ai_1 _2286_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit9.Q ),
    .Y(_0910_),
    .A1(_1049_),
    .A2(_0908_));
 sg13g2_a21oi_2 _2287_ (.B1(_0910_),
    .Y(_0911_),
    .A2(_0909_),
    .A1(_1049_));
 sg13g2_nor2_2 _2288_ (.A(_0907_),
    .B(_0911_),
    .Y(\Inst_LUT4AB_switch_matrix.E6BEG1 ));
 sg13g2_mux4_1 _2289_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit2.Q ),
    .A0(net1214),
    .A1(net1003),
    .A2(net978),
    .A3(net973),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit3.Q ),
    .X(_0912_));
 sg13g2_mux4_1 _2290_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit2.Q ),
    .A0(net943),
    .A1(net948),
    .A2(net965),
    .A3(net960),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit3.Q ),
    .X(_0913_));
 sg13g2_mux4_1 _2291_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit2.Q ),
    .A0(net953),
    .A1(net936),
    .A2(net930),
    .A3(net928),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit3.Q ),
    .X(_0914_));
 sg13g2_mux4_1 _2292_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit2.Q ),
    .A0(_1084_),
    .A1(_0148_),
    .A2(_0308_),
    .A3(net981),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit3.Q ),
    .X(_0915_));
 sg13g2_mux4_1 _2293_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit4.Q ),
    .A0(_0912_),
    .A1(_0913_),
    .A2(_0914_),
    .A3(_0915_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit5.Q ),
    .X(\Inst_LUT4AB_switch_matrix.E6BEG0 ));
 sg13g2_mux4_1 _2294_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit31.Q ),
    .A0(net1009),
    .A1(net1216),
    .A2(net60),
    .A3(net948),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit0.Q ),
    .X(_0916_));
 sg13g2_nor2_1 _2295_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit1.Q ),
    .B(_0916_),
    .Y(_0917_));
 sg13g2_nand2_1 _2296_ (.Y(_0918_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit31.Q ),
    .B(_1119_));
 sg13g2_o21ai_1 _2297_ (.B1(_0918_),
    .Y(_0919_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit31.Q ),
    .A2(_0556_));
 sg13g2_nand2_2 _2298_ (.Y(_0920_),
    .A(_0276_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit31.Q ));
 sg13g2_o21ai_1 _2299_ (.B1(_0920_),
    .Y(_0921_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit31.Q ),
    .A2(net967));
 sg13g2_o21ai_1 _2300_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit1.Q ),
    .Y(_0922_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit0.Q ),
    .A2(_0921_));
 sg13g2_a21oi_2 _2301_ (.B1(_0922_),
    .Y(_0923_),
    .A2(_0919_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit0.Q ));
 sg13g2_nor2_2 _2302_ (.A(_0917_),
    .B(_0923_),
    .Y(\Inst_LUT4AB_switch_matrix.EE4BEG3 ));
 sg13g2_mux4_1 _2303_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit28.Q ),
    .A0(net943),
    .A1(_0308_),
    .A2(net980),
    .A3(_0366_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit29.Q ),
    .X(_0924_));
 sg13g2_inv_1 _2304_ (.Y(_0925_),
    .A(_0924_));
 sg13g2_a21oi_1 _2305_ (.A1(_1016_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit28.Q ),
    .Y(_0926_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit29.Q ));
 sg13g2_o21ai_1 _2306_ (.B1(_0926_),
    .Y(_0927_),
    .A1(net1010),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit28.Q ));
 sg13g2_mux2_1 _2307_ (.A0(net59),
    .A1(net973),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit28.Q ),
    .X(_0928_));
 sg13g2_a21oi_1 _2308_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit29.Q ),
    .A2(_0928_),
    .Y(_0929_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit30.Q ));
 sg13g2_a22oi_1 _2309_ (.Y(\Inst_LUT4AB_switch_matrix.EE4BEG2 ),
    .B1(_0927_),
    .B2(_0929_),
    .A2(_0925_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit30.Q ));
 sg13g2_mux4_1 _2310_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit25.Q ),
    .A0(net937),
    .A1(_1157_),
    .A2(_0197_),
    .A3(_0239_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit26.Q ),
    .X(_0930_));
 sg13g2_mux4_1 _2311_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit25.Q ),
    .A0(net1007),
    .A1(net1214),
    .A2(net62),
    .A3(net978),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit26.Q ),
    .X(_0931_));
 sg13g2_mux2_1 _2312_ (.A0(_0931_),
    .A1(_0930_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit27.Q ),
    .X(\Inst_LUT4AB_switch_matrix.EE4BEG1 ));
 sg13g2_o21ai_1 _2313_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit23.Q ),
    .Y(_0932_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit22.Q ),
    .A2(_0148_));
 sg13g2_a21oi_1 _2314_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit22.Q ),
    .A2(_0529_),
    .Y(_0933_),
    .B1(_0932_));
 sg13g2_nor2b_1 _2315_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit22.Q ),
    .B_N(net954),
    .Y(_0934_));
 sg13g2_a21oi_1 _2316_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit22.Q ),
    .A2(_1084_),
    .Y(_0935_),
    .B1(_0934_));
 sg13g2_o21ai_1 _2317_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit24.Q ),
    .Y(_0936_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit23.Q ),
    .A2(_0935_));
 sg13g2_nor2_1 _2318_ (.A(_0933_),
    .B(_0936_),
    .Y(_0937_));
 sg13g2_mux4_1 _2319_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit23.Q ),
    .A0(net1008),
    .A1(net61),
    .A2(net1215),
    .A3(net960),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit22.Q ),
    .X(_0938_));
 sg13g2_nor2_1 _2320_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit24.Q ),
    .B(_0938_),
    .Y(_0939_));
 sg13g2_nor2_1 _2321_ (.A(_0937_),
    .B(_0939_),
    .Y(\Inst_LUT4AB_switch_matrix.EE4BEG0 ));
 sg13g2_mux2_1 _2322_ (.A0(net1009),
    .A1(net1216),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit11.Q ),
    .X(_0940_));
 sg13g2_mux2_1 _2323_ (.A0(net1006),
    .A1(net948),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit11.Q ),
    .X(_0941_));
 sg13g2_nor2_1 _2324_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit11.Q ),
    .B(net967),
    .Y(_0942_));
 sg13g2_a21oi_2 _2325_ (.B1(_0942_),
    .Y(_0943_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit11.Q ),
    .A1(_0276_));
 sg13g2_nand2_1 _2326_ (.Y(_0944_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit11.Q ),
    .B(_1066_));
 sg13g2_o21ai_1 _2327_ (.B1(_0944_),
    .Y(_0945_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit11.Q ),
    .A2(_0556_));
 sg13g2_mux4_1 _2328_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit12.Q ),
    .A0(_0940_),
    .A1(_0941_),
    .A2(_0943_),
    .A3(_0945_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit13.Q ),
    .X(\Inst_LUT4AB_switch_matrix.NN4BEG3 ));
 sg13g2_or2_1 _2329_ (.X(_0946_),
    .B(net980),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit8.Q ));
 sg13g2_nand2b_1 _2330_ (.Y(_0947_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit8.Q ),
    .A_N(_0130_));
 sg13g2_nand3_1 _2331_ (.B(_0946_),
    .C(_0947_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit9.Q ),
    .Y(_0948_));
 sg13g2_nor2b_1 _2332_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit8.Q ),
    .B_N(net943),
    .Y(_0949_));
 sg13g2_a21oi_1 _2333_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit8.Q ),
    .A2(_0308_),
    .Y(_0950_),
    .B1(_0949_));
 sg13g2_o21ai_1 _2334_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit10.Q ),
    .Y(_0951_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit9.Q ),
    .A2(_0950_));
 sg13g2_inv_1 _2335_ (.Y(_0952_),
    .A(_0951_));
 sg13g2_mux4_1 _2336_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit9.Q ),
    .A0(net1010),
    .A1(net87),
    .A2(net1217),
    .A3(net973),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit8.Q ),
    .X(_0953_));
 sg13g2_nor2_1 _2337_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit10.Q ),
    .B(_0953_),
    .Y(_0954_));
 sg13g2_a21oi_2 _2338_ (.B1(_0954_),
    .Y(\Inst_LUT4AB_switch_matrix.NN4BEG2 ),
    .A2(_0948_),
    .A1(_0952_));
 sg13g2_mux4_1 _2339_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit5.Q ),
    .A0(net932),
    .A1(_1158_),
    .A2(_0196_),
    .A3(_0290_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit6.Q ),
    .X(_0955_));
 sg13g2_mux4_1 _2340_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit5.Q ),
    .A0(net1007),
    .A1(net1214),
    .A2(net1003),
    .A3(net978),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit6.Q ),
    .X(_0956_));
 sg13g2_nand2_1 _2341_ (.Y(_0957_),
    .A(_1050_),
    .B(_0956_));
 sg13g2_o21ai_1 _2342_ (.B1(_0957_),
    .Y(\Inst_LUT4AB_switch_matrix.NN4BEG1 ),
    .A1(_1050_),
    .A2(_0955_));
 sg13g2_o21ai_1 _2343_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit3.Q ),
    .Y(_0958_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit2.Q ),
    .A2(_0148_));
 sg13g2_a21oi_1 _2344_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit2.Q ),
    .A2(_0589_),
    .Y(_0959_),
    .B1(_0958_));
 sg13g2_nor2b_1 _2345_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit2.Q ),
    .B_N(net954),
    .Y(_0960_));
 sg13g2_a21oi_1 _2346_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit2.Q ),
    .A2(_1084_),
    .Y(_0961_),
    .B1(_0960_));
 sg13g2_o21ai_1 _2347_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit4.Q ),
    .Y(_0962_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit3.Q ),
    .A2(_0961_));
 sg13g2_nor2_1 _2348_ (.A(_0959_),
    .B(_0962_),
    .Y(_0963_));
 sg13g2_mux4_1 _2349_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit3.Q ),
    .A0(net1008),
    .A1(net1005),
    .A2(net1215),
    .A3(net960),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit2.Q ),
    .X(_0964_));
 sg13g2_nor2_1 _2350_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit4.Q ),
    .B(_0964_),
    .Y(_0965_));
 sg13g2_nor2_1 _2351_ (.A(_0963_),
    .B(_0965_),
    .Y(\Inst_LUT4AB_switch_matrix.NN4BEG0 ));
 sg13g2_mux4_1 _2352_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit12.Q ),
    .A0(A),
    .A1(_1159_),
    .A2(\Inst_LUT4AB_switch_matrix.JS2BEG2 ),
    .A3(_1118_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit13.Q ),
    .X(\Inst_LUT4AB_switch_matrix.W1BEG3 ));
 sg13g2_mux4_1 _2353_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit11.Q ),
    .A0(net934),
    .A1(\Inst_LUT4AB_switch_matrix.JS2BEG1 ),
    .A2(net980),
    .A3(_0623_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit10.Q ),
    .X(\Inst_LUT4AB_switch_matrix.W1BEG2 ));
 sg13g2_mux4_1 _2354_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit8.Q ),
    .A0(net950),
    .A1(_0237_),
    .A2(\Inst_LUT4AB_switch_matrix.JS2BEG0 ),
    .A3(net376),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit9.Q ),
    .X(\Inst_LUT4AB_switch_matrix.W1BEG1 ));
 sg13g2_mux4_1 _2355_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit7.Q ),
    .A0(net955),
    .A1(\Inst_LUT4AB_switch_matrix.JS2BEG3 ),
    .A2(_0453_),
    .A3(_0129_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit6.Q ),
    .X(\Inst_LUT4AB_switch_matrix.W1BEG0 ));
 sg13g2_mux4_1 _2356_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit24.Q ),
    .A0(net64),
    .A1(net79),
    .A2(net106),
    .A3(net945),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit25.Q ),
    .X(\Inst_LUT4AB_switch_matrix.S4BEG3 ));
 sg13g2_mux4_1 _2357_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit23.Q ),
    .A0(net63),
    .A1(net107),
    .A2(net82),
    .A3(net940),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit22.Q ),
    .X(\Inst_LUT4AB_switch_matrix.S4BEG2 ));
 sg13g2_mux4_1 _2358_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit21.Q ),
    .A0(net1212),
    .A1(net81),
    .A2(net66),
    .A3(net970),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit20.Q ),
    .X(\Inst_LUT4AB_switch_matrix.S4BEG1 ));
 sg13g2_mux4_1 _2359_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit19.Q ),
    .A0(net1210),
    .A1(net80),
    .A2(net65),
    .A3(net975),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit18.Q ),
    .X(\Inst_LUT4AB_switch_matrix.S4BEG0 ));
 sg13g2_mux4_1 _2360_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit16.Q ),
    .A0(net934),
    .A1(_1159_),
    .A2(\Inst_LUT4AB_switch_matrix.E2BEG2 ),
    .A3(_1118_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit17.Q ),
    .X(\Inst_LUT4AB_switch_matrix.S1BEG3 ));
 sg13g2_mux4_1 _2361_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit15.Q ),
    .A0(net952),
    .A1(net382),
    .A2(net980),
    .A3(_0623_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit14.Q ),
    .X(\Inst_LUT4AB_switch_matrix.S1BEG2 ));
 sg13g2_mux4_1 _2362_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit12.Q ),
    .A0(net957),
    .A1(_0237_),
    .A2(\Inst_LUT4AB_switch_matrix.E2BEG0 ),
    .A3(net376),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit13.Q ),
    .X(\Inst_LUT4AB_switch_matrix.S1BEG1 ));
 sg13g2_mux4_1 _2363_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit11.Q ),
    .A0(net962),
    .A1(\Inst_LUT4AB_switch_matrix.E2BEG3 ),
    .A2(_0453_),
    .A3(_0129_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit10.Q ),
    .X(\Inst_LUT4AB_switch_matrix.S1BEG0 ));
 sg13g2_mux4_1 _2364_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit20.Q ),
    .A0(net952),
    .A1(_1159_),
    .A2(\Inst_LUT4AB_switch_matrix.JN2BEG2 ),
    .A3(_1118_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit21.Q ),
    .X(\Inst_LUT4AB_switch_matrix.E1BEG3 ));
 sg13g2_mux4_1 _2365_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit19.Q ),
    .A0(net957),
    .A1(\Inst_LUT4AB_switch_matrix.JN2BEG1 ),
    .A2(net980),
    .A3(_0623_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit18.Q ),
    .X(\Inst_LUT4AB_switch_matrix.E1BEG2 ));
 sg13g2_mux4_1 _2366_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit16.Q ),
    .A0(net964),
    .A1(_0237_),
    .A2(\Inst_LUT4AB_switch_matrix.JN2BEG0 ),
    .A3(_0248_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit17.Q ),
    .X(\Inst_LUT4AB_switch_matrix.E1BEG1 ));
 sg13g2_mux4_1 _2367_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit15.Q ),
    .A0(net945),
    .A1(\Inst_LUT4AB_switch_matrix.JN2BEG3 ),
    .A2(_0453_),
    .A3(_0129_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit14.Q ),
    .X(\Inst_LUT4AB_switch_matrix.E1BEG0 ));
 sg13g2_mux4_1 _2368_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit1.Q ),
    .A0(net36),
    .A1(net106),
    .A2(net51),
    .A3(net935),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit0.Q ),
    .X(\Inst_LUT4AB_switch_matrix.N4BEG3 ));
 sg13g2_mux4_1 _2369_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit30.Q ),
    .A0(net35),
    .A1(net54),
    .A2(net107),
    .A3(net951),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit31.Q ),
    .X(\Inst_LUT4AB_switch_matrix.N4BEG2 ));
 sg13g2_mux4_1 _2370_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit28.Q ),
    .A0(net38),
    .A1(net53),
    .A2(net1213),
    .A3(net958),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit29.Q ),
    .X(\Inst_LUT4AB_switch_matrix.N4BEG1 ));
 sg13g2_mux4_1 _2371_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit26.Q ),
    .A0(net37),
    .A1(net52),
    .A2(net1211),
    .A3(net963),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit27.Q ),
    .X(\Inst_LUT4AB_switch_matrix.N4BEG0 ));
 sg13g2_mux4_1 _2372_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit24.Q ),
    .A0(net957),
    .A1(_1159_),
    .A2(net384),
    .A3(_1118_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit25.Q ),
    .X(\Inst_LUT4AB_switch_matrix.N1BEG3 ));
 sg13g2_mux4_1 _2373_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit23.Q ),
    .A0(net963),
    .A1(\Inst_LUT4AB_switch_matrix.JW2BEG1 ),
    .A2(net980),
    .A3(_0623_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit22.Q ),
    .X(\Inst_LUT4AB_switch_matrix.N1BEG2 ));
 sg13g2_mux4_1 _2374_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit20.Q ),
    .A0(net947),
    .A1(_0237_),
    .A2(\Inst_LUT4AB_switch_matrix.JW2BEG0 ),
    .A3(net375),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit21.Q ),
    .X(\Inst_LUT4AB_switch_matrix.N1BEG1 ));
 sg13g2_mux4_1 _2375_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit19.Q ),
    .A0(net939),
    .A1(\Inst_LUT4AB_switch_matrix.JW2BEG3 ),
    .A2(_0453_),
    .A3(_0129_),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit18.Q ),
    .X(\Inst_LUT4AB_switch_matrix.N1BEG0 ));
 sg13g2_o21ai_1 _2376_ (.B1(_0651_),
    .Y(net112),
    .A1(_0652_),
    .A2(_0639_));
 sg13g2_nand2b_1 _2377_ (.Y(_0966_),
    .B(_0617_),
    .A_N(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit29.Q ));
 sg13g2_a21oi_1 _2378_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit29.Q ),
    .A2(_0048_),
    .Y(_0967_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit30.Q ));
 sg13g2_nor2_1 _2379_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit29.Q ),
    .B(_0453_),
    .Y(_0968_));
 sg13g2_a21oi_1 _2380_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit29.Q ),
    .A2(_0334_),
    .Y(_0969_),
    .B1(_0968_));
 sg13g2_mux4_1 _2381_ (.S0(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit30.Q ),
    .A0(\Inst_LUT4AB_switch_matrix.JN2BEG2 ),
    .A1(\Inst_LUT4AB_switch_matrix.JS2BEG2 ),
    .A2(\Inst_LUT4AB_switch_matrix.E2BEG2 ),
    .A3(net384),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit29.Q ),
    .X(_0970_));
 sg13g2_nand2_1 _2382_ (.Y(_0971_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit31.Q ),
    .B(_0970_));
 sg13g2_a22oi_1 _2383_ (.Y(_0972_),
    .B1(_0969_),
    .B2(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit30.Q ),
    .A2(_0967_),
    .A1(_0966_));
 sg13g2_o21ai_1 _2384_ (.B1(_0971_),
    .Y(_0973_),
    .A1(_0972_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit31.Q ));
 sg13g2_nand2b_1 _2385_ (.Y(_0974_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit8.Q ),
    .A_N(_0973_));
 sg13g2_nand3b_1 _2386_ (.B(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit8.Q ),
    .C(net397),
    .Y(_0975_),
    .A_N(_0973_));
 sg13g2_nand2b_1 _2387_ (.Y(_0976_),
    .B(net385),
    .A_N(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q ));
 sg13g2_a21oi_1 _2388_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q ),
    .A2(_1104_),
    .Y(_0977_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit27.Q ));
 sg13g2_mux2_1 _2389_ (.A0(_0390_),
    .A1(_0237_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q ),
    .X(_0978_));
 sg13g2_a221oi_1 _2390_ (.B2(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit27.Q ),
    .C1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit28.Q ),
    .B1(_0978_),
    .A1(_0976_),
    .Y(_0979_),
    .A2(_0977_));
 sg13g2_o21ai_1 _2391_ (.B1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit27.Q ),
    .Y(_0980_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q ),
    .A2(\Inst_LUT4AB_switch_matrix.JS2BEG1 ));
 sg13g2_a21oi_1 _2392_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q ),
    .A2(_0021_),
    .Y(_0981_),
    .B1(_0980_));
 sg13g2_a21oi_1 _2393_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q ),
    .A2(_1064_),
    .Y(_0982_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit27.Q ));
 sg13g2_o21ai_1 _2394_ (.B1(_0982_),
    .Y(_0983_),
    .A1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q ),
    .A2(\Inst_LUT4AB_switch_matrix.JN2BEG1 ));
 sg13g2_nor2b_1 _2395_ (.A(_0981_),
    .B_N(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit28.Q ),
    .Y(_0984_));
 sg13g2_a21oi_2 _2396_ (.B1(_0979_),
    .Y(_0985_),
    .A2(_0984_),
    .A1(_0983_));
 sg13g2_nand2_1 _2397_ (.Y(_0986_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit17.Q ),
    .B(_0985_));
 sg13g2_a221oi_1 _2398_ (.B2(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit17.Q ),
    .C1(_0659_),
    .B1(_0985_),
    .A1(_0665_),
    .Y(_0987_),
    .A2(_0661_));
 sg13g2_o21ai_1 _2399_ (.B1(_0974_),
    .Y(_0988_),
    .A1(\Inst_LH_LUT4c_frame_config_dffesr.c_reset_value ),
    .A2(_0986_));
 sg13g2_o21ai_1 _2400_ (.B1(_0975_),
    .Y(_0000_),
    .A1(_0988_),
    .A2(_0987_));
 sg13g2_nand2_1 _2401_ (.Y(_0989_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit11.Q ),
    .B(net925));
 sg13g2_nand2b_1 _2402_ (.Y(_0990_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit2.Q ),
    .A_N(net927));
 sg13g2_mux2_1 _2403_ (.A0(\Inst_LA_LUT4c_frame_config_dffesr.c_reset_value ),
    .A1(_0069_),
    .S(_0989_),
    .X(_0991_));
 sg13g2_mux2_1 _2404_ (.A0(net394),
    .A1(_0991_),
    .S(_0990_),
    .X(_0001_));
 sg13g2_nand2b_1 _2405_ (.Y(_0992_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit12.Q ),
    .A_N(net927));
 sg13g2_nand2_1 _2406_ (.Y(_0993_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit21.Q ),
    .B(net925));
 sg13g2_mux2_1 _2407_ (.A0(\Inst_LB_LUT4c_frame_config_dffesr.c_reset_value ),
    .A1(_0109_),
    .S(_0993_),
    .X(_0994_));
 sg13g2_mux2_1 _2408_ (.A0(net395),
    .A1(_0994_),
    .S(_0992_),
    .X(_0002_));
 sg13g2_nand2b_1 _2409_ (.Y(_0995_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit22.Q ),
    .A_N(net927));
 sg13g2_nand2_1 _2410_ (.Y(_0996_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit31.Q ),
    .B(net925));
 sg13g2_mux2_1 _2411_ (.A0(\Inst_LC_LUT4c_frame_config_dffesr.c_reset_value ),
    .A1(_0467_),
    .S(_0996_),
    .X(_0997_));
 sg13g2_mux2_1 _2412_ (.A0(net392),
    .A1(_0997_),
    .S(_0995_),
    .X(_0003_));
 sg13g2_nand2b_1 _2413_ (.Y(_0998_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit0.Q ),
    .A_N(net927));
 sg13g2_nand2_1 _2414_ (.Y(_0999_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit9.Q ),
    .B(net925));
 sg13g2_mux2_1 _2415_ (.A0(\Inst_LD_LUT4c_frame_config_dffesr.c_reset_value ),
    .A1(_0688_),
    .S(_0999_),
    .X(_1000_));
 sg13g2_mux2_1 _2416_ (.A0(net391),
    .A1(_1000_),
    .S(_0998_),
    .X(_0004_));
 sg13g2_nand2b_1 _2417_ (.Y(_1001_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit10.Q ),
    .A_N(net927));
 sg13g2_nand2_1 _2418_ (.Y(_1002_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit19.Q ),
    .B(net925));
 sg13g2_mux2_1 _2419_ (.A0(\Inst_LE_LUT4c_frame_config_dffesr.c_reset_value ),
    .A1(net389),
    .S(_1002_),
    .X(_1003_));
 sg13g2_mux2_1 _2420_ (.A0(net396),
    .A1(_1003_),
    .S(_1001_),
    .X(_0005_));
 sg13g2_nand2b_1 _2421_ (.Y(_1004_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit20.Q ),
    .A_N(net927));
 sg13g2_nand2_1 _2422_ (.Y(_1005_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit29.Q ),
    .B(net925));
 sg13g2_mux2_1 _2423_ (.A0(\Inst_LF_LUT4c_frame_config_dffesr.c_reset_value ),
    .A1(_0496_),
    .S(_1005_),
    .X(_1006_));
 sg13g2_mux2_1 _2424_ (.A0(net393),
    .A1(_1006_),
    .S(_1004_),
    .X(_0006_));
 sg13g2_nand2b_1 _2425_ (.Y(_1007_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit30.Q ),
    .A_N(net927));
 sg13g2_nand3b_1 _2426_ (.B(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit30.Q ),
    .C(net390),
    .Y(_1008_),
    .A_N(net927));
 sg13g2_nand2_1 _2427_ (.Y(_1009_),
    .A(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit7.Q ),
    .B(net925));
 sg13g2_a221oi_1 _2428_ (.B2(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit7.Q ),
    .C1(_0630_),
    .B1(net925),
    .A1(_0632_),
    .Y(_1010_),
    .A2(_0635_));
 sg13g2_o21ai_1 _2429_ (.B1(_1007_),
    .Y(_1011_),
    .A1(\Inst_LG_LUT4c_frame_config_dffesr.c_reset_value ),
    .A2(_1009_));
 sg13g2_o21ai_1 _2430_ (.B1(_1008_),
    .Y(_0007_),
    .A1(_1010_),
    .A2(_1011_));
 sg13g2_dlhq_1 _2431_ (.D(net1160),
    .GATE(net1059),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ));
 sg13g2_dlhq_1 _2432_ (.D(net1157),
    .GATE(net1059),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ));
 sg13g2_dlhq_1 _2433_ (.D(net1153),
    .GATE(net1059),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ));
 sg13g2_dlhq_1 _2434_ (.D(net1150),
    .GATE(net1059),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ));
 sg13g2_dlhq_1 _2435_ (.D(net1147),
    .GATE(net1059),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ));
 sg13g2_dlhq_1 _2436_ (.D(net1144),
    .GATE(net28),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ));
 sg13g2_dlhq_1 _2437_ (.D(net1139),
    .GATE(net1059),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ));
 sg13g2_dlhq_1 _2438_ (.D(net1136),
    .GATE(net1059),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ));
 sg13g2_dlhq_1 _2439_ (.D(net1209),
    .GATE(net1060),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ));
 sg13g2_dlhq_1 _2440_ (.D(net1175),
    .GATE(net1060),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ));
 sg13g2_dlhq_1 _2441_ (.D(net1143),
    .GATE(net1061),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ));
 sg13g2_dlhq_1 _2442_ (.D(net1134),
    .GATE(net1061),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ));
 sg13g2_dlhq_1 _2443_ (.D(net1131),
    .GATE(net1060),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ));
 sg13g2_dlhq_1 _2444_ (.D(net1128),
    .GATE(net1060),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ));
 sg13g2_dlhq_1 _2445_ (.D(net1124),
    .GATE(net1060),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ));
 sg13g2_dlhq_1 _2446_ (.D(net1121),
    .GATE(net1060),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ));
 sg13g2_dlhq_1 _2447_ (.D(net1117),
    .GATE(net1062),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.c_out_mux ));
 sg13g2_dlhq_1 _2448_ (.D(net1114),
    .GATE(net1062),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.c_I0mux ));
 sg13g2_dlhq_1 _2449_ (.D(net1204),
    .GATE(net1062),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.c_reset_value ));
 sg13g2_dlhq_1 _2450_ (.D(net1202),
    .GATE(net1061),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ));
 sg13g2_dlhq_1 _2451_ (.D(net1199),
    .GATE(net1061),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ));
 sg13g2_dlhq_1 _2452_ (.D(net1196),
    .GATE(net1061),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ));
 sg13g2_dlhq_1 _2453_ (.D(net1193),
    .GATE(net1063),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ));
 sg13g2_dlhq_1 _2454_ (.D(net1190),
    .GATE(net1061),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ));
 sg13g2_dlhq_1 _2455_ (.D(net1187),
    .GATE(net1063),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ));
 sg13g2_dlhq_1 _2456_ (.D(net1184),
    .GATE(net1060),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ));
 sg13g2_dlhq_1 _2457_ (.D(net1181),
    .GATE(net1060),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ));
 sg13g2_dlhq_1 _2458_ (.D(net1178),
    .GATE(net1063),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ));
 sg13g2_dlhq_1 _2459_ (.D(net1172),
    .GATE(net1063),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ));
 sg13g2_dlhq_1 _2460_ (.D(net1169),
    .GATE(net1063),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ));
 sg13g2_dlhq_1 _2461_ (.D(net1166),
    .GATE(net1064),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ));
 sg13g2_dlhq_1 _2462_ (.D(net1163),
    .GATE(net1063),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ));
 sg13g2_dlhq_1 _2463_ (.D(net1160),
    .GATE(net1063),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ));
 sg13g2_dlhq_1 _2464_ (.D(net1157),
    .GATE(net1064),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ));
 sg13g2_dlhq_1 _2465_ (.D(net1153),
    .GATE(net1063),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ));
 sg13g2_dlhq_1 _2466_ (.D(net1150),
    .GATE(net1065),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.c_out_mux ));
 sg13g2_dlhq_1 _2467_ (.D(net1147),
    .GATE(net1065),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.c_I0mux ));
 sg13g2_dlhq_1 _2468_ (.D(net1144),
    .GATE(net1065),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.c_reset_value ));
 sg13g2_dlhq_1 _2469_ (.D(net1139),
    .GATE(net1064),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ));
 sg13g2_dlhq_1 _2470_ (.D(net1136),
    .GATE(net1064),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ));
 sg13g2_dlhq_1 _2471_ (.D(net1209),
    .GATE(net1067),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ));
 sg13g2_dlhq_1 _2472_ (.D(net1175),
    .GATE(net1067),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ));
 sg13g2_dlhq_1 _2473_ (.D(net1143),
    .GATE(net1067),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ));
 sg13g2_dlhq_1 _2474_ (.D(net1134),
    .GATE(net1067),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ));
 sg13g2_dlhq_1 _2475_ (.D(net1131),
    .GATE(net1067),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ));
 sg13g2_dlhq_1 _2476_ (.D(net1128),
    .GATE(net1066),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ));
 sg13g2_dlhq_1 _2477_ (.D(net1124),
    .GATE(net1066),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ));
 sg13g2_dlhq_1 _2478_ (.D(net1121),
    .GATE(net1066),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ));
 sg13g2_dlhq_1 _2479_ (.D(net1117),
    .GATE(net1066),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ));
 sg13g2_dlhq_1 _2480_ (.D(net1114),
    .GATE(net1066),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ));
 sg13g2_dlhq_1 _2481_ (.D(net1204),
    .GATE(net1066),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ));
 sg13g2_dlhq_1 _2482_ (.D(net1202),
    .GATE(net1066),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ));
 sg13g2_dlhq_1 _2483_ (.D(net1199),
    .GATE(net1066),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ));
 sg13g2_dlhq_1 _2484_ (.D(net1196),
    .GATE(net1067),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ));
 sg13g2_dlhq_1 _2485_ (.D(net1193),
    .GATE(net1068),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.c_out_mux ));
 sg13g2_dlhq_1 _2486_ (.D(net1190),
    .GATE(net1068),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.c_I0mux ));
 sg13g2_dlhq_1 _2487_ (.D(net1187),
    .GATE(net1068),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.c_reset_value ));
 sg13g2_dlhq_1 _2488_ (.D(net1184),
    .GATE(net1070),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ));
 sg13g2_dlhq_1 _2489_ (.D(net1181),
    .GATE(net1069),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ));
 sg13g2_dlhq_1 _2490_ (.D(net1178),
    .GATE(net1070),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ));
 sg13g2_dlhq_1 _2491_ (.D(net1172),
    .GATE(net1070),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ));
 sg13g2_dlhq_1 _2492_ (.D(net1169),
    .GATE(net1070),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ));
 sg13g2_dlhq_1 _2493_ (.D(net1166),
    .GATE(net1069),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ));
 sg13g2_dlhq_1 _2494_ (.D(net1163),
    .GATE(net1070),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ));
 sg13g2_dlhq_1 _2495_ (.D(net1161),
    .GATE(net1069),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ));
 sg13g2_dlhq_1 _2496_ (.D(net1158),
    .GATE(net1069),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ));
 sg13g2_dlhq_1 _2497_ (.D(net1154),
    .GATE(net1069),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ));
 sg13g2_dlhq_1 _2498_ (.D(net1150),
    .GATE(net1069),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ));
 sg13g2_dlhq_1 _2499_ (.D(net1148),
    .GATE(net1070),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ));
 sg13g2_dlhq_1 _2500_ (.D(net1144),
    .GATE(net1069),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ));
 sg13g2_dlhq_1 _2501_ (.D(net1140),
    .GATE(net1070),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ));
 sg13g2_dlhq_1 _2502_ (.D(net1136),
    .GATE(net1069),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ));
 sg13g2_dlhq_1 _2503_ (.D(net1208),
    .GATE(net1074),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ));
 sg13g2_dlhq_1 _2504_ (.D(net1176),
    .GATE(net1074),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.c_out_mux ));
 sg13g2_dlhq_1 _2505_ (.D(net1142),
    .GATE(net1074),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.c_I0mux ));
 sg13g2_dlhq_1 _2506_ (.D(net1133),
    .GATE(net1074),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.c_reset_value ));
 sg13g2_dlhq_1 _2507_ (.D(net1129),
    .GATE(net1071),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ));
 sg13g2_dlhq_1 _2508_ (.D(net1127),
    .GATE(net1071),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ));
 sg13g2_dlhq_1 _2509_ (.D(net1125),
    .GATE(net1071),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ));
 sg13g2_dlhq_1 _2510_ (.D(net1122),
    .GATE(net1071),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ));
 sg13g2_dlhq_1 _2511_ (.D(net1118),
    .GATE(net1071),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ));
 sg13g2_dlhq_1 _2512_ (.D(net1115),
    .GATE(net1071),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ));
 sg13g2_dlhq_1 _2513_ (.D(net1205),
    .GATE(net1071),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ));
 sg13g2_dlhq_1 _2514_ (.D(net1203),
    .GATE(net1071),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ));
 sg13g2_dlhq_1 _2515_ (.D(net1199),
    .GATE(net1072),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ));
 sg13g2_dlhq_1 _2516_ (.D(net1197),
    .GATE(net1072),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ));
 sg13g2_dlhq_1 _2517_ (.D(net1194),
    .GATE(net1072),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ));
 sg13g2_dlhq_1 _2518_ (.D(net1191),
    .GATE(net1072),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ));
 sg13g2_dlhq_1 _2519_ (.D(net1188),
    .GATE(net1072),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ));
 sg13g2_dlhq_1 _2520_ (.D(net1185),
    .GATE(net1072),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ));
 sg13g2_dlhq_1 _2521_ (.D(net1182),
    .GATE(net1072),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ));
 sg13g2_dlhq_1 _2522_ (.D(net1179),
    .GATE(net1072),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ));
 sg13g2_dlhq_1 _2523_ (.D(net1172),
    .GATE(net1073),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.c_out_mux ));
 sg13g2_dlhq_1 _2524_ (.D(net1169),
    .GATE(net1073),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.c_I0mux ));
 sg13g2_dlhq_1 _2525_ (.D(net1166),
    .GATE(net1073),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.c_reset_value ));
 sg13g2_dlhq_1 _2526_ (.D(net1163),
    .GATE(net1075),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ));
 sg13g2_dlhq_1 _2527_ (.D(net1160),
    .GATE(net1075),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ));
 sg13g2_dlhq_1 _2528_ (.D(net1158),
    .GATE(net1075),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ));
 sg13g2_dlhq_1 _2529_ (.D(net1154),
    .GATE(net1075),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ));
 sg13g2_dlhq_1 _2530_ (.D(net1151),
    .GATE(net1075),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ));
 sg13g2_dlhq_1 _2531_ (.D(net1148),
    .GATE(net1075),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ));
 sg13g2_dlhq_1 _2532_ (.D(net1145),
    .GATE(net1075),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ));
 sg13g2_dlhq_1 _2533_ (.D(net1140),
    .GATE(net1076),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ));
 sg13g2_dlhq_1 _2534_ (.D(net1137),
    .GATE(net1076),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ));
 sg13g2_dlhq_1 _2535_ (.D(net1209),
    .GATE(net1078),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ));
 sg13g2_dlhq_1 _2536_ (.D(net26),
    .GATE(net1078),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ));
 sg13g2_dlhq_1 _2537_ (.D(net1142),
    .GATE(net1077),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ));
 sg13g2_dlhq_1 _2538_ (.D(net1133),
    .GATE(net1077),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ));
 sg13g2_dlhq_1 _2539_ (.D(net1129),
    .GATE(net1077),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ));
 sg13g2_dlhq_1 _2540_ (.D(net1127),
    .GATE(net1077),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ));
 sg13g2_dlhq_1 _2541_ (.D(net1125),
    .GATE(net1078),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ));
 sg13g2_dlhq_1 _2542_ (.D(net1121),
    .GATE(net1081),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.c_out_mux ));
 sg13g2_dlhq_1 _2543_ (.D(net1118),
    .GATE(net1078),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.c_I0mux ));
 sg13g2_dlhq_1 _2544_ (.D(net1115),
    .GATE(net1080),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.c_reset_value ));
 sg13g2_dlhq_1 _2545_ (.D(net1205),
    .GATE(net1077),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ));
 sg13g2_dlhq_1 _2546_ (.D(net1202),
    .GATE(net1079),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ));
 sg13g2_dlhq_1 _2547_ (.D(net1199),
    .GATE(net1077),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ));
 sg13g2_dlhq_1 _2548_ (.D(net1196),
    .GATE(net1079),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ));
 sg13g2_dlhq_1 _2549_ (.D(net1193),
    .GATE(net1077),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ));
 sg13g2_dlhq_1 _2550_ (.D(net1191),
    .GATE(net1079),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ));
 sg13g2_dlhq_1 _2551_ (.D(net1187),
    .GATE(net1077),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ));
 sg13g2_dlhq_1 _2552_ (.D(net1185),
    .GATE(net1079),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ));
 sg13g2_dlhq_1 _2553_ (.D(net1182),
    .GATE(net1080),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ));
 sg13g2_dlhq_1 _2554_ (.D(net1179),
    .GATE(net1081),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ));
 sg13g2_dlhq_1 _2555_ (.D(net1172),
    .GATE(net1080),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ));
 sg13g2_dlhq_1 _2556_ (.D(net1169),
    .GATE(net1080),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ));
 sg13g2_dlhq_1 _2557_ (.D(net1166),
    .GATE(net1080),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ));
 sg13g2_dlhq_1 _2558_ (.D(net1163),
    .GATE(net1080),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ));
 sg13g2_dlhq_1 _2559_ (.D(net1160),
    .GATE(net1080),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ));
 sg13g2_dlhq_1 _2560_ (.D(net1157),
    .GATE(net1080),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ));
 sg13g2_dlhq_1 _2561_ (.D(net1154),
    .GATE(net1081),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.c_out_mux ));
 sg13g2_dlhq_1 _2562_ (.D(net1151),
    .GATE(net1079),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.c_I0mux ));
 sg13g2_dlhq_1 _2563_ (.D(net1148),
    .GATE(net1081),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.c_reset_value ));
 sg13g2_dlhq_1 _2564_ (.D(net1145),
    .GATE(net1081),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ));
 sg13g2_dlhq_1 _2565_ (.D(net1140),
    .GATE(net1079),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ));
 sg13g2_dlhq_1 _2566_ (.D(net1137),
    .GATE(net1081),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ));
 sg13g2_dlhq_1 _2567_ (.D(net1208),
    .GATE(net1086),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ));
 sg13g2_dlhq_1 _2568_ (.D(net1176),
    .GATE(net1083),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ));
 sg13g2_dlhq_1 _2569_ (.D(net1142),
    .GATE(net1083),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ));
 sg13g2_dlhq_1 _2570_ (.D(net1132),
    .GATE(net1083),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ));
 sg13g2_dlhq_1 _2571_ (.D(net1130),
    .GATE(net1083),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ));
 sg13g2_dlhq_1 _2572_ (.D(net1127),
    .GATE(net1084),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ));
 sg13g2_dlhq_1 _2573_ (.D(net1124),
    .GATE(net1083),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ));
 sg13g2_dlhq_1 _2574_ (.D(net1122),
    .GATE(net1084),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ));
 sg13g2_dlhq_1 _2575_ (.D(net1118),
    .GATE(net1084),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ));
 sg13g2_dlhq_1 _2576_ (.D(net1114),
    .GATE(net1084),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ));
 sg13g2_dlhq_1 _2577_ (.D(net1205),
    .GATE(net1083),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ));
 sg13g2_dlhq_1 _2578_ (.D(net1202),
    .GATE(net1084),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ));
 sg13g2_dlhq_1 _2579_ (.D(net1200),
    .GATE(net1084),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ));
 sg13g2_dlhq_1 _2580_ (.D(net1196),
    .GATE(net1083),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.c_out_mux ));
 sg13g2_dlhq_1 _2581_ (.D(net1194),
    .GATE(net1083),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.c_I0mux ));
 sg13g2_dlhq_1 _2582_ (.D(net1191),
    .GATE(net1084),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.c_reset_value ));
 sg13g2_dlhq_1 _2583_ (.D(net1188),
    .GATE(net1085),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit16.Q ));
 sg13g2_dlhq_1 _2584_ (.D(net1185),
    .GATE(net1085),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit17.Q ));
 sg13g2_dlhq_1 _2585_ (.D(net1180),
    .GATE(net1082),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit18.Q ));
 sg13g2_dlhq_1 _2586_ (.D(net1177),
    .GATE(net1082),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit19.Q ));
 sg13g2_dlhq_1 _2587_ (.D(net1171),
    .GATE(net1085),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit20.Q ));
 sg13g2_dlhq_1 _2588_ (.D(net1168),
    .GATE(net1085),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit21.Q ));
 sg13g2_dlhq_1 _2589_ (.D(net1165),
    .GATE(net1082),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit22.Q ));
 sg13g2_dlhq_1 _2590_ (.D(net1162),
    .GATE(net1082),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit23.Q ));
 sg13g2_dlhq_1 _2591_ (.D(net1159),
    .GATE(net1082),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit24.Q ));
 sg13g2_dlhq_1 _2592_ (.D(net1156),
    .GATE(net1086),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit25.Q ));
 sg13g2_dlhq_1 _2593_ (.D(net1155),
    .GATE(net1082),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit26.Q ));
 sg13g2_dlhq_1 _2594_ (.D(net1152),
    .GATE(net1086),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit27.Q ));
 sg13g2_dlhq_1 _2595_ (.D(net1149),
    .GATE(net1085),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit28.Q ));
 sg13g2_dlhq_1 _2596_ (.D(net1146),
    .GATE(net1085),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit29.Q ));
 sg13g2_dlhq_1 _2597_ (.D(net1138),
    .GATE(net1082),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit30.Q ));
 sg13g2_dlhq_1 _2598_ (.D(net1135),
    .GATE(net1082),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit31.Q ));
 sg13g2_dlhq_1 _2599_ (.D(net1207),
    .GATE(net1087),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit0.Q ));
 sg13g2_dlhq_1 _2600_ (.D(net1174),
    .GATE(net1087),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit1.Q ));
 sg13g2_dlhq_1 _2601_ (.D(net1141),
    .GATE(net1090),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit2.Q ));
 sg13g2_dlhq_1 _2602_ (.D(net1132),
    .GATE(net1091),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit3.Q ));
 sg13g2_dlhq_1 _2603_ (.D(net1129),
    .GATE(net1091),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit4.Q ));
 sg13g2_dlhq_1 _2604_ (.D(net1127),
    .GATE(net1090),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit5.Q ));
 sg13g2_dlhq_1 _2605_ (.D(net1125),
    .GATE(net1090),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit6.Q ));
 sg13g2_dlhq_1 _2606_ (.D(net1120),
    .GATE(net1090),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit7.Q ));
 sg13g2_dlhq_1 _2607_ (.D(net1118),
    .GATE(net1088),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit8.Q ));
 sg13g2_dlhq_1 _2608_ (.D(net1116),
    .GATE(net1088),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit9.Q ));
 sg13g2_dlhq_1 _2609_ (.D(net1205),
    .GATE(net1088),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit10.Q ));
 sg13g2_dlhq_1 _2610_ (.D(net1201),
    .GATE(net1090),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit11.Q ));
 sg13g2_dlhq_1 _2611_ (.D(net1198),
    .GATE(net1090),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit12.Q ));
 sg13g2_dlhq_1 _2612_ (.D(net1195),
    .GATE(net1090),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit13.Q ));
 sg13g2_dlhq_1 _2613_ (.D(net1193),
    .GATE(net1092),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit14.Q ));
 sg13g2_dlhq_1 _2614_ (.D(net1190),
    .GATE(net1087),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit15.Q ));
 sg13g2_dlhq_1 _2615_ (.D(net1187),
    .GATE(net1087),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit16.Q ));
 sg13g2_dlhq_1 _2616_ (.D(net1184),
    .GATE(net1087),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit17.Q ));
 sg13g2_dlhq_1 _2617_ (.D(net1181),
    .GATE(net1087),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit18.Q ));
 sg13g2_dlhq_1 _2618_ (.D(net1178),
    .GATE(net1092),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit19.Q ));
 sg13g2_dlhq_1 _2619_ (.D(net1172),
    .GATE(net1087),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit20.Q ));
 sg13g2_dlhq_1 _2620_ (.D(net1169),
    .GATE(net1087),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit21.Q ));
 sg13g2_dlhq_1 _2621_ (.D(net1166),
    .GATE(net1088),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit22.Q ));
 sg13g2_dlhq_1 _2622_ (.D(net1164),
    .GATE(net1089),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit23.Q ));
 sg13g2_dlhq_1 _2623_ (.D(net1160),
    .GATE(net1089),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit24.Q ));
 sg13g2_dlhq_1 _2624_ (.D(net1158),
    .GATE(net1089),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit25.Q ));
 sg13g2_dlhq_1 _2625_ (.D(net1155),
    .GATE(net1089),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit26.Q ));
 sg13g2_dlhq_1 _2626_ (.D(net1152),
    .GATE(net1089),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit27.Q ));
 sg13g2_dlhq_1 _2627_ (.D(net1148),
    .GATE(net1088),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit28.Q ));
 sg13g2_dlhq_1 _2628_ (.D(net1145),
    .GATE(net1088),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit29.Q ));
 sg13g2_dlhq_1 _2629_ (.D(net1140),
    .GATE(net1088),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit30.Q ));
 sg13g2_dlhq_1 _2630_ (.D(net1137),
    .GATE(net1088),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit31.Q ));
 sg13g2_dlhq_1 _2631_ (.D(net1208),
    .GATE(net1097),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit0.Q ));
 sg13g2_dlhq_1 _2632_ (.D(net1176),
    .GATE(net1097),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit1.Q ));
 sg13g2_dlhq_1 _2633_ (.D(net1141),
    .GATE(net1096),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit2.Q ));
 sg13g2_dlhq_1 _2634_ (.D(net1132),
    .GATE(net1096),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit3.Q ));
 sg13g2_dlhq_1 _2635_ (.D(net1129),
    .GATE(net1096),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit4.Q ));
 sg13g2_dlhq_1 _2636_ (.D(net1127),
    .GATE(net1096),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit5.Q ));
 sg13g2_dlhq_1 _2637_ (.D(net1123),
    .GATE(net1096),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit6.Q ));
 sg13g2_dlhq_1 _2638_ (.D(net1122),
    .GATE(net1096),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit7.Q ));
 sg13g2_dlhq_1 _2639_ (.D(net1119),
    .GATE(net1096),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit8.Q ));
 sg13g2_dlhq_1 _2640_ (.D(net1116),
    .GATE(net1096),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit9.Q ));
 sg13g2_dlhq_1 _2641_ (.D(net1206),
    .GATE(net1093),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit10.Q ));
 sg13g2_dlhq_1 _2642_ (.D(net1201),
    .GATE(net1093),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit11.Q ));
 sg13g2_dlhq_1 _2643_ (.D(net1198),
    .GATE(net1093),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit12.Q ));
 sg13g2_dlhq_1 _2644_ (.D(net1195),
    .GATE(net1093),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit13.Q ));
 sg13g2_dlhq_1 _2645_ (.D(net1192),
    .GATE(net1093),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit14.Q ));
 sg13g2_dlhq_1 _2646_ (.D(net1189),
    .GATE(net1094),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit15.Q ));
 sg13g2_dlhq_1 _2647_ (.D(net1186),
    .GATE(net1093),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit16.Q ));
 sg13g2_dlhq_1 _2648_ (.D(net1183),
    .GATE(net1093),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit17.Q ));
 sg13g2_dlhq_1 _2649_ (.D(net1180),
    .GATE(net1094),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit18.Q ));
 sg13g2_dlhq_1 _2650_ (.D(net1177),
    .GATE(net1094),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit19.Q ));
 sg13g2_dlhq_1 _2651_ (.D(net1171),
    .GATE(net1095),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit20.Q ));
 sg13g2_dlhq_1 _2652_ (.D(net1168),
    .GATE(net1095),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit21.Q ));
 sg13g2_dlhq_1 _2653_ (.D(net1166),
    .GATE(net1095),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit22.Q ));
 sg13g2_dlhq_1 _2654_ (.D(net1162),
    .GATE(net1095),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit23.Q ));
 sg13g2_dlhq_1 _2655_ (.D(net1159),
    .GATE(net1093),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit24.Q ));
 sg13g2_dlhq_1 _2656_ (.D(net1157),
    .GATE(net1094),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit25.Q ));
 sg13g2_dlhq_1 _2657_ (.D(net1153),
    .GATE(net1094),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit26.Q ));
 sg13g2_dlhq_1 _2658_ (.D(net1150),
    .GATE(net1094),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit27.Q ));
 sg13g2_dlhq_1 _2659_ (.D(net1147),
    .GATE(net1094),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit28.Q ));
 sg13g2_dlhq_1 _2660_ (.D(net1146),
    .GATE(net1095),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit29.Q ));
 sg13g2_dlhq_1 _2661_ (.D(net1139),
    .GATE(net1095),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit30.Q ));
 sg13g2_dlhq_1 _2662_ (.D(net1135),
    .GATE(net1095),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit31.Q ));
 sg13g2_dlhq_1 _2663_ (.D(net1209),
    .GATE(net1102),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit0.Q ));
 sg13g2_dlhq_1 _2664_ (.D(net1175),
    .GATE(net1102),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit1.Q ));
 sg13g2_dlhq_1 _2665_ (.D(net1143),
    .GATE(net1102),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit2.Q ));
 sg13g2_dlhq_1 _2666_ (.D(net1133),
    .GATE(net1102),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit3.Q ));
 sg13g2_dlhq_1 _2667_ (.D(net1130),
    .GATE(net1102),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit4.Q ));
 sg13g2_dlhq_1 _2668_ (.D(net1128),
    .GATE(net1102),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit5.Q ));
 sg13g2_dlhq_1 _2669_ (.D(net1123),
    .GATE(net1101),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit6.Q ));
 sg13g2_dlhq_1 _2670_ (.D(net1120),
    .GATE(net1101),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit7.Q ));
 sg13g2_dlhq_1 _2671_ (.D(net1119),
    .GATE(net1101),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit8.Q ));
 sg13g2_dlhq_1 _2672_ (.D(net1116),
    .GATE(net1101),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit9.Q ));
 sg13g2_dlhq_1 _2673_ (.D(net1206),
    .GATE(net1101),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit10.Q ));
 sg13g2_dlhq_1 _2674_ (.D(net1201),
    .GATE(net1101),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit11.Q ));
 sg13g2_dlhq_1 _2675_ (.D(net1198),
    .GATE(net1101),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit12.Q ));
 sg13g2_dlhq_1 _2676_ (.D(net1195),
    .GATE(net27),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit13.Q ));
 sg13g2_dlhq_1 _2677_ (.D(net1194),
    .GATE(net1098),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit14.Q ));
 sg13g2_dlhq_1 _2678_ (.D(net1191),
    .GATE(net1098),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit15.Q ));
 sg13g2_dlhq_1 _2679_ (.D(net1186),
    .GATE(net1098),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit16.Q ));
 sg13g2_dlhq_1 _2680_ (.D(net1183),
    .GATE(net1099),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit17.Q ));
 sg13g2_dlhq_1 _2681_ (.D(net1180),
    .GATE(net1099),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit18.Q ));
 sg13g2_dlhq_1 _2682_ (.D(net1177),
    .GATE(net1098),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit19.Q ));
 sg13g2_dlhq_1 _2683_ (.D(net1171),
    .GATE(net1099),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit20.Q ));
 sg13g2_dlhq_1 _2684_ (.D(net1168),
    .GATE(net1099),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit21.Q ));
 sg13g2_dlhq_1 _2685_ (.D(net1165),
    .GATE(net1099),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit22.Q ));
 sg13g2_dlhq_1 _2686_ (.D(net1162),
    .GATE(net1100),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit23.Q ));
 sg13g2_dlhq_1 _2687_ (.D(net1161),
    .GATE(net1100),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit24.Q ));
 sg13g2_dlhq_1 _2688_ (.D(net1158),
    .GATE(net1100),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit25.Q ));
 sg13g2_dlhq_1 _2689_ (.D(net1155),
    .GATE(net1098),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit26.Q ));
 sg13g2_dlhq_1 _2690_ (.D(net1152),
    .GATE(net1098),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit27.Q ));
 sg13g2_dlhq_1 _2691_ (.D(net1149),
    .GATE(net1098),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit28.Q ));
 sg13g2_dlhq_1 _2692_ (.D(net1146),
    .GATE(net1098),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit29.Q ));
 sg13g2_dlhq_1 _2693_ (.D(net1138),
    .GATE(net1099),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit30.Q ));
 sg13g2_dlhq_1 _2694_ (.D(net1135),
    .GATE(net1100),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit31.Q ));
 sg13g2_dlhq_1 _2695_ (.D(net1208),
    .GATE(net1108),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit0.Q ));
 sg13g2_dlhq_1 _2696_ (.D(net1174),
    .GATE(net1108),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit1.Q ));
 sg13g2_dlhq_1 _2697_ (.D(net1143),
    .GATE(net1104),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit2.Q ));
 sg13g2_dlhq_1 _2698_ (.D(net1134),
    .GATE(net1103),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit3.Q ));
 sg13g2_dlhq_1 _2699_ (.D(net1131),
    .GATE(net1103),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit4.Q ));
 sg13g2_dlhq_1 _2700_ (.D(net1126),
    .GATE(net1105),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit5.Q ));
 sg13g2_dlhq_1 _2701_ (.D(net1124),
    .GATE(net1105),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit6.Q ));
 sg13g2_dlhq_1 _2702_ (.D(net1121),
    .GATE(net1107),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit7.Q ));
 sg13g2_dlhq_1 _2703_ (.D(net1117),
    .GATE(net1106),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit8.Q ));
 sg13g2_dlhq_1 _2704_ (.D(net1114),
    .GATE(net1104),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit9.Q ));
 sg13g2_dlhq_1 _2705_ (.D(net1204),
    .GATE(net1104),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit10.Q ));
 sg13g2_dlhq_1 _2706_ (.D(net1202),
    .GATE(net1104),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit11.Q ));
 sg13g2_dlhq_1 _2707_ (.D(net1199),
    .GATE(net1103),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit12.Q ));
 sg13g2_dlhq_1 _2708_ (.D(net1196),
    .GATE(net1103),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit13.Q ));
 sg13g2_dlhq_1 _2709_ (.D(net1193),
    .GATE(net1103),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit14.Q ));
 sg13g2_dlhq_1 _2710_ (.D(net1190),
    .GATE(net1105),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit15.Q ));
 sg13g2_dlhq_1 _2711_ (.D(net1187),
    .GATE(net1105),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit16.Q ));
 sg13g2_dlhq_1 _2712_ (.D(net1184),
    .GATE(net1107),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit17.Q ));
 sg13g2_dlhq_1 _2713_ (.D(net1181),
    .GATE(net1106),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit18.Q ));
 sg13g2_dlhq_1 _2714_ (.D(net1178),
    .GATE(net1103),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit19.Q ));
 sg13g2_dlhq_1 _2715_ (.D(net1172),
    .GATE(net1103),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit20.Q ));
 sg13g2_dlhq_1 _2716_ (.D(net1169),
    .GATE(net1103),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit21.Q ));
 sg13g2_dlhq_1 _2717_ (.D(net1166),
    .GATE(net1106),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit22.Q ));
 sg13g2_dlhq_1 _2718_ (.D(net1163),
    .GATE(net1106),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit23.Q ));
 sg13g2_dlhq_1 _2719_ (.D(net1161),
    .GATE(net1106),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit24.Q ));
 sg13g2_dlhq_1 _2720_ (.D(net1157),
    .GATE(net1107),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit25.Q ));
 sg13g2_dlhq_1 _2721_ (.D(net1153),
    .GATE(net1107),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit26.Q ));
 sg13g2_dlhq_1 _2722_ (.D(net1151),
    .GATE(net1106),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit27.Q ));
 sg13g2_dlhq_1 _2723_ (.D(net1148),
    .GATE(net1107),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit28.Q ));
 sg13g2_dlhq_1 _2724_ (.D(net1144),
    .GATE(net1104),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit29.Q ));
 sg13g2_dlhq_1 _2725_ (.D(net1139),
    .GATE(net1104),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit30.Q ));
 sg13g2_dlhq_1 _2726_ (.D(net1136),
    .GATE(net1106),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit31.Q ));
 sg13g2_dlhq_1 _2727_ (.D(net1208),
    .GATE(net1014),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit0.Q ));
 sg13g2_dlhq_1 _2728_ (.D(net1176),
    .GATE(net1011),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit1.Q ));
 sg13g2_dlhq_1 _2729_ (.D(net1142),
    .GATE(net1011),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit2.Q ));
 sg13g2_dlhq_1 _2730_ (.D(net1134),
    .GATE(net1012),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit3.Q ));
 sg13g2_dlhq_1 _2731_ (.D(net1130),
    .GATE(net1012),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit4.Q ));
 sg13g2_dlhq_1 _2732_ (.D(net1128),
    .GATE(net1012),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit5.Q ));
 sg13g2_dlhq_1 _2733_ (.D(net1124),
    .GATE(net1012),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit6.Q ));
 sg13g2_dlhq_1 _2734_ (.D(net1121),
    .GATE(net1011),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit7.Q ));
 sg13g2_dlhq_1 _2735_ (.D(net1117),
    .GATE(net1011),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit8.Q ));
 sg13g2_dlhq_1 _2736_ (.D(net1115),
    .GATE(net1014),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit9.Q ));
 sg13g2_dlhq_1 _2737_ (.D(net1204),
    .GATE(net1013),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit10.Q ));
 sg13g2_dlhq_1 _2738_ (.D(net1202),
    .GATE(net1014),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit11.Q ));
 sg13g2_dlhq_1 _2739_ (.D(net1199),
    .GATE(net1014),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit12.Q ));
 sg13g2_dlhq_1 _2740_ (.D(net1196),
    .GATE(net1013),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit13.Q ));
 sg13g2_dlhq_1 _2741_ (.D(net1193),
    .GATE(net1013),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit14.Q ));
 sg13g2_dlhq_1 _2742_ (.D(net1190),
    .GATE(net1014),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit15.Q ));
 sg13g2_dlhq_1 _2743_ (.D(net1188),
    .GATE(net1014),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit16.Q ));
 sg13g2_dlhq_1 _2744_ (.D(net1184),
    .GATE(net1011),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit17.Q ));
 sg13g2_dlhq_1 _2745_ (.D(net1181),
    .GATE(net1011),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit18.Q ));
 sg13g2_dlhq_1 _2746_ (.D(net1178),
    .GATE(net1013),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit19.Q ));
 sg13g2_dlhq_1 _2747_ (.D(net1172),
    .GATE(net1015),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit20.Q ));
 sg13g2_dlhq_1 _2748_ (.D(net1170),
    .GATE(net1015),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit21.Q ));
 sg13g2_dlhq_1 _2749_ (.D(net1167),
    .GATE(net1013),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit22.Q ));
 sg13g2_dlhq_1 _2750_ (.D(net1163),
    .GATE(net1013),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit23.Q ));
 sg13g2_dlhq_1 _2751_ (.D(net1160),
    .GATE(net1013),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit24.Q ));
 sg13g2_dlhq_1 _2752_ (.D(net1157),
    .GATE(net1013),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit25.Q ));
 sg13g2_dlhq_1 _2753_ (.D(net1154),
    .GATE(net1014),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit26.Q ));
 sg13g2_dlhq_1 _2754_ (.D(net1150),
    .GATE(net1011),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit27.Q ));
 sg13g2_dlhq_1 _2755_ (.D(net1147),
    .GATE(net1011),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit28.Q ));
 sg13g2_dlhq_1 _2756_ (.D(net1145),
    .GATE(net1015),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit29.Q ));
 sg13g2_dlhq_1 _2757_ (.D(net1140),
    .GATE(net1015),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit30.Q ));
 sg13g2_dlhq_1 _2758_ (.D(net1137),
    .GATE(net1015),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit31.Q ));
 sg13g2_dlhq_1 _2759_ (.D(net1208),
    .GATE(net1017),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit0.Q ));
 sg13g2_dlhq_1 _2760_ (.D(net1176),
    .GATE(net1017),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit1.Q ));
 sg13g2_dlhq_1 _2761_ (.D(net1141),
    .GATE(net1017),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit2.Q ));
 sg13g2_dlhq_1 _2762_ (.D(net1132),
    .GATE(net1018),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit3.Q ));
 sg13g2_dlhq_1 _2763_ (.D(net1130),
    .GATE(net1018),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit4.Q ));
 sg13g2_dlhq_1 _2764_ (.D(net1126),
    .GATE(net1016),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit5.Q ));
 sg13g2_dlhq_1 _2765_ (.D(net1124),
    .GATE(net1016),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit6.Q ));
 sg13g2_dlhq_1 _2766_ (.D(net1121),
    .GATE(net1018),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit7.Q ));
 sg13g2_dlhq_1 _2767_ (.D(net1117),
    .GATE(net1018),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit8.Q ));
 sg13g2_dlhq_1 _2768_ (.D(net1115),
    .GATE(net1017),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit9.Q ));
 sg13g2_dlhq_1 _2769_ (.D(net1204),
    .GATE(net1017),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit10.Q ));
 sg13g2_dlhq_1 _2770_ (.D(net1203),
    .GATE(net1017),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit11.Q ));
 sg13g2_dlhq_1 _2771_ (.D(net1199),
    .GATE(net1017),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit12.Q ));
 sg13g2_dlhq_1 _2772_ (.D(net1197),
    .GATE(net1018),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit13.Q ));
 sg13g2_dlhq_1 _2773_ (.D(net1194),
    .GATE(net1018),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit14.Q ));
 sg13g2_dlhq_1 _2774_ (.D(net1190),
    .GATE(net1020),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit15.Q ));
 sg13g2_dlhq_1 _2775_ (.D(net1187),
    .GATE(net1016),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit16.Q ));
 sg13g2_dlhq_1 _2776_ (.D(net1184),
    .GATE(net1017),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit17.Q ));
 sg13g2_dlhq_1 _2777_ (.D(net1182),
    .GATE(net1019),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit18.Q ));
 sg13g2_dlhq_1 _2778_ (.D(net1179),
    .GATE(net1019),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit19.Q ));
 sg13g2_dlhq_1 _2779_ (.D(net1173),
    .GATE(net1019),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit20.Q ));
 sg13g2_dlhq_1 _2780_ (.D(net1170),
    .GATE(net1019),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit21.Q ));
 sg13g2_dlhq_1 _2781_ (.D(net1165),
    .GATE(net1019),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit22.Q ));
 sg13g2_dlhq_1 _2782_ (.D(net1164),
    .GATE(net1019),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit23.Q ));
 sg13g2_dlhq_1 _2783_ (.D(net1161),
    .GATE(net1019),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit24.Q ));
 sg13g2_dlhq_1 _2784_ (.D(net1158),
    .GATE(net1019),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit25.Q ));
 sg13g2_dlhq_1 _2785_ (.D(net1153),
    .GATE(net1020),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit26.Q ));
 sg13g2_dlhq_1 _2786_ (.D(net1150),
    .GATE(net1016),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit27.Q ));
 sg13g2_dlhq_1 _2787_ (.D(net1147),
    .GATE(net1016),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit28.Q ));
 sg13g2_dlhq_1 _2788_ (.D(net1144),
    .GATE(net1016),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit29.Q ));
 sg13g2_dlhq_1 _2789_ (.D(net1138),
    .GATE(net1016),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit30.Q ));
 sg13g2_dlhq_1 _2790_ (.D(net1136),
    .GATE(net1016),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit31.Q ));
 sg13g2_dlhq_1 _2791_ (.D(net1207),
    .GATE(net1021),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit0.Q ));
 sg13g2_dlhq_1 _2792_ (.D(net1174),
    .GATE(net1021),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit1.Q ));
 sg13g2_dlhq_1 _2793_ (.D(net1141),
    .GATE(net1024),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit2.Q ));
 sg13g2_dlhq_1 _2794_ (.D(net1132),
    .GATE(net1024),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit3.Q ));
 sg13g2_dlhq_1 _2795_ (.D(net1129),
    .GATE(net1022),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit4.Q ));
 sg13g2_dlhq_1 _2796_ (.D(net1126),
    .GATE(net30),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit5.Q ));
 sg13g2_dlhq_1 _2797_ (.D(net1125),
    .GATE(net1023),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit6.Q ));
 sg13g2_dlhq_1 _2798_ (.D(net1122),
    .GATE(net1023),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit7.Q ));
 sg13g2_dlhq_1 _2799_ (.D(net1119),
    .GATE(net1022),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit8.Q ));
 sg13g2_dlhq_1 _2800_ (.D(net1114),
    .GATE(net1022),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit9.Q ));
 sg13g2_dlhq_1 _2801_ (.D(net1206),
    .GATE(net1023),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit10.Q ));
 sg13g2_dlhq_1 _2802_ (.D(net1201),
    .GATE(net1023),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit11.Q ));
 sg13g2_dlhq_1 _2803_ (.D(net1200),
    .GATE(net1023),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit12.Q ));
 sg13g2_dlhq_1 _2804_ (.D(net1195),
    .GATE(net1024),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit13.Q ));
 sg13g2_dlhq_1 _2805_ (.D(net1192),
    .GATE(net1023),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit14.Q ));
 sg13g2_dlhq_1 _2806_ (.D(net1189),
    .GATE(net1023),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit15.Q ));
 sg13g2_dlhq_1 _2807_ (.D(net1187),
    .GATE(net1021),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit16.Q ));
 sg13g2_dlhq_1 _2808_ (.D(net1184),
    .GATE(net1021),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit17.Q ));
 sg13g2_dlhq_1 _2809_ (.D(net1180),
    .GATE(net1025),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit18.Q ));
 sg13g2_dlhq_1 _2810_ (.D(net1178),
    .GATE(net1025),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit19.Q ));
 sg13g2_dlhq_1 _2811_ (.D(net1173),
    .GATE(net1025),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit20.Q ));
 sg13g2_dlhq_1 _2812_ (.D(net1168),
    .GATE(net1025),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit21.Q ));
 sg13g2_dlhq_1 _2813_ (.D(net1167),
    .GATE(net1024),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit22.Q ));
 sg13g2_dlhq_1 _2814_ (.D(net1164),
    .GATE(net1023),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit23.Q ));
 sg13g2_dlhq_1 _2815_ (.D(net1159),
    .GATE(net1021),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit24.Q ));
 sg13g2_dlhq_1 _2816_ (.D(net1156),
    .GATE(net1021),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit25.Q ));
 sg13g2_dlhq_1 _2817_ (.D(net1153),
    .GATE(net1022),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit26.Q ));
 sg13g2_dlhq_1 _2818_ (.D(net1150),
    .GATE(net1022),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit27.Q ));
 sg13g2_dlhq_1 _2819_ (.D(net1147),
    .GATE(net1021),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit28.Q ));
 sg13g2_dlhq_1 _2820_ (.D(net1144),
    .GATE(net1021),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit29.Q ));
 sg13g2_dlhq_1 _2821_ (.D(net1139),
    .GATE(net1022),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit30.Q ));
 sg13g2_dlhq_1 _2822_ (.D(net1136),
    .GATE(net1022),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit31.Q ));
 sg13g2_dlhq_1 _2823_ (.D(net1207),
    .GATE(net1027),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit0.Q ));
 sg13g2_dlhq_1 _2824_ (.D(net1175),
    .GATE(net1026),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit1.Q ));
 sg13g2_dlhq_1 _2825_ (.D(net1143),
    .GATE(net1029),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit2.Q ));
 sg13g2_dlhq_1 _2826_ (.D(net1134),
    .GATE(net1029),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit3.Q ));
 sg13g2_dlhq_1 _2827_ (.D(net1131),
    .GATE(net1026),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit4.Q ));
 sg13g2_dlhq_1 _2828_ (.D(net1126),
    .GATE(net1026),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit5.Q ));
 sg13g2_dlhq_1 _2829_ (.D(net1124),
    .GATE(net1030),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit6.Q ));
 sg13g2_dlhq_1 _2830_ (.D(net1121),
    .GATE(net1030),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit7.Q ));
 sg13g2_dlhq_1 _2831_ (.D(net1117),
    .GATE(net1027),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit8.Q ));
 sg13g2_dlhq_1 _2832_ (.D(net1114),
    .GATE(net1027),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit9.Q ));
 sg13g2_dlhq_1 _2833_ (.D(net1204),
    .GATE(net1029),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit10.Q ));
 sg13g2_dlhq_1 _2834_ (.D(net1202),
    .GATE(net1029),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit11.Q ));
 sg13g2_dlhq_1 _2835_ (.D(net1198),
    .GATE(net1026),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit12.Q ));
 sg13g2_dlhq_1 _2836_ (.D(net1196),
    .GATE(net1026),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit13.Q ));
 sg13g2_dlhq_1 _2837_ (.D(net1193),
    .GATE(net1030),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit14.Q ));
 sg13g2_dlhq_1 _2838_ (.D(net1190),
    .GATE(net1030),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit15.Q ));
 sg13g2_dlhq_1 _2839_ (.D(net1187),
    .GATE(net1026),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit16.Q ));
 sg13g2_dlhq_1 _2840_ (.D(net1184),
    .GATE(net1026),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit17.Q ));
 sg13g2_dlhq_1 _2841_ (.D(net1181),
    .GATE(net1029),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit18.Q ));
 sg13g2_dlhq_1 _2842_ (.D(net1178),
    .GATE(net1029),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit19.Q ));
 sg13g2_dlhq_1 _2843_ (.D(net1171),
    .GATE(net1028),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit20.Q ));
 sg13g2_dlhq_1 _2844_ (.D(net1169),
    .GATE(net1028),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit21.Q ));
 sg13g2_dlhq_1 _2845_ (.D(net1167),
    .GATE(net1030),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit22.Q ));
 sg13g2_dlhq_1 _2846_ (.D(net1163),
    .GATE(net1030),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit23.Q ));
 sg13g2_dlhq_1 _2847_ (.D(net1160),
    .GATE(net1027),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit24.Q ));
 sg13g2_dlhq_1 _2848_ (.D(net1157),
    .GATE(net1026),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit25.Q ));
 sg13g2_dlhq_1 _2849_ (.D(net1154),
    .GATE(net1029),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit26.Q ));
 sg13g2_dlhq_1 _2850_ (.D(net1151),
    .GATE(net1029),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit27.Q ));
 sg13g2_dlhq_1 _2851_ (.D(net1149),
    .GATE(net1031),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit28.Q ));
 sg13g2_dlhq_1 _2852_ (.D(net1146),
    .GATE(net1031),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit29.Q ));
 sg13g2_dlhq_1 _2853_ (.D(net1139),
    .GATE(net1031),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit30.Q ));
 sg13g2_dlhq_1 _2854_ (.D(net1136),
    .GATE(net1031),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit31.Q ));
 sg13g2_dlhq_1 _2855_ (.D(net1208),
    .GATE(net1034),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit0.Q ));
 sg13g2_dlhq_1 _2856_ (.D(net26),
    .GATE(net1034),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit1.Q ));
 sg13g2_dlhq_1 _2857_ (.D(net1141),
    .GATE(net1034),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit2.Q ));
 sg13g2_dlhq_1 _2858_ (.D(net1132),
    .GATE(net1034),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit3.Q ));
 sg13g2_dlhq_1 _2859_ (.D(net1131),
    .GATE(net29),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit4.Q ));
 sg13g2_dlhq_1 _2860_ (.D(net1126),
    .GATE(net1034),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit5.Q ));
 sg13g2_dlhq_1 _2861_ (.D(net1123),
    .GATE(net1033),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit6.Q ));
 sg13g2_dlhq_1 _2862_ (.D(net1120),
    .GATE(net1033),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit7.Q ));
 sg13g2_dlhq_1 _2863_ (.D(net1119),
    .GATE(net1034),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit8.Q ));
 sg13g2_dlhq_1 _2864_ (.D(net1116),
    .GATE(net1034),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit9.Q ));
 sg13g2_dlhq_1 _2865_ (.D(net1206),
    .GATE(net1035),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit10.Q ));
 sg13g2_dlhq_1 _2866_ (.D(net1203),
    .GATE(net1035),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit11.Q ));
 sg13g2_dlhq_1 _2867_ (.D(net1200),
    .GATE(net1035),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit12.Q ));
 sg13g2_dlhq_1 _2868_ (.D(net1195),
    .GATE(net1035),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit13.Q ));
 sg13g2_dlhq_1 _2869_ (.D(net1192),
    .GATE(net1036),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit14.Q ));
 sg13g2_dlhq_1 _2870_ (.D(net1189),
    .GATE(net1036),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit15.Q ));
 sg13g2_dlhq_1 _2871_ (.D(net1186),
    .GATE(net1032),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit16.Q ));
 sg13g2_dlhq_1 _2872_ (.D(net1183),
    .GATE(net1032),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit17.Q ));
 sg13g2_dlhq_1 _2873_ (.D(net1180),
    .GATE(net1035),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit18.Q ));
 sg13g2_dlhq_1 _2874_ (.D(net1177),
    .GATE(net1035),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit19.Q ));
 sg13g2_dlhq_1 _2875_ (.D(net1173),
    .GATE(net1035),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit20.Q ));
 sg13g2_dlhq_1 _2876_ (.D(net1170),
    .GATE(net1035),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit21.Q ));
 sg13g2_dlhq_1 _2877_ (.D(net1165),
    .GATE(net1036),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit22.Q ));
 sg13g2_dlhq_1 _2878_ (.D(net1162),
    .GATE(net1036),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit23.Q ));
 sg13g2_dlhq_1 _2879_ (.D(net1159),
    .GATE(net1033),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit24.Q ));
 sg13g2_dlhq_1 _2880_ (.D(net1156),
    .GATE(net1032),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit25.Q ));
 sg13g2_dlhq_1 _2881_ (.D(net1155),
    .GATE(net1032),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit26.Q ));
 sg13g2_dlhq_1 _2882_ (.D(net1152),
    .GATE(net1032),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit27.Q ));
 sg13g2_dlhq_1 _2883_ (.D(net1149),
    .GATE(net1032),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit28.Q ));
 sg13g2_dlhq_1 _2884_ (.D(net1146),
    .GATE(net1032),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit29.Q ));
 sg13g2_dlhq_1 _2885_ (.D(net1138),
    .GATE(net1032),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit30.Q ));
 sg13g2_dlhq_1 _2886_ (.D(net1135),
    .GATE(net1033),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit31.Q ));
 sg13g2_dlhq_1 _2887_ (.D(net1207),
    .GATE(net1038),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit0.Q ));
 sg13g2_dlhq_1 _2888_ (.D(net1174),
    .GATE(net1038),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit1.Q ));
 sg13g2_dlhq_1 _2889_ (.D(net1141),
    .GATE(net1041),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit2.Q ));
 sg13g2_dlhq_1 _2890_ (.D(net1132),
    .GATE(net1041),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit3.Q ));
 sg13g2_dlhq_1 _2891_ (.D(net1129),
    .GATE(net1041),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit4.Q ));
 sg13g2_dlhq_1 _2892_ (.D(net1127),
    .GATE(net1041),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit5.Q ));
 sg13g2_dlhq_1 _2893_ (.D(net1123),
    .GATE(net1037),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit6.Q ));
 sg13g2_dlhq_1 _2894_ (.D(net1120),
    .GATE(net1037),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit7.Q ));
 sg13g2_dlhq_1 _2895_ (.D(net1119),
    .GATE(net1037),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit8.Q ));
 sg13g2_dlhq_1 _2896_ (.D(net1116),
    .GATE(net1037),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit9.Q ));
 sg13g2_dlhq_1 _2897_ (.D(net1206),
    .GATE(net1039),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit10.Q ));
 sg13g2_dlhq_1 _2898_ (.D(net1201),
    .GATE(net1039),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit11.Q ));
 sg13g2_dlhq_1 _2899_ (.D(net1198),
    .GATE(net1039),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit12.Q ));
 sg13g2_dlhq_1 _2900_ (.D(net1197),
    .GATE(net1039),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit13.Q ));
 sg13g2_dlhq_1 _2901_ (.D(net1192),
    .GATE(net1039),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit14.Q ));
 sg13g2_dlhq_1 _2902_ (.D(net1189),
    .GATE(net1040),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit15.Q ));
 sg13g2_dlhq_1 _2903_ (.D(net1186),
    .GATE(net1040),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit16.Q ));
 sg13g2_dlhq_1 _2904_ (.D(net1183),
    .GATE(net1040),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit17.Q ));
 sg13g2_dlhq_1 _2905_ (.D(net1180),
    .GATE(net1041),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit18.Q ));
 sg13g2_dlhq_1 _2906_ (.D(net1177),
    .GATE(net1039),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit19.Q ));
 sg13g2_dlhq_1 _2907_ (.D(net1171),
    .GATE(net1039),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit20.Q ));
 sg13g2_dlhq_1 _2908_ (.D(net1168),
    .GATE(net1039),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit21.Q ));
 sg13g2_dlhq_1 _2909_ (.D(net1165),
    .GATE(net1040),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit22.Q ));
 sg13g2_dlhq_1 _2910_ (.D(net1162),
    .GATE(net1040),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit23.Q ));
 sg13g2_dlhq_1 _2911_ (.D(net1161),
    .GATE(net1040),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit24.Q ));
 sg13g2_dlhq_1 _2912_ (.D(net1156),
    .GATE(net1040),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit25.Q ));
 sg13g2_dlhq_1 _2913_ (.D(net1155),
    .GATE(net1037),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit26.Q ));
 sg13g2_dlhq_1 _2914_ (.D(net1152),
    .GATE(net1037),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit27.Q ));
 sg13g2_dlhq_1 _2915_ (.D(net1149),
    .GATE(net1037),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit28.Q ));
 sg13g2_dlhq_1 _2916_ (.D(net1146),
    .GATE(net1037),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit29.Q ));
 sg13g2_dlhq_1 _2917_ (.D(net1138),
    .GATE(net1038),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit30.Q ));
 sg13g2_dlhq_1 _2918_ (.D(net1135),
    .GATE(net1038),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit31.Q ));
 sg13g2_dlhq_1 _2919_ (.D(net1207),
    .GATE(net1046),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit0.Q ));
 sg13g2_dlhq_1 _2920_ (.D(net1174),
    .GATE(net1043),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit1.Q ));
 sg13g2_dlhq_1 _2921_ (.D(net1143),
    .GATE(net1043),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit2.Q ));
 sg13g2_dlhq_1 _2922_ (.D(net1134),
    .GATE(net1043),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit3.Q ));
 sg13g2_dlhq_1 _2923_ (.D(net1131),
    .GATE(net1043),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit4.Q ));
 sg13g2_dlhq_1 _2924_ (.D(net1126),
    .GATE(net1043),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit5.Q ));
 sg13g2_dlhq_1 _2925_ (.D(net1123),
    .GATE(net1042),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit6.Q ));
 sg13g2_dlhq_1 _2926_ (.D(net1120),
    .GATE(net1042),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit7.Q ));
 sg13g2_dlhq_1 _2927_ (.D(net1119),
    .GATE(net1042),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit8.Q ));
 sg13g2_dlhq_1 _2928_ (.D(net1116),
    .GATE(net1042),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit9.Q ));
 sg13g2_dlhq_1 _2929_ (.D(net1206),
    .GATE(net1045),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit10.Q ));
 sg13g2_dlhq_1 _2930_ (.D(net1201),
    .GATE(net1045),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit11.Q ));
 sg13g2_dlhq_1 _2931_ (.D(net1198),
    .GATE(net1045),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit12.Q ));
 sg13g2_dlhq_1 _2932_ (.D(net1197),
    .GATE(net1045),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit13.Q ));
 sg13g2_dlhq_1 _2933_ (.D(net1192),
    .GATE(net1045),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit14.Q ));
 sg13g2_dlhq_1 _2934_ (.D(net1189),
    .GATE(net1045),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit15.Q ));
 sg13g2_dlhq_1 _2935_ (.D(net1186),
    .GATE(net1046),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit16.Q ));
 sg13g2_dlhq_1 _2936_ (.D(net1183),
    .GATE(net1044),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit17.Q ));
 sg13g2_dlhq_1 _2937_ (.D(net1180),
    .GATE(net1045),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit18.Q ));
 sg13g2_dlhq_1 _2938_ (.D(net1177),
    .GATE(net1045),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit19.Q ));
 sg13g2_dlhq_1 _2939_ (.D(net1171),
    .GATE(net1044),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit20.Q ));
 sg13g2_dlhq_1 _2940_ (.D(net1168),
    .GATE(net1044),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit21.Q ));
 sg13g2_dlhq_1 _2941_ (.D(net1165),
    .GATE(net1044),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit22.Q ));
 sg13g2_dlhq_1 _2942_ (.D(net1162),
    .GATE(net1044),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit23.Q ));
 sg13g2_dlhq_1 _2943_ (.D(net1159),
    .GATE(net1044),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit24.Q ));
 sg13g2_dlhq_1 _2944_ (.D(net1156),
    .GATE(net1044),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit25.Q ));
 sg13g2_dlhq_1 _2945_ (.D(net1155),
    .GATE(net1043),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit26.Q ));
 sg13g2_dlhq_1 _2946_ (.D(net1152),
    .GATE(net1042),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit27.Q ));
 sg13g2_dlhq_1 _2947_ (.D(net1149),
    .GATE(net1042),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit28.Q ));
 sg13g2_dlhq_1 _2948_ (.D(net1146),
    .GATE(net1042),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit29.Q ));
 sg13g2_dlhq_1 _2949_ (.D(net1138),
    .GATE(net1043),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit30.Q ));
 sg13g2_dlhq_1 _2950_ (.D(net1135),
    .GATE(net1042),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit31.Q ));
 sg13g2_dlhq_1 _2951_ (.D(net1207),
    .GATE(net1048),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit0.Q ));
 sg13g2_dlhq_1 _2952_ (.D(net1174),
    .GATE(net1048),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit1.Q ));
 sg13g2_dlhq_1 _2953_ (.D(net1141),
    .GATE(net1049),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit2.Q ));
 sg13g2_dlhq_1 _2954_ (.D(net1132),
    .GATE(net1050),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit3.Q ));
 sg13g2_dlhq_1 _2955_ (.D(net1129),
    .GATE(net1052),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit4.Q ));
 sg13g2_dlhq_1 _2956_ (.D(net1127),
    .GATE(net1049),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit5.Q ));
 sg13g2_dlhq_1 _2957_ (.D(net1123),
    .GATE(net1047),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit6.Q ));
 sg13g2_dlhq_1 _2958_ (.D(net1120),
    .GATE(net1047),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit7.Q ));
 sg13g2_dlhq_1 _2959_ (.D(net1119),
    .GATE(net1047),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit8.Q ));
 sg13g2_dlhq_1 _2960_ (.D(net1116),
    .GATE(net1047),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit9.Q ));
 sg13g2_dlhq_1 _2961_ (.D(net1206),
    .GATE(net1051),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit10.Q ));
 sg13g2_dlhq_1 _2962_ (.D(net1201),
    .GATE(net1051),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit11.Q ));
 sg13g2_dlhq_1 _2963_ (.D(net1200),
    .GATE(net1051),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit12.Q ));
 sg13g2_dlhq_1 _2964_ (.D(net1195),
    .GATE(net1050),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit13.Q ));
 sg13g2_dlhq_1 _2965_ (.D(net1192),
    .GATE(net1050),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit14.Q ));
 sg13g2_dlhq_1 _2966_ (.D(net1189),
    .GATE(net1050),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit15.Q ));
 sg13g2_dlhq_1 _2967_ (.D(net1186),
    .GATE(net1050),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit16.Q ));
 sg13g2_dlhq_1 _2968_ (.D(net1183),
    .GATE(net1050),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit17.Q ));
 sg13g2_dlhq_1 _2969_ (.D(net1180),
    .GATE(net1050),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit18.Q ));
 sg13g2_dlhq_1 _2970_ (.D(net1177),
    .GATE(net1050),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit19.Q ));
 sg13g2_dlhq_1 _2971_ (.D(net1171),
    .GATE(net1051),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit20.Q ));
 sg13g2_dlhq_1 _2972_ (.D(net1168),
    .GATE(net1051),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit21.Q ));
 sg13g2_dlhq_1 _2973_ (.D(net1165),
    .GATE(net1049),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit22.Q ));
 sg13g2_dlhq_1 _2974_ (.D(net1162),
    .GATE(net1049),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit23.Q ));
 sg13g2_dlhq_1 _2975_ (.D(net1159),
    .GATE(net1049),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit24.Q ));
 sg13g2_dlhq_1 _2976_ (.D(net1156),
    .GATE(net1049),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit25.Q ));
 sg13g2_dlhq_1 _2977_ (.D(net1155),
    .GATE(net1047),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit26.Q ));
 sg13g2_dlhq_1 _2978_ (.D(net1152),
    .GATE(net1047),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit27.Q ));
 sg13g2_dlhq_1 _2979_ (.D(net1149),
    .GATE(net1047),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit28.Q ));
 sg13g2_dlhq_1 _2980_ (.D(net1146),
    .GATE(net1047),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit29.Q ));
 sg13g2_dlhq_1 _2981_ (.D(net1138),
    .GATE(net1048),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit30.Q ));
 sg13g2_dlhq_1 _2982_ (.D(net1135),
    .GATE(net1048),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit31.Q ));
 sg13g2_dlhq_1 _2983_ (.D(net1207),
    .GATE(net1053),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit0.Q ));
 sg13g2_dlhq_1 _2984_ (.D(net1174),
    .GATE(net1053),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit1.Q ));
 sg13g2_dlhq_1 _2985_ (.D(net1143),
    .GATE(net1054),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit2.Q ));
 sg13g2_dlhq_1 _2986_ (.D(net1134),
    .GATE(net1054),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit3.Q ));
 sg13g2_dlhq_1 _2987_ (.D(net1131),
    .GATE(net1053),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit4.Q ));
 sg13g2_dlhq_1 _2988_ (.D(net1126),
    .GATE(net1053),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit5.Q ));
 sg13g2_dlhq_1 _2989_ (.D(net1123),
    .GATE(net1053),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit6.Q ));
 sg13g2_dlhq_1 _2990_ (.D(net1120),
    .GATE(net1053),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit7.Q ));
 sg13g2_dlhq_1 _2991_ (.D(net1119),
    .GATE(net1053),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit8.Q ));
 sg13g2_dlhq_1 _2992_ (.D(net1116),
    .GATE(net1053),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit9.Q ));
 sg13g2_dlhq_1 _2993_ (.D(net1206),
    .GATE(net1056),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit10.Q ));
 sg13g2_dlhq_1 _2994_ (.D(net1201),
    .GATE(net1056),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit11.Q ));
 sg13g2_dlhq_1 _2995_ (.D(net1198),
    .GATE(net1056),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit12.Q ));
 sg13g2_dlhq_1 _2996_ (.D(net1195),
    .GATE(net1056),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit13.Q ));
 sg13g2_dlhq_1 _2997_ (.D(net1192),
    .GATE(net1056),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit14.Q ));
 sg13g2_dlhq_1 _2998_ (.D(net1189),
    .GATE(net1056),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit15.Q ));
 sg13g2_dlhq_1 _2999_ (.D(net1186),
    .GATE(net1056),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit16.Q ));
 sg13g2_dlhq_1 _3000_ (.D(net1183),
    .GATE(net1056),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit17.Q ));
 sg13g2_dlhq_1 _3001_ (.D(net1182),
    .GATE(net1057),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit18.Q ));
 sg13g2_dlhq_1 _3002_ (.D(net1177),
    .GATE(net1057),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit19.Q ));
 sg13g2_dlhq_1 _3003_ (.D(net1171),
    .GATE(net1057),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit20.Q ));
 sg13g2_dlhq_1 _3004_ (.D(net1168),
    .GATE(net1057),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit21.Q ));
 sg13g2_dlhq_1 _3005_ (.D(net1165),
    .GATE(net1055),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit22.Q ));
 sg13g2_dlhq_1 _3006_ (.D(net1162),
    .GATE(net1054),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit23.Q ));
 sg13g2_dlhq_1 _3007_ (.D(net1159),
    .GATE(net1054),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit24.Q ));
 sg13g2_dlhq_1 _3008_ (.D(net1156),
    .GATE(net1054),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit25.Q ));
 sg13g2_dlhq_1 _3009_ (.D(net1153),
    .GATE(net1055),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit26.Q ));
 sg13g2_dlhq_1 _3010_ (.D(net1152),
    .GATE(net1055),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit27.Q ));
 sg13g2_dlhq_1 _3011_ (.D(net1147),
    .GATE(net1055),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit28.Q ));
 sg13g2_dlhq_1 _3012_ (.D(net1144),
    .GATE(net1055),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit29.Q ));
 sg13g2_dlhq_1 _3013_ (.D(net1138),
    .GATE(net1054),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit30.Q ));
 sg13g2_dlhq_1 _3014_ (.D(net1135),
    .GATE(net1054),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit31.Q ));
 sg13g2_dlhq_1 _3015_ (.D(net1207),
    .GATE(net1109),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit0.Q ));
 sg13g2_dlhq_1 _3016_ (.D(net1174),
    .GATE(net1109),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit1.Q ));
 sg13g2_dlhq_1 _3017_ (.D(net1143),
    .GATE(net1111),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit2.Q ));
 sg13g2_dlhq_1 _3018_ (.D(net1134),
    .GATE(net1111),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit3.Q ));
 sg13g2_dlhq_1 _3019_ (.D(net1131),
    .GATE(net1111),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit4.Q ));
 sg13g2_dlhq_1 _3020_ (.D(net1126),
    .GATE(net1111),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit5.Q ));
 sg13g2_dlhq_1 _3021_ (.D(net1123),
    .GATE(net1111),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit6.Q ));
 sg13g2_dlhq_1 _3022_ (.D(net1120),
    .GATE(net1111),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit7.Q ));
 sg13g2_dlhq_1 _3023_ (.D(net1117),
    .GATE(net1110),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit8.Q ));
 sg13g2_dlhq_1 _3024_ (.D(net1114),
    .GATE(net1110),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit9.Q ));
 sg13g2_dlhq_1 _3025_ (.D(net1204),
    .GATE(net1113),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit10.Q ));
 sg13g2_dlhq_1 _3026_ (.D(net1203),
    .GATE(net1113),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit11.Q ));
 sg13g2_dlhq_1 _3027_ (.D(net1198),
    .GATE(net1109),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit12.Q ));
 sg13g2_dlhq_1 _3028_ (.D(net1195),
    .GATE(net1109),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit13.Q ));
 sg13g2_dlhq_1 _3029_ (.D(net1192),
    .GATE(net1111),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit14.Q ));
 sg13g2_dlhq_1 _3030_ (.D(net1189),
    .GATE(net1111),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit15.Q ));
 sg13g2_dlhq_1 _3031_ (.D(net1186),
    .GATE(net1109),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit16.Q ));
 sg13g2_dlhq_1 _3032_ (.D(net1183),
    .GATE(net1109),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit17.Q ));
 sg13g2_dlhq_1 _3033_ (.D(net1181),
    .GATE(net1113),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit18.Q ));
 sg13g2_dlhq_1 _3034_ (.D(net1179),
    .GATE(net1113),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit19.Q ));
 sg13g2_dlhq_1 _3035_ (.D(net1173),
    .GATE(net1113),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit20.Q ));
 sg13g2_dlhq_1 _3036_ (.D(net1170),
    .GATE(net1113),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit21.Q ));
 sg13g2_dlhq_1 _3037_ (.D(net1167),
    .GATE(net1113),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit22.Q ));
 sg13g2_dlhq_1 _3038_ (.D(net1164),
    .GATE(net1113),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit23.Q ));
 sg13g2_dlhq_1 _3039_ (.D(net1159),
    .GATE(net1109),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit24.Q ));
 sg13g2_dlhq_1 _3040_ (.D(net1156),
    .GATE(net1109),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit25.Q ));
 sg13g2_dlhq_1 _3041_ (.D(net1153),
    .GATE(net1112),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q ));
 sg13g2_dlhq_1 _3042_ (.D(net1150),
    .GATE(net1112),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit27.Q ));
 sg13g2_dlhq_1 _3043_ (.D(net1147),
    .GATE(net1112),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit28.Q ));
 sg13g2_dlhq_1 _3044_ (.D(net1144),
    .GATE(net1110),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit29.Q ));
 sg13g2_dlhq_1 _3045_ (.D(net1139),
    .GATE(net1110),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit30.Q ));
 sg13g2_dlhq_1 _3046_ (.D(net1137),
    .GATE(net1110),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit31.Q ));
 sg13g2_dfrbp_1 _3047_ (.CLK(UserCLK),
    .RESET_B(net371),
    .D(_0000_),
    .Q_N(_1170_),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.LUT_flop ));
 sg13g2_dfrbp_1 _3048_ (.CLK(UserCLK),
    .RESET_B(net370),
    .D(_0001_),
    .Q_N(_1169_),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.LUT_flop ));
 sg13g2_dfrbp_1 _3049_ (.CLK(UserCLK),
    .RESET_B(net369),
    .D(_0002_),
    .Q_N(_1168_),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.LUT_flop ));
 sg13g2_dfrbp_1 _3050_ (.CLK(UserCLK),
    .RESET_B(net368),
    .D(_0003_),
    .Q_N(_1167_),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.LUT_flop ));
 sg13g2_dfrbp_1 _3051_ (.CLK(UserCLK),
    .RESET_B(net367),
    .D(_0004_),
    .Q_N(_1166_),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.LUT_flop ));
 sg13g2_dfrbp_1 _3052_ (.CLK(UserCLK),
    .RESET_B(net366),
    .D(_0005_),
    .Q_N(_1165_),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.LUT_flop ));
 sg13g2_dfrbp_1 _3053_ (.CLK(UserCLK),
    .RESET_B(net373),
    .D(_0006_),
    .Q_N(_1164_),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.LUT_flop ));
 sg13g2_dfrbp_1 _3054_ (.CLK(UserCLK),
    .RESET_B(net372),
    .D(_0007_),
    .Q_N(_1163_),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.LUT_flop ));
 sg13g2_tiehi _3051__367 (.L_HI(net367));
 sg13g2_tiehi _3050__368 (.L_HI(net368));
 sg13g2_tiehi _3049__369 (.L_HI(net369));
 sg13g2_tiehi _3048__370 (.L_HI(net370));
 sg13g2_tiehi _3047__371 (.L_HI(net371));
 sg13g2_tiehi _3054__372 (.L_HI(net372));
 sg13g2_tiehi _3053__373 (.L_HI(net373));
 sg13g2_dlygate4sd1_1 rebuffer1 (.A(_0565_),
    .X(net374));
 sg13g2_buf_1 _3063_ (.A(\Inst_LUT4AB_switch_matrix.E1BEG0 ),
    .X(net113));
 sg13g2_buf_1 _3064_ (.A(\Inst_LUT4AB_switch_matrix.E1BEG1 ),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold24 (.A(\Inst_LH_LUT4c_frame_config_dffesr.LUT_flop ),
    .X(net397));
 sg13g2_fill_1 FILLER_0_2 ();
 sg13g2_buf_2 _3067_ (.A(\Inst_LUT4AB_switch_matrix.E2BEG0 ),
    .X(net117));
 sg13g2_buf_1 _3068_ (.A(net382),
    .X(net118));
 sg13g2_buf_1 _3069_ (.A(\Inst_LUT4AB_switch_matrix.E2BEG2 ),
    .X(net119));
 sg13g2_buf_1 _3070_ (.A(\Inst_LUT4AB_switch_matrix.E2BEG3 ),
    .X(net120));
 sg13g2_buf_2 _3071_ (.A(\Inst_LUT4AB_switch_matrix.E2BEG4 ),
    .X(net121));
 sg13g2_fill_1 FILLER_0_197 ();
 sg13g2_buf_2 _3073_ (.A(\Inst_LUT4AB_switch_matrix.E2BEG6 ),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold23 (.A(\Inst_LE_LUT4c_frame_config_dffesr.LUT_flop ),
    .X(net396));
 sg13g2_buf_1 _3075_ (.A(net14),
    .X(net125));
 sg13g2_buf_1 _3076_ (.A(net15),
    .X(net126));
 sg13g2_buf_1 _3077_ (.A(net16),
    .X(net127));
 sg13g2_buf_1 _3078_ (.A(net17),
    .X(net128));
 sg13g2_buf_1 _3079_ (.A(net18),
    .X(net129));
 sg13g2_buf_1 _3080_ (.A(net19),
    .X(net130));
 sg13g2_buf_1 _3081_ (.A(net20),
    .X(net131));
 sg13g2_buf_1 _3082_ (.A(net21),
    .X(net132));
 sg13g2_buf_1 _3083_ (.A(E6END[2]),
    .X(net133));
 sg13g2_buf_1 _3084_ (.A(E6END[3]),
    .X(net136));
 sg13g2_buf_1 _3085_ (.A(E6END[4]),
    .X(net137));
 sg13g2_buf_1 _3086_ (.A(E6END[5]),
    .X(net138));
 sg13g2_buf_1 _3087_ (.A(E6END[6]),
    .X(net139));
 sg13g2_buf_1 _3088_ (.A(E6END[7]),
    .X(net140));
 sg13g2_buf_1 _3089_ (.A(E6END[8]),
    .X(net141));
 sg13g2_buf_1 _3090_ (.A(E6END[9]),
    .X(net142));
 sg13g2_buf_1 _3091_ (.A(E6END[10]),
    .X(net143));
 sg13g2_buf_1 _3092_ (.A(E6END[11]),
    .X(net144));
 sg13g2_buf_1 _3093_ (.A(\Inst_LUT4AB_switch_matrix.E6BEG0 ),
    .X(net134));
 sg13g2_buf_2 rebuffer13 (.A(_0479_),
    .X(net386));
 sg13g2_buf_1 _3095_ (.A(EE4END[4]),
    .X(net145));
 sg13g2_buf_1 _3096_ (.A(EE4END[5]),
    .X(net152));
 sg13g2_buf_1 _3097_ (.A(EE4END[6]),
    .X(net153));
 sg13g2_buf_1 _3098_ (.A(EE4END[7]),
    .X(net154));
 sg13g2_buf_1 _3099_ (.A(EE4END[8]),
    .X(net155));
 sg13g2_buf_1 _3100_ (.A(EE4END[9]),
    .X(net156));
 sg13g2_buf_1 _3101_ (.A(EE4END[10]),
    .X(net157));
 sg13g2_buf_1 _3102_ (.A(EE4END[11]),
    .X(net158));
 sg13g2_buf_1 _3103_ (.A(EE4END[12]),
    .X(net159));
 sg13g2_buf_1 _3104_ (.A(EE4END[13]),
    .X(net160));
 sg13g2_buf_1 _3105_ (.A(EE4END[14]),
    .X(net146));
 sg13g2_buf_1 _3106_ (.A(EE4END[15]),
    .X(net147));
 sg13g2_buf_1 _3107_ (.A(\Inst_LUT4AB_switch_matrix.EE4BEG0 ),
    .X(net148));
 sg13g2_buf_1 _3108_ (.A(\Inst_LUT4AB_switch_matrix.EE4BEG1 ),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold19 (.A(\Inst_LC_LUT4c_frame_config_dffesr.LUT_flop ),
    .X(net392));
 sg13g2_fill_1 FILLER_0_260 ();
 sg13g2_buf_1 _3111_ (.A(net1208),
    .X(net161));
 sg13g2_buf_1 _3112_ (.A(net1176),
    .X(net172));
 sg13g2_buf_1 _3113_ (.A(net1141),
    .X(net183));
 sg13g2_buf_1 _3114_ (.A(net1133),
    .X(net186));
 sg13g2_buf_1 _3115_ (.A(net1129),
    .X(net187));
 sg13g2_buf_1 _3116_ (.A(net1127),
    .X(net188));
 sg13g2_buf_1 _3117_ (.A(net1124),
    .X(net189));
 sg13g2_buf_1 _3118_ (.A(net1121),
    .X(net190));
 sg13g2_buf_1 _3119_ (.A(net1117),
    .X(net191));
 sg13g2_buf_1 _3120_ (.A(net1114),
    .X(net192));
 sg13g2_buf_1 _3121_ (.A(net1204),
    .X(net162));
 sg13g2_buf_1 _3122_ (.A(net1202),
    .X(net163));
 sg13g2_buf_1 _3123_ (.A(net1199),
    .X(net164));
 sg13g2_buf_1 _3124_ (.A(net1196),
    .X(net165));
 sg13g2_buf_1 _3125_ (.A(net1193),
    .X(net166));
 sg13g2_buf_1 _3126_ (.A(net1190),
    .X(net167));
 sg13g2_buf_1 _3127_ (.A(net1188),
    .X(net168));
 sg13g2_buf_1 _3128_ (.A(net1185),
    .X(net169));
 sg13g2_buf_1 _3129_ (.A(net1181),
    .X(net170));
 sg13g2_buf_1 _3130_ (.A(net1178),
    .X(net171));
 sg13g2_buf_1 _3131_ (.A(net1172),
    .X(net173));
 sg13g2_buf_1 _3132_ (.A(net1169),
    .X(net174));
 sg13g2_buf_1 _3133_ (.A(net1166),
    .X(net175));
 sg13g2_buf_1 _3134_ (.A(net1163),
    .X(net176));
 sg13g2_buf_1 _3135_ (.A(net1160),
    .X(net177));
 sg13g2_buf_1 _3136_ (.A(net1157),
    .X(net178));
 sg13g2_buf_1 _3137_ (.A(net1154),
    .X(net179));
 sg13g2_buf_1 _3138_ (.A(net1151),
    .X(net180));
 sg13g2_buf_1 _3139_ (.A(net1148),
    .X(net181));
 sg13g2_buf_1 _3140_ (.A(net1145),
    .X(net182));
 sg13g2_buf_1 _3141_ (.A(net1140),
    .X(net184));
 sg13g2_buf_1 _3142_ (.A(net1137),
    .X(net185));
 sg13g2_buf_1 _3143_ (.A(FrameStrobe[0]),
    .X(net193));
 sg13g2_buf_1 _3144_ (.A(net1058),
    .X(net204));
 sg13g2_buf_1 _3145_ (.A(net1052),
    .X(net205));
 sg13g2_buf_1 _3146_ (.A(net1044),
    .X(net206));
 sg13g2_buf_1 _3147_ (.A(net1041),
    .X(net207));
 sg13g2_buf_1 _3148_ (.A(net1036),
    .X(net208));
 sg13g2_buf_1 _3149_ (.A(net1030),
    .X(net209));
 sg13g2_buf_1 _3150_ (.A(net1025),
    .X(net210));
 sg13g2_buf_1 _3151_ (.A(net1018),
    .X(net211));
 sg13g2_buf_1 _3152_ (.A(net1015),
    .X(net212));
 sg13g2_buf_1 _3153_ (.A(net1106),
    .X(net194));
 sg13g2_buf_1 _3154_ (.A(net1102),
    .X(net195));
 sg13g2_buf_1 _3155_ (.A(net1097),
    .X(net196));
 sg13g2_buf_1 _3156_ (.A(net1090),
    .X(net197));
 sg13g2_buf_1 _3157_ (.A(net1084),
    .X(net198));
 sg13g2_buf_1 _3158_ (.A(net1081),
    .X(net199));
 sg13g2_buf_1 _3159_ (.A(net1075),
    .X(net200));
 sg13g2_buf_1 _3160_ (.A(FrameStrobe[17]),
    .X(net201));
 sg13g2_buf_1 _3161_ (.A(net1065),
    .X(net202));
 sg13g2_buf_1 _3162_ (.A(net1059),
    .X(net203));
 sg13g2_fill_2 FILLER_0_219 ();
 sg13g2_buf_1 _3164_ (.A(\Inst_LUT4AB_switch_matrix.N1BEG1 ),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold22 (.A(\Inst_LB_LUT4c_frame_config_dffesr.LUT_flop ),
    .X(net395));
 sg13g2_fill_2 FILLER_0_44 ();
 sg13g2_buf_2 _3167_ (.A(\Inst_LUT4AB_switch_matrix.JN2BEG0 ),
    .X(net217));
 sg13g2_buf_8 _3168_ (.A(\Inst_LUT4AB_switch_matrix.JN2BEG1 ),
    .X(net218));
 sg13g2_buf_8 _3169_ (.A(\Inst_LUT4AB_switch_matrix.JN2BEG2 ),
    .X(net219));
 sg13g2_buf_1 _3170_ (.A(\Inst_LUT4AB_switch_matrix.JN2BEG3 ),
    .X(net220));
 sg13g2_buf_2 _3171_ (.A(\Inst_LUT4AB_switch_matrix.JN2BEG4 ),
    .X(net221));
 sg13g2_fill_1 FILLER_0_46 ();
 sg13g2_buf_1 _3173_ (.A(\Inst_LUT4AB_switch_matrix.JN2BEG6 ),
    .X(net223));
 sg13g2_buf_1 _3174_ (.A(\Inst_LUT4AB_switch_matrix.JN2BEG7 ),
    .X(net224));
 sg13g2_buf_1 _3175_ (.A(net43),
    .X(net225));
 sg13g2_buf_1 _3176_ (.A(net44),
    .X(net226));
 sg13g2_buf_1 _3177_ (.A(net45),
    .X(net227));
 sg13g2_buf_1 _3178_ (.A(net46),
    .X(net228));
 sg13g2_buf_1 _3179_ (.A(net47),
    .X(net229));
 sg13g2_buf_1 _3180_ (.A(net48),
    .X(net230));
 sg13g2_buf_1 _3181_ (.A(net49),
    .X(net231));
 sg13g2_buf_1 _3182_ (.A(net50),
    .X(net232));
 sg13g2_buf_1 _3183_ (.A(N4END[4]),
    .X(net233));
 sg13g2_buf_1 _3184_ (.A(N4END[5]),
    .X(net240));
 sg13g2_buf_1 _3185_ (.A(N4END[6]),
    .X(net241));
 sg13g2_buf_1 _3186_ (.A(N4END[7]),
    .X(net242));
 sg13g2_buf_1 _3187_ (.A(N4END[8]),
    .X(net243));
 sg13g2_buf_1 _3188_ (.A(N4END[9]),
    .X(net244));
 sg13g2_buf_1 _3189_ (.A(N4END[10]),
    .X(net245));
 sg13g2_buf_1 _3190_ (.A(N4END[11]),
    .X(net246));
 sg13g2_buf_1 _3191_ (.A(N4END[12]),
    .X(net247));
 sg13g2_buf_1 _3192_ (.A(N4END[13]),
    .X(net248));
 sg13g2_buf_1 _3193_ (.A(N4END[14]),
    .X(net234));
 sg13g2_buf_1 _3194_ (.A(N4END[15]),
    .X(net235));
 sg13g2_buf_1 _3195_ (.A(\Inst_LUT4AB_switch_matrix.N4BEG0 ),
    .X(net236));
 sg13g2_buf_1 _3196_ (.A(\Inst_LUT4AB_switch_matrix.N4BEG1 ),
    .X(net237));
 sg13g2_buf_1 _3197_ (.A(\Inst_LUT4AB_switch_matrix.N4BEG2 ),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold18 (.A(\Inst_LD_LUT4c_frame_config_dffesr.LUT_flop ),
    .X(net391));
 sg13g2_buf_1 _3199_ (.A(NN4END[4]),
    .X(net249));
 sg13g2_buf_1 _3200_ (.A(NN4END[5]),
    .X(net256));
 sg13g2_buf_1 _3201_ (.A(NN4END[6]),
    .X(net257));
 sg13g2_buf_1 _3202_ (.A(NN4END[7]),
    .X(net258));
 sg13g2_buf_1 _3203_ (.A(NN4END[8]),
    .X(net259));
 sg13g2_buf_1 _3204_ (.A(NN4END[9]),
    .X(net260));
 sg13g2_buf_1 _3205_ (.A(NN4END[10]),
    .X(net261));
 sg13g2_buf_1 _3206_ (.A(NN4END[11]),
    .X(net262));
 sg13g2_buf_1 _3207_ (.A(NN4END[12]),
    .X(net263));
 sg13g2_buf_1 _3208_ (.A(NN4END[13]),
    .X(net264));
 sg13g2_buf_1 _3209_ (.A(NN4END[14]),
    .X(net250));
 sg13g2_buf_1 _3210_ (.A(NN4END[15]),
    .X(net251));
 sg13g2_buf_1 _3211_ (.A(\Inst_LUT4AB_switch_matrix.NN4BEG0 ),
    .X(net252));
 sg13g2_buf_1 _3212_ (.A(\Inst_LUT4AB_switch_matrix.NN4BEG1 ),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold20 (.A(\Inst_LF_LUT4c_frame_config_dffesr.LUT_flop ),
    .X(net393));
 sg13g2_fill_1 FILLER_0_221 ();
 sg13g2_buf_1 _3215_ (.A(\Inst_LUT4AB_switch_matrix.S1BEG0 ),
    .X(net265));
 sg13g2_buf_1 _3216_ (.A(\Inst_LUT4AB_switch_matrix.S1BEG1 ),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold21 (.A(\Inst_LA_LUT4c_frame_config_dffesr.LUT_flop ),
    .X(net394));
 sg13g2_fill_2 FILLER_0_0 ();
 sg13g2_buf_1 _3219_ (.A(\Inst_LUT4AB_switch_matrix.JS2BEG0 ),
    .X(net269));
 sg13g2_buf_1 _3220_ (.A(\Inst_LUT4AB_switch_matrix.JS2BEG1 ),
    .X(net270));
 sg13g2_buf_1 _3221_ (.A(\Inst_LUT4AB_switch_matrix.JS2BEG2 ),
    .X(net271));
 sg13g2_buf_1 _3222_ (.A(\Inst_LUT4AB_switch_matrix.JS2BEG3 ),
    .X(net272));
 sg13g2_buf_1 _3223_ (.A(\Inst_LUT4AB_switch_matrix.JS2BEG4 ),
    .X(net273));
 sg13g2_fill_1 FILLER_0_157 ();
 sg13g2_buf_1 _3225_ (.A(\Inst_LUT4AB_switch_matrix.JS2BEG6 ),
    .X(net275));
 sg13g2_buf_1 _3226_ (.A(\Inst_LUT4AB_switch_matrix.JS2BEG7 ),
    .X(net276));
 sg13g2_buf_1 _3227_ (.A(net71),
    .X(net277));
 sg13g2_buf_1 _3228_ (.A(net72),
    .X(net278));
 sg13g2_buf_1 _3229_ (.A(net73),
    .X(net279));
 sg13g2_buf_1 _3230_ (.A(net74),
    .X(net280));
 sg13g2_buf_1 _3231_ (.A(net75),
    .X(net281));
 sg13g2_buf_1 _3232_ (.A(net76),
    .X(net282));
 sg13g2_buf_1 _3233_ (.A(net77),
    .X(net283));
 sg13g2_buf_1 _3234_ (.A(net78),
    .X(net284));
 sg13g2_buf_1 _3235_ (.A(S4END[4]),
    .X(net285));
 sg13g2_buf_1 _3236_ (.A(S4END[5]),
    .X(net292));
 sg13g2_buf_1 _3237_ (.A(S4END[6]),
    .X(net293));
 sg13g2_buf_1 _3238_ (.A(S4END[7]),
    .X(net294));
 sg13g2_buf_1 _3239_ (.A(S4END[8]),
    .X(net295));
 sg13g2_buf_1 _3240_ (.A(S4END[9]),
    .X(net296));
 sg13g2_buf_1 _3241_ (.A(S4END[10]),
    .X(net297));
 sg13g2_buf_1 _3242_ (.A(S4END[11]),
    .X(net298));
 sg13g2_buf_1 _3243_ (.A(S4END[12]),
    .X(net299));
 sg13g2_buf_1 _3244_ (.A(S4END[13]),
    .X(net300));
 sg13g2_buf_1 _3245_ (.A(S4END[14]),
    .X(net286));
 sg13g2_buf_1 _3246_ (.A(S4END[15]),
    .X(net287));
 sg13g2_buf_1 _3247_ (.A(\Inst_LUT4AB_switch_matrix.S4BEG0 ),
    .X(net288));
 sg13g2_buf_1 _3248_ (.A(\Inst_LUT4AB_switch_matrix.S4BEG1 ),
    .X(net289));
 sg13g2_buf_1 _3249_ (.A(\Inst_LUT4AB_switch_matrix.S4BEG2 ),
    .X(net290));
 sg13g2_buf_1 _3250_ (.A(\Inst_LUT4AB_switch_matrix.S4BEG3 ),
    .X(net291));
 sg13g2_buf_1 _3251_ (.A(SS4END[4]),
    .X(net301));
 sg13g2_buf_1 _3252_ (.A(SS4END[5]),
    .X(net308));
 sg13g2_buf_1 _3253_ (.A(SS4END[6]),
    .X(net309));
 sg13g2_buf_1 _3254_ (.A(SS4END[7]),
    .X(net310));
 sg13g2_buf_1 _3255_ (.A(SS4END[8]),
    .X(net311));
 sg13g2_buf_1 _3256_ (.A(SS4END[9]),
    .X(net312));
 sg13g2_buf_1 _3257_ (.A(SS4END[10]),
    .X(net313));
 sg13g2_buf_1 _3258_ (.A(SS4END[11]),
    .X(net314));
 sg13g2_buf_1 _3259_ (.A(SS4END[12]),
    .X(net315));
 sg13g2_buf_1 _3260_ (.A(SS4END[13]),
    .X(net316));
 sg13g2_buf_1 _3261_ (.A(SS4END[14]),
    .X(net302));
 sg13g2_buf_1 _3262_ (.A(SS4END[15]),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold17 (.A(\Inst_LG_LUT4c_frame_config_dffesr.LUT_flop ),
    .X(net390));
 sg13g2_buf_1 _3264_ (.A(\Inst_LUT4AB_switch_matrix.SS4BEG1 ),
    .X(net305));
 sg13g2_buf_1 _3265_ (.A(\Inst_LUT4AB_switch_matrix.SS4BEG2 ),
    .X(net306));
 sg13g2_fill_1 FILLER_0_294 ();
 sg13g2_buf_1 _3267_ (.A(UserCLK),
    .X(net317));
 sg13g2_buf_1 _3268_ (.A(\Inst_LUT4AB_switch_matrix.W1BEG0 ),
    .X(net318));
 sg13g2_buf_1 _3269_ (.A(\Inst_LUT4AB_switch_matrix.W1BEG1 ),
    .X(net319));
 sg13g2_buf_1 _3270_ (.A(\Inst_LUT4AB_switch_matrix.W1BEG2 ),
    .X(net320));
 sg13g2_fill_1 FILLER_0_175 ();
 sg13g2_buf_1 _3272_ (.A(\Inst_LUT4AB_switch_matrix.JW2BEG0 ),
    .X(net322));
 sg13g2_buf_1 _3273_ (.A(\Inst_LUT4AB_switch_matrix.JW2BEG1 ),
    .X(net323));
 sg13g2_buf_1 _3274_ (.A(\Inst_LUT4AB_switch_matrix.JW2BEG2 ),
    .X(net324));
 sg13g2_buf_1 _3275_ (.A(\Inst_LUT4AB_switch_matrix.JW2BEG3 ),
    .X(net325));
 sg13g2_buf_1 _3276_ (.A(\Inst_LUT4AB_switch_matrix.JW2BEG4 ),
    .X(net326));
 sg13g2_buf_1 _3277_ (.A(net377),
    .X(net327));
 sg13g2_buf_8 _3278_ (.A(\Inst_LUT4AB_switch_matrix.JW2BEG6 ),
    .X(net328));
 sg13g2_buf_1 _3279_ (.A(\Inst_LUT4AB_switch_matrix.JW2BEG7 ),
    .X(net329));
 sg13g2_buf_1 _3280_ (.A(net98),
    .X(net330));
 sg13g2_buf_1 _3281_ (.A(net99),
    .X(net331));
 sg13g2_buf_1 _3282_ (.A(net100),
    .X(net332));
 sg13g2_buf_1 _3283_ (.A(net101),
    .X(net333));
 sg13g2_buf_1 _3284_ (.A(net102),
    .X(net334));
 sg13g2_buf_1 _3285_ (.A(net103),
    .X(net335));
 sg13g2_buf_1 _3286_ (.A(net104),
    .X(net336));
 sg13g2_buf_1 _3287_ (.A(net105),
    .X(net337));
 sg13g2_buf_1 _3288_ (.A(W6END[2]),
    .X(net338));
 sg13g2_buf_1 _3289_ (.A(W6END[3]),
    .X(net341));
 sg13g2_buf_1 _3290_ (.A(W6END[4]),
    .X(net342));
 sg13g2_buf_1 _3291_ (.A(W6END[5]),
    .X(net343));
 sg13g2_buf_1 _3292_ (.A(W6END[6]),
    .X(net344));
 sg13g2_buf_1 _3293_ (.A(W6END[7]),
    .X(net345));
 sg13g2_buf_1 _3294_ (.A(W6END[8]),
    .X(net346));
 sg13g2_buf_1 _3295_ (.A(W6END[9]),
    .X(net347));
 sg13g2_buf_1 _3296_ (.A(W6END[10]),
    .X(net348));
 sg13g2_buf_1 _3297_ (.A(W6END[11]),
    .X(net349));
 sg13g2_fill_2 FILLER_0_155 ();
 sg13g2_fill_2 FILLER_0_332 ();
 sg13g2_buf_1 _3300_ (.A(WW4END[4]),
    .X(net350));
 sg13g2_buf_1 _3301_ (.A(WW4END[5]),
    .X(net357));
 sg13g2_buf_1 _3302_ (.A(WW4END[6]),
    .X(net358));
 sg13g2_buf_1 _3303_ (.A(WW4END[7]),
    .X(net359));
 sg13g2_buf_1 _3304_ (.A(WW4END[8]),
    .X(net360));
 sg13g2_buf_1 _3305_ (.A(WW4END[9]),
    .X(net361));
 sg13g2_buf_1 _3306_ (.A(WW4END[10]),
    .X(net362));
 sg13g2_buf_1 _3307_ (.A(WW4END[11]),
    .X(net363));
 sg13g2_buf_1 _3308_ (.A(WW4END[12]),
    .X(net364));
 sg13g2_buf_1 _3309_ (.A(WW4END[13]),
    .X(net365));
 sg13g2_buf_1 _3310_ (.A(WW4END[14]),
    .X(net351));
 sg13g2_buf_1 _3311_ (.A(WW4END[15]),
    .X(net352));
 sg13g2_buf_1 _3312_ (.A(\Inst_LUT4AB_switch_matrix.WW4BEG0 ),
    .X(net353));
 sg13g2_buf_1 _3313_ (.A(\Inst_LUT4AB_switch_matrix.WW4BEG1 ),
    .X(net354));
 sg13g2_buf_1 _3314_ (.A(\Inst_LUT4AB_switch_matrix.WW4BEG2 ),
    .X(net355));
 sg13g2_fill_1 FILLER_0_251 ();
 sg13g2_buf_2 fanout925 (.A(_0985_),
    .X(net925));
 sg13g2_buf_1 fanout926 (.A(_0395_),
    .X(net926));
 sg13g2_buf_8 fanout927 (.A(_0973_),
    .X(net927));
 sg13g2_buf_1 fanout928 (.A(\Inst_LUT4AB_switch_matrix.M_AH ),
    .X(net928));
 sg13g2_buf_2 fanout929 (.A(\Inst_LUT4AB_switch_matrix.M_EF ),
    .X(net929));
 sg13g2_buf_4 fanout930 (.X(net930),
    .A(\Inst_LUT4AB_switch_matrix.M_AB ));
 sg13g2_buf_1 fanout931 (.A(\Inst_LUT4AB_switch_matrix.M_AD ),
    .X(net931));
 sg13g2_buf_1 fanout932 (.A(_1052_),
    .X(net932));
 sg13g2_buf_1 fanout933 (.A(_1052_),
    .X(net933));
 sg13g2_buf_16 fanout934 (.X(net934),
    .A(net935));
 sg13g2_buf_8 fanout935 (.A(H),
    .X(net935));
 sg13g2_buf_1 fanout936 (.A(net937),
    .X(net936));
 sg13g2_buf_1 fanout937 (.A(H),
    .X(net937));
 sg13g2_buf_2 fanout938 (.A(net939),
    .X(net938));
 sg13g2_buf_2 fanout939 (.A(net940),
    .X(net939));
 sg13g2_buf_1 fanout940 (.A(C),
    .X(net940));
 sg13g2_buf_1 fanout941 (.A(net942),
    .X(net941));
 sg13g2_buf_16 fanout942 (.X(net942),
    .A(net943));
 sg13g2_buf_8 fanout943 (.A(C),
    .X(net943));
 sg13g2_buf_2 fanout944 (.A(net945),
    .X(net944));
 sg13g2_buf_1 fanout945 (.A(D),
    .X(net945));
 sg13g2_buf_16 fanout946 (.X(net946),
    .A(net947));
 sg13g2_buf_16 fanout947 (.X(net947),
    .A(net948));
 sg13g2_buf_16 fanout948 (.X(net948),
    .A(D));
 sg13g2_dlygate4sd1_1 rebuffer7 (.A(\Inst_LUT4AB_switch_matrix.JS2BEG4 ),
    .X(net380));
 sg13g2_buf_1 fanout950 (.A(net952),
    .X(net950));
 sg13g2_buf_16 fanout951 (.X(net951),
    .A(net952));
 sg13g2_buf_8 fanout952 (.A(G),
    .X(net952));
 sg13g2_buf_1 fanout953 (.A(net954),
    .X(net953));
 sg13g2_buf_1 fanout954 (.A(G),
    .X(net954));
 sg13g2_buf_16 fanout955 (.X(net955),
    .A(net956));
 sg13g2_buf_16 fanout956 (.X(net956),
    .A(net957));
 sg13g2_buf_16 fanout957 (.X(net957),
    .A(F));
 sg13g2_buf_2 fanout958 (.A(net959),
    .X(net958));
 sg13g2_buf_2 fanout959 (.A(net960),
    .X(net959));
 sg13g2_buf_1 fanout960 (.A(F),
    .X(net960));
 sg13g2_buf_1 fanout961 (.A(net963),
    .X(net961));
 sg13g2_buf_16 fanout962 (.X(net962),
    .A(net963));
 sg13g2_buf_16 fanout963 (.X(net963),
    .A(net964));
 sg13g2_buf_8 fanout964 (.A(E),
    .X(net964));
 sg13g2_buf_1 fanout965 (.A(net966),
    .X(net965));
 sg13g2_buf_1 fanout966 (.A(net967),
    .X(net966));
 sg13g2_buf_1 fanout967 (.A(E),
    .X(net967));
 sg13g2_buf_1 fanout968 (.A(net970),
    .X(net968));
 sg13g2_buf_16 fanout969 (.X(net969),
    .A(net970));
 sg13g2_buf_8 fanout970 (.A(B),
    .X(net970));
 sg13g2_buf_1 fanout971 (.A(net972),
    .X(net971));
 sg13g2_buf_1 fanout972 (.A(net973),
    .X(net972));
 sg13g2_buf_1 fanout973 (.A(B),
    .X(net973));
 sg13g2_buf_16 fanout974 (.X(net974),
    .A(net975));
 sg13g2_buf_16 fanout975 (.X(net975),
    .A(A));
 sg13g2_buf_1 fanout976 (.A(net977),
    .X(net976));
 sg13g2_buf_1 fanout977 (.A(net979),
    .X(net977));
 sg13g2_buf_1 fanout978 (.A(net979),
    .X(net978));
 sg13g2_buf_1 fanout979 (.A(A),
    .X(net979));
 sg13g2_buf_1 fanout980 (.A(_0586_),
    .X(net980));
 sg13g2_buf_1 fanout981 (.A(_0586_),
    .X(net981));
 sg13g2_buf_8 fanout982 (.A(_1121_),
    .X(net982));
 sg13g2_buf_1 fanout983 (.A(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit18.Q ),
    .X(net983));
 sg13g2_buf_1 fanout984 (.A(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit10.Q ),
    .X(net984));
 sg13g2_buf_1 fanout985 (.A(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit2.Q ),
    .X(net985));
 sg13g2_buf_1 fanout986 (.A(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit26.Q ),
    .X(net986));
 sg13g2_buf_1 fanout987 (.A(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit14.Q ),
    .X(net987));
 sg13g2_buf_1 fanout988 (.A(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit10.Q ),
    .X(net988));
 sg13g2_buf_1 fanout989 (.A(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit10.Q ),
    .X(net989));
 sg13g2_buf_1 fanout990 (.A(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit2.Q ),
    .X(net990));
 sg13g2_buf_1 fanout991 (.A(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit26.Q ),
    .X(net991));
 sg13g2_buf_1 fanout992 (.A(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit18.Q ),
    .X(net992));
 sg13g2_buf_1 fanout993 (.A(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit2.Q ),
    .X(net993));
 sg13g2_buf_1 fanout994 (.A(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit26.Q ),
    .X(net994));
 sg13g2_buf_1 fanout995 (.A(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit26.Q ),
    .X(net995));
 sg13g2_buf_1 fanout996 (.A(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit18.Q ),
    .X(net996));
 sg13g2_buf_1 fanout997 (.A(net998),
    .X(net997));
 sg13g2_buf_1 fanout998 (.A(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit14.Q ),
    .X(net998));
 sg13g2_buf_1 fanout999 (.A(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit10.Q ),
    .X(net999));
 sg13g2_buf_1 fanout1000 (.A(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit6.Q ),
    .X(net1000));
 sg13g2_buf_1 fanout1001 (.A(net1002),
    .X(net1001));
 sg13g2_buf_1 fanout1002 (.A(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit26.Q ),
    .X(net1002));
 sg13g2_buf_1 fanout1003 (.A(net89),
    .X(net1003));
 sg13g2_buf_1 fanout1004 (.A(net1005),
    .X(net1004));
 sg13g2_buf_1 fanout1005 (.A(W1END[2]),
    .X(net1005));
 sg13g2_buf_1 fanout1006 (.A(net88),
    .X(net1006));
 sg13g2_buf_1 fanout1007 (.A(net34),
    .X(net1007));
 sg13g2_buf_1 fanout1008 (.A(net33),
    .X(net1008));
 sg13g2_buf_1 fanout1009 (.A(net32),
    .X(net1009));
 sg13g2_buf_1 fanout1010 (.A(net31),
    .X(net1010));
 sg13g2_buf_1 fanout1011 (.A(FrameStrobe[9]),
    .X(net1011));
 sg13g2_buf_1 fanout1012 (.A(FrameStrobe[9]),
    .X(net1012));
 sg13g2_buf_1 fanout1013 (.A(net1014),
    .X(net1013));
 sg13g2_buf_1 fanout1014 (.A(net1015),
    .X(net1014));
 sg13g2_buf_1 fanout1015 (.A(FrameStrobe[9]),
    .X(net1015));
 sg13g2_buf_1 fanout1016 (.A(net1020),
    .X(net1016));
 sg13g2_buf_1 fanout1017 (.A(net1018),
    .X(net1017));
 sg13g2_buf_1 fanout1018 (.A(net1020),
    .X(net1018));
 sg13g2_buf_1 fanout1019 (.A(net1020),
    .X(net1019));
 sg13g2_buf_1 fanout1020 (.A(FrameStrobe[8]),
    .X(net1020));
 sg13g2_buf_1 fanout1021 (.A(net1022),
    .X(net1021));
 sg13g2_buf_1 fanout1022 (.A(net30),
    .X(net1022));
 sg13g2_buf_1 fanout1023 (.A(net1024),
    .X(net1023));
 sg13g2_buf_1 fanout1024 (.A(net1025),
    .X(net1024));
 sg13g2_buf_1 fanout1025 (.A(net30),
    .X(net1025));
 sg13g2_buf_1 fanout1026 (.A(net1028),
    .X(net1026));
 sg13g2_buf_1 fanout1027 (.A(net1028),
    .X(net1027));
 sg13g2_buf_1 fanout1028 (.A(FrameStrobe[6]),
    .X(net1028));
 sg13g2_buf_1 fanout1029 (.A(net1030),
    .X(net1029));
 sg13g2_buf_1 fanout1030 (.A(net1031),
    .X(net1030));
 sg13g2_buf_1 fanout1031 (.A(FrameStrobe[6]),
    .X(net1031));
 sg13g2_buf_1 fanout1032 (.A(net1033),
    .X(net1032));
 sg13g2_buf_1 fanout1033 (.A(net1034),
    .X(net1033));
 sg13g2_buf_1 fanout1034 (.A(net29),
    .X(net1034));
 sg13g2_buf_1 fanout1035 (.A(net1036),
    .X(net1035));
 sg13g2_buf_1 fanout1036 (.A(net29),
    .X(net1036));
 sg13g2_buf_1 fanout1037 (.A(FrameStrobe[4]),
    .X(net1037));
 sg13g2_buf_1 fanout1038 (.A(FrameStrobe[4]),
    .X(net1038));
 sg13g2_buf_1 fanout1039 (.A(net1040),
    .X(net1039));
 sg13g2_buf_1 fanout1040 (.A(net1041),
    .X(net1040));
 sg13g2_buf_1 fanout1041 (.A(FrameStrobe[4]),
    .X(net1041));
 sg13g2_buf_1 fanout1042 (.A(net1043),
    .X(net1042));
 sg13g2_buf_1 fanout1043 (.A(net1046),
    .X(net1043));
 sg13g2_buf_1 fanout1044 (.A(net1046),
    .X(net1044));
 sg13g2_buf_1 fanout1045 (.A(net1046),
    .X(net1045));
 sg13g2_buf_1 fanout1046 (.A(FrameStrobe[3]),
    .X(net1046));
 sg13g2_buf_1 fanout1047 (.A(net1049),
    .X(net1047));
 sg13g2_buf_1 fanout1048 (.A(net1049),
    .X(net1048));
 sg13g2_buf_1 fanout1049 (.A(FrameStrobe[2]),
    .X(net1049));
 sg13g2_buf_1 fanout1050 (.A(net1052),
    .X(net1050));
 sg13g2_buf_1 fanout1051 (.A(net1052),
    .X(net1051));
 sg13g2_buf_1 fanout1052 (.A(FrameStrobe[2]),
    .X(net1052));
 sg13g2_buf_1 fanout1053 (.A(net1054),
    .X(net1053));
 sg13g2_buf_1 fanout1054 (.A(net1055),
    .X(net1054));
 sg13g2_buf_1 fanout1055 (.A(net1058),
    .X(net1055));
 sg13g2_buf_1 fanout1056 (.A(net1058),
    .X(net1056));
 sg13g2_buf_1 fanout1057 (.A(net1058),
    .X(net1057));
 sg13g2_buf_1 fanout1058 (.A(FrameStrobe[1]),
    .X(net1058));
 sg13g2_buf_1 fanout1059 (.A(net28),
    .X(net1059));
 sg13g2_buf_1 fanout1060 (.A(net1062),
    .X(net1060));
 sg13g2_buf_1 fanout1061 (.A(net1062),
    .X(net1061));
 sg13g2_buf_1 fanout1062 (.A(FrameStrobe[18]),
    .X(net1062));
 sg13g2_buf_1 fanout1063 (.A(net1064),
    .X(net1063));
 sg13g2_buf_1 fanout1064 (.A(net1065),
    .X(net1064));
 sg13g2_buf_1 fanout1065 (.A(FrameStrobe[18]),
    .X(net1065));
 sg13g2_buf_1 fanout1066 (.A(net1067),
    .X(net1066));
 sg13g2_buf_1 fanout1067 (.A(net1068),
    .X(net1067));
 sg13g2_buf_1 fanout1068 (.A(FrameStrobe[17]),
    .X(net1068));
 sg13g2_buf_1 fanout1069 (.A(net1070),
    .X(net1069));
 sg13g2_buf_1 fanout1070 (.A(FrameStrobe[17]),
    .X(net1070));
 sg13g2_buf_1 fanout1071 (.A(net1073),
    .X(net1071));
 sg13g2_buf_1 fanout1072 (.A(net1073),
    .X(net1072));
 sg13g2_buf_1 fanout1073 (.A(net1074),
    .X(net1073));
 sg13g2_buf_1 fanout1074 (.A(net1076),
    .X(net1074));
 sg13g2_buf_1 fanout1075 (.A(net1076),
    .X(net1075));
 sg13g2_buf_1 fanout1076 (.A(FrameStrobe[16]),
    .X(net1076));
 sg13g2_buf_1 fanout1077 (.A(net1078),
    .X(net1077));
 sg13g2_buf_1 fanout1078 (.A(net1079),
    .X(net1078));
 sg13g2_buf_1 fanout1079 (.A(FrameStrobe[15]),
    .X(net1079));
 sg13g2_buf_1 fanout1080 (.A(net1081),
    .X(net1080));
 sg13g2_buf_1 fanout1081 (.A(FrameStrobe[15]),
    .X(net1081));
 sg13g2_buf_1 fanout1082 (.A(net1086),
    .X(net1082));
 sg13g2_buf_1 fanout1083 (.A(net1085),
    .X(net1083));
 sg13g2_buf_1 fanout1084 (.A(net1085),
    .X(net1084));
 sg13g2_buf_1 fanout1085 (.A(net1086),
    .X(net1085));
 sg13g2_buf_1 fanout1086 (.A(FrameStrobe[14]),
    .X(net1086));
 sg13g2_buf_1 fanout1087 (.A(net1092),
    .X(net1087));
 sg13g2_buf_1 fanout1088 (.A(net1089),
    .X(net1088));
 sg13g2_buf_1 fanout1089 (.A(net1091),
    .X(net1089));
 sg13g2_buf_1 fanout1090 (.A(net1091),
    .X(net1090));
 sg13g2_buf_1 fanout1091 (.A(net1092),
    .X(net1091));
 sg13g2_buf_1 fanout1092 (.A(FrameStrobe[13]),
    .X(net1092));
 sg13g2_buf_1 fanout1093 (.A(net1094),
    .X(net1093));
 sg13g2_buf_1 fanout1094 (.A(net1095),
    .X(net1094));
 sg13g2_buf_1 fanout1095 (.A(FrameStrobe[12]),
    .X(net1095));
 sg13g2_buf_1 fanout1096 (.A(net1097),
    .X(net1096));
 sg13g2_buf_1 fanout1097 (.A(FrameStrobe[12]),
    .X(net1097));
 sg13g2_buf_1 fanout1098 (.A(net1099),
    .X(net1098));
 sg13g2_buf_1 fanout1099 (.A(net1100),
    .X(net1099));
 sg13g2_buf_1 fanout1100 (.A(net1101),
    .X(net1100));
 sg13g2_buf_1 fanout1101 (.A(net1102),
    .X(net1101));
 sg13g2_buf_1 fanout1102 (.A(net27),
    .X(net1102));
 sg13g2_buf_1 fanout1103 (.A(net1104),
    .X(net1103));
 sg13g2_buf_1 fanout1104 (.A(net1105),
    .X(net1104));
 sg13g2_buf_1 fanout1105 (.A(net1108),
    .X(net1105));
 sg13g2_buf_1 fanout1106 (.A(net1107),
    .X(net1106));
 sg13g2_buf_1 fanout1107 (.A(net1108),
    .X(net1107));
 sg13g2_buf_1 fanout1108 (.A(FrameStrobe[10]),
    .X(net1108));
 sg13g2_buf_1 fanout1109 (.A(net1112),
    .X(net1109));
 sg13g2_buf_1 fanout1110 (.A(net1112),
    .X(net1110));
 sg13g2_buf_1 fanout1111 (.A(net1112),
    .X(net1111));
 sg13g2_buf_1 fanout1112 (.A(FrameStrobe[0]),
    .X(net1112));
 sg13g2_buf_1 fanout1113 (.A(FrameStrobe[0]),
    .X(net1113));
 sg13g2_buf_1 fanout1114 (.A(FrameData[9]),
    .X(net1114));
 sg13g2_buf_1 fanout1115 (.A(FrameData[9]),
    .X(net1115));
 sg13g2_buf_1 fanout1116 (.A(FrameData[9]),
    .X(net1116));
 sg13g2_buf_1 fanout1117 (.A(FrameData[8]),
    .X(net1117));
 sg13g2_buf_1 fanout1118 (.A(FrameData[8]),
    .X(net1118));
 sg13g2_buf_1 fanout1119 (.A(FrameData[8]),
    .X(net1119));
 sg13g2_buf_1 fanout1120 (.A(net1122),
    .X(net1120));
 sg13g2_buf_1 fanout1121 (.A(net1122),
    .X(net1121));
 sg13g2_buf_1 fanout1122 (.A(FrameData[7]),
    .X(net1122));
 sg13g2_buf_1 fanout1123 (.A(net1125),
    .X(net1123));
 sg13g2_buf_1 fanout1124 (.A(net1125),
    .X(net1124));
 sg13g2_buf_1 fanout1125 (.A(FrameData[6]),
    .X(net1125));
 sg13g2_buf_1 fanout1126 (.A(net1128),
    .X(net1126));
 sg13g2_buf_1 fanout1127 (.A(net1128),
    .X(net1127));
 sg13g2_buf_1 fanout1128 (.A(FrameData[5]),
    .X(net1128));
 sg13g2_buf_1 fanout1129 (.A(FrameData[4]),
    .X(net1129));
 sg13g2_buf_1 fanout1130 (.A(FrameData[4]),
    .X(net1130));
 sg13g2_buf_1 fanout1131 (.A(FrameData[4]),
    .X(net1131));
 sg13g2_buf_1 fanout1132 (.A(FrameData[3]),
    .X(net1132));
 sg13g2_buf_1 fanout1133 (.A(FrameData[3]),
    .X(net1133));
 sg13g2_buf_1 fanout1134 (.A(FrameData[3]),
    .X(net1134));
 sg13g2_buf_1 fanout1135 (.A(net1136),
    .X(net1135));
 sg13g2_buf_1 fanout1136 (.A(net1137),
    .X(net1136));
 sg13g2_buf_1 fanout1137 (.A(FrameData[31]),
    .X(net1137));
 sg13g2_buf_1 fanout1138 (.A(net1139),
    .X(net1138));
 sg13g2_buf_1 fanout1139 (.A(net1140),
    .X(net1139));
 sg13g2_buf_1 fanout1140 (.A(FrameData[30]),
    .X(net1140));
 sg13g2_buf_1 fanout1141 (.A(FrameData[2]),
    .X(net1141));
 sg13g2_buf_1 fanout1142 (.A(FrameData[2]),
    .X(net1142));
 sg13g2_buf_1 fanout1143 (.A(FrameData[2]),
    .X(net1143));
 sg13g2_buf_1 fanout1144 (.A(FrameData[29]),
    .X(net1144));
 sg13g2_buf_1 fanout1145 (.A(FrameData[29]),
    .X(net1145));
 sg13g2_buf_1 fanout1146 (.A(FrameData[29]),
    .X(net1146));
 sg13g2_buf_1 fanout1147 (.A(net1148),
    .X(net1147));
 sg13g2_buf_1 fanout1148 (.A(net1149),
    .X(net1148));
 sg13g2_buf_1 fanout1149 (.A(FrameData[28]),
    .X(net1149));
 sg13g2_buf_1 fanout1150 (.A(net1151),
    .X(net1150));
 sg13g2_buf_1 fanout1151 (.A(FrameData[27]),
    .X(net1151));
 sg13g2_buf_1 fanout1152 (.A(FrameData[27]),
    .X(net1152));
 sg13g2_buf_1 fanout1153 (.A(FrameData[26]),
    .X(net1153));
 sg13g2_buf_1 fanout1154 (.A(net1155),
    .X(net1154));
 sg13g2_buf_1 fanout1155 (.A(FrameData[26]),
    .X(net1155));
 sg13g2_buf_1 fanout1156 (.A(net1158),
    .X(net1156));
 sg13g2_buf_1 fanout1157 (.A(net1158),
    .X(net1157));
 sg13g2_buf_1 fanout1158 (.A(FrameData[25]),
    .X(net1158));
 sg13g2_buf_1 fanout1159 (.A(net1161),
    .X(net1159));
 sg13g2_buf_1 fanout1160 (.A(net1161),
    .X(net1160));
 sg13g2_buf_1 fanout1161 (.A(FrameData[24]),
    .X(net1161));
 sg13g2_buf_1 fanout1162 (.A(net1164),
    .X(net1162));
 sg13g2_buf_1 fanout1163 (.A(net1164),
    .X(net1163));
 sg13g2_buf_1 fanout1164 (.A(FrameData[23]),
    .X(net1164));
 sg13g2_buf_1 fanout1165 (.A(net1167),
    .X(net1165));
 sg13g2_buf_1 fanout1166 (.A(net1167),
    .X(net1166));
 sg13g2_buf_1 fanout1167 (.A(FrameData[22]),
    .X(net1167));
 sg13g2_buf_1 fanout1168 (.A(net1170),
    .X(net1168));
 sg13g2_buf_1 fanout1169 (.A(net1170),
    .X(net1169));
 sg13g2_buf_1 fanout1170 (.A(FrameData[21]),
    .X(net1170));
 sg13g2_buf_1 fanout1171 (.A(net1173),
    .X(net1171));
 sg13g2_buf_1 fanout1172 (.A(net1173),
    .X(net1172));
 sg13g2_buf_1 fanout1173 (.A(FrameData[20]),
    .X(net1173));
 sg13g2_buf_1 fanout1174 (.A(net1176),
    .X(net1174));
 sg13g2_buf_1 fanout1175 (.A(net1176),
    .X(net1175));
 sg13g2_buf_1 fanout1176 (.A(net26),
    .X(net1176));
 sg13g2_buf_1 fanout1177 (.A(net1179),
    .X(net1177));
 sg13g2_buf_1 fanout1178 (.A(net1179),
    .X(net1178));
 sg13g2_buf_1 fanout1179 (.A(FrameData[19]),
    .X(net1179));
 sg13g2_buf_1 fanout1180 (.A(net1182),
    .X(net1180));
 sg13g2_buf_1 fanout1181 (.A(net1182),
    .X(net1181));
 sg13g2_buf_1 fanout1182 (.A(FrameData[18]),
    .X(net1182));
 sg13g2_buf_1 fanout1183 (.A(net1185),
    .X(net1183));
 sg13g2_buf_1 fanout1184 (.A(net1185),
    .X(net1184));
 sg13g2_buf_1 fanout1185 (.A(FrameData[17]),
    .X(net1185));
 sg13g2_buf_1 fanout1186 (.A(net1188),
    .X(net1186));
 sg13g2_buf_1 fanout1187 (.A(net1188),
    .X(net1187));
 sg13g2_buf_1 fanout1188 (.A(FrameData[16]),
    .X(net1188));
 sg13g2_buf_1 fanout1189 (.A(net1191),
    .X(net1189));
 sg13g2_buf_1 fanout1190 (.A(net1191),
    .X(net1190));
 sg13g2_buf_1 fanout1191 (.A(FrameData[15]),
    .X(net1191));
 sg13g2_buf_1 fanout1192 (.A(net1194),
    .X(net1192));
 sg13g2_buf_1 fanout1193 (.A(net1194),
    .X(net1193));
 sg13g2_buf_1 fanout1194 (.A(FrameData[14]),
    .X(net1194));
 sg13g2_buf_1 fanout1195 (.A(net1197),
    .X(net1195));
 sg13g2_buf_1 fanout1196 (.A(net1197),
    .X(net1196));
 sg13g2_buf_1 fanout1197 (.A(FrameData[13]),
    .X(net1197));
 sg13g2_buf_1 fanout1198 (.A(net1200),
    .X(net1198));
 sg13g2_buf_1 fanout1199 (.A(net1200),
    .X(net1199));
 sg13g2_buf_1 fanout1200 (.A(FrameData[12]),
    .X(net1200));
 sg13g2_buf_1 fanout1201 (.A(net1203),
    .X(net1201));
 sg13g2_buf_1 fanout1202 (.A(net1203),
    .X(net1202));
 sg13g2_buf_1 fanout1203 (.A(FrameData[11]),
    .X(net1203));
 sg13g2_buf_1 fanout1204 (.A(FrameData[10]),
    .X(net1204));
 sg13g2_buf_1 fanout1205 (.A(FrameData[10]),
    .X(net1205));
 sg13g2_buf_1 fanout1206 (.A(FrameData[10]),
    .X(net1206));
 sg13g2_buf_1 fanout1207 (.A(net1209),
    .X(net1207));
 sg13g2_buf_1 fanout1208 (.A(net1209),
    .X(net1208));
 sg13g2_buf_1 fanout1209 (.A(FrameData[0]),
    .X(net1209));
 sg13g2_buf_1 fanout1210 (.A(net1211),
    .X(net1210));
 sg13g2_buf_1 fanout1211 (.A(E6END[1]),
    .X(net1211));
 sg13g2_buf_1 fanout1212 (.A(net1213),
    .X(net1212));
 sg13g2_buf_1 fanout1213 (.A(E6END[0]),
    .X(net1213));
 sg13g2_buf_1 fanout1214 (.A(net5),
    .X(net1214));
 sg13g2_buf_1 fanout1215 (.A(net4),
    .X(net1215));
 sg13g2_buf_1 fanout1216 (.A(net3),
    .X(net1216));
 sg13g2_buf_1 fanout1217 (.A(net2),
    .X(net1217));
 sg13g2_buf_2 input1 (.A(Ci),
    .X(net1));
 sg13g2_buf_1 input2 (.A(E1END[0]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(E1END[1]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(E1END[2]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(E1END[3]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(E2END[0]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(E2END[1]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(E2END[2]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(E2END[3]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(E2END[4]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(E2END[5]),
    .X(net11));
 sg13g2_buf_1 input12 (.A(E2END[6]),
    .X(net12));
 sg13g2_buf_1 input13 (.A(E2END[7]),
    .X(net13));
 sg13g2_buf_1 input14 (.A(E2MID[0]),
    .X(net14));
 sg13g2_buf_16 input15 (.X(net15),
    .A(E2MID[1]));
 sg13g2_buf_1 input16 (.A(E2MID[2]),
    .X(net16));
 sg13g2_buf_1 input17 (.A(E2MID[3]),
    .X(net17));
 sg13g2_buf_1 input18 (.A(E2MID[4]),
    .X(net18));
 sg13g2_buf_1 input19 (.A(E2MID[5]),
    .X(net19));
 sg13g2_buf_1 input20 (.A(E2MID[6]),
    .X(net20));
 sg13g2_buf_1 input21 (.A(E2MID[7]),
    .X(net21));
 sg13g2_buf_1 input22 (.A(EE4END[0]),
    .X(net22));
 sg13g2_buf_1 input23 (.A(EE4END[1]),
    .X(net23));
 sg13g2_buf_1 input24 (.A(EE4END[2]),
    .X(net24));
 sg13g2_buf_1 input25 (.A(EE4END[3]),
    .X(net25));
 sg13g2_buf_1 input26 (.A(FrameData[1]),
    .X(net26));
 sg13g2_buf_1 input27 (.A(FrameStrobe[11]),
    .X(net27));
 sg13g2_buf_1 input28 (.A(FrameStrobe[19]),
    .X(net28));
 sg13g2_buf_1 input29 (.A(FrameStrobe[5]),
    .X(net29));
 sg13g2_buf_1 input30 (.A(FrameStrobe[7]),
    .X(net30));
 sg13g2_buf_1 input31 (.A(N1END[0]),
    .X(net31));
 sg13g2_buf_1 input32 (.A(N1END[1]),
    .X(net32));
 sg13g2_buf_1 input33 (.A(N1END[2]),
    .X(net33));
 sg13g2_buf_1 input34 (.A(N1END[3]),
    .X(net34));
 sg13g2_buf_1 input35 (.A(N2END[0]),
    .X(net35));
 sg13g2_buf_1 input36 (.A(N2END[1]),
    .X(net36));
 sg13g2_buf_1 input37 (.A(N2END[2]),
    .X(net37));
 sg13g2_buf_1 input38 (.A(N2END[3]),
    .X(net38));
 sg13g2_buf_1 input39 (.A(N2END[4]),
    .X(net39));
 sg13g2_buf_1 input40 (.A(N2END[5]),
    .X(net40));
 sg13g2_buf_1 input41 (.A(N2END[6]),
    .X(net41));
 sg13g2_buf_1 input42 (.A(N2END[7]),
    .X(net42));
 sg13g2_buf_1 input43 (.A(N2MID[0]),
    .X(net43));
 sg13g2_buf_8 input44 (.A(N2MID[1]),
    .X(net44));
 sg13g2_buf_1 input45 (.A(N2MID[2]),
    .X(net45));
 sg13g2_buf_1 input46 (.A(N2MID[3]),
    .X(net46));
 sg13g2_buf_1 input47 (.A(N2MID[4]),
    .X(net47));
 sg13g2_buf_1 input48 (.A(N2MID[5]),
    .X(net48));
 sg13g2_buf_1 input49 (.A(N2MID[6]),
    .X(net49));
 sg13g2_buf_1 input50 (.A(N2MID[7]),
    .X(net50));
 sg13g2_buf_1 input51 (.A(N4END[0]),
    .X(net51));
 sg13g2_buf_1 input52 (.A(N4END[1]),
    .X(net52));
 sg13g2_buf_1 input53 (.A(N4END[2]),
    .X(net53));
 sg13g2_buf_1 input54 (.A(N4END[3]),
    .X(net54));
 sg13g2_buf_1 input55 (.A(NN4END[0]),
    .X(net55));
 sg13g2_buf_1 input56 (.A(NN4END[1]),
    .X(net56));
 sg13g2_buf_1 input57 (.A(NN4END[2]),
    .X(net57));
 sg13g2_buf_1 input58 (.A(NN4END[3]),
    .X(net58));
 sg13g2_buf_1 input59 (.A(S1END[0]),
    .X(net59));
 sg13g2_buf_1 input60 (.A(S1END[1]),
    .X(net60));
 sg13g2_buf_1 input61 (.A(S1END[2]),
    .X(net61));
 sg13g2_buf_1 input62 (.A(S1END[3]),
    .X(net62));
 sg13g2_buf_1 input63 (.A(S2END[0]),
    .X(net63));
 sg13g2_buf_1 input64 (.A(S2END[1]),
    .X(net64));
 sg13g2_buf_1 input65 (.A(S2END[2]),
    .X(net65));
 sg13g2_buf_1 input66 (.A(S2END[3]),
    .X(net66));
 sg13g2_buf_1 input67 (.A(S2END[4]),
    .X(net67));
 sg13g2_buf_1 input68 (.A(S2END[5]),
    .X(net68));
 sg13g2_buf_1 input69 (.A(S2END[6]),
    .X(net69));
 sg13g2_buf_1 input70 (.A(S2END[7]),
    .X(net70));
 sg13g2_buf_1 input71 (.A(S2MID[0]),
    .X(net71));
 sg13g2_buf_2 input72 (.A(S2MID[1]),
    .X(net72));
 sg13g2_buf_1 input73 (.A(S2MID[2]),
    .X(net73));
 sg13g2_buf_1 input74 (.A(S2MID[3]),
    .X(net74));
 sg13g2_buf_1 input75 (.A(S2MID[4]),
    .X(net75));
 sg13g2_buf_1 input76 (.A(S2MID[5]),
    .X(net76));
 sg13g2_buf_1 input77 (.A(S2MID[6]),
    .X(net77));
 sg13g2_buf_1 input78 (.A(S2MID[7]),
    .X(net78));
 sg13g2_buf_1 input79 (.A(S4END[0]),
    .X(net79));
 sg13g2_buf_1 input80 (.A(S4END[1]),
    .X(net80));
 sg13g2_buf_1 input81 (.A(S4END[2]),
    .X(net81));
 sg13g2_buf_1 input82 (.A(S4END[3]),
    .X(net82));
 sg13g2_buf_1 input83 (.A(SS4END[0]),
    .X(net83));
 sg13g2_buf_1 input84 (.A(SS4END[1]),
    .X(net84));
 sg13g2_buf_1 input85 (.A(SS4END[2]),
    .X(net85));
 sg13g2_buf_1 input86 (.A(SS4END[3]),
    .X(net86));
 sg13g2_buf_1 input87 (.A(W1END[0]),
    .X(net87));
 sg13g2_buf_1 input88 (.A(W1END[1]),
    .X(net88));
 sg13g2_buf_1 input89 (.A(W1END[3]),
    .X(net89));
 sg13g2_buf_1 input90 (.A(W2END[0]),
    .X(net90));
 sg13g2_buf_1 input91 (.A(W2END[1]),
    .X(net91));
 sg13g2_buf_1 input92 (.A(W2END[2]),
    .X(net92));
 sg13g2_buf_1 input93 (.A(W2END[3]),
    .X(net93));
 sg13g2_buf_1 input94 (.A(W2END[4]),
    .X(net94));
 sg13g2_buf_1 input95 (.A(W2END[5]),
    .X(net95));
 sg13g2_buf_1 input96 (.A(W2END[6]),
    .X(net96));
 sg13g2_buf_1 input97 (.A(W2END[7]),
    .X(net97));
 sg13g2_buf_1 input98 (.A(W2MID[0]),
    .X(net98));
 sg13g2_buf_1 input99 (.A(W2MID[1]),
    .X(net99));
 sg13g2_buf_1 input100 (.A(W2MID[2]),
    .X(net100));
 sg13g2_buf_1 input101 (.A(W2MID[3]),
    .X(net101));
 sg13g2_buf_1 input102 (.A(W2MID[4]),
    .X(net102));
 sg13g2_buf_1 input103 (.A(W2MID[5]),
    .X(net103));
 sg13g2_buf_1 input104 (.A(W2MID[6]),
    .X(net104));
 sg13g2_buf_1 input105 (.A(W2MID[7]),
    .X(net105));
 sg13g2_buf_1 input106 (.A(W6END[0]),
    .X(net106));
 sg13g2_buf_1 input107 (.A(W6END[1]),
    .X(net107));
 sg13g2_buf_1 input108 (.A(WW4END[0]),
    .X(net108));
 sg13g2_buf_1 input109 (.A(WW4END[1]),
    .X(net109));
 sg13g2_buf_1 input110 (.A(WW4END[2]),
    .X(net110));
 sg13g2_buf_1 input111 (.A(WW4END[3]),
    .X(net111));
 sg13g2_buf_1 output112 (.A(net112),
    .X(Co));
 sg13g2_buf_1 output113 (.A(net113),
    .X(E1BEG[0]));
 sg13g2_buf_1 output114 (.A(net114),
    .X(E1BEG[1]));
 sg13g2_buf_1 output115 (.A(\Inst_LUT4AB_switch_matrix.E1BEG2 ),
    .X(E1BEG[2]));
 sg13g2_buf_1 output116 (.A(\Inst_LUT4AB_switch_matrix.E1BEG3 ),
    .X(E1BEG[3]));
 sg13g2_buf_1 output117 (.A(net117),
    .X(E2BEG[0]));
 sg13g2_buf_1 output118 (.A(net118),
    .X(E2BEG[1]));
 sg13g2_buf_1 output119 (.A(net119),
    .X(E2BEG[2]));
 sg13g2_buf_1 output120 (.A(net120),
    .X(E2BEG[3]));
 sg13g2_buf_1 output121 (.A(net121),
    .X(E2BEG[4]));
 sg13g2_buf_1 output122 (.A(\Inst_LUT4AB_switch_matrix.E2BEG5 ),
    .X(E2BEG[5]));
 sg13g2_buf_1 output123 (.A(net123),
    .X(E2BEG[6]));
 sg13g2_buf_1 output124 (.A(\Inst_LUT4AB_switch_matrix.E2BEG7 ),
    .X(E2BEG[7]));
 sg13g2_buf_1 output125 (.A(net125),
    .X(E2BEGb[0]));
 sg13g2_buf_1 output126 (.A(net126),
    .X(E2BEGb[1]));
 sg13g2_buf_1 output127 (.A(net127),
    .X(E2BEGb[2]));
 sg13g2_buf_1 output128 (.A(net128),
    .X(E2BEGb[3]));
 sg13g2_buf_1 output129 (.A(net129),
    .X(E2BEGb[4]));
 sg13g2_buf_1 output130 (.A(net130),
    .X(E2BEGb[5]));
 sg13g2_buf_1 output131 (.A(net131),
    .X(E2BEGb[6]));
 sg13g2_buf_1 output132 (.A(net132),
    .X(E2BEGb[7]));
 sg13g2_buf_1 output133 (.A(net133),
    .X(E6BEG[0]));
 sg13g2_buf_1 output134 (.A(net134),
    .X(E6BEG[10]));
 sg13g2_buf_1 output135 (.A(\Inst_LUT4AB_switch_matrix.E6BEG1 ),
    .X(E6BEG[11]));
 sg13g2_buf_1 output136 (.A(net136),
    .X(E6BEG[1]));
 sg13g2_buf_1 output137 (.A(net137),
    .X(E6BEG[2]));
 sg13g2_buf_1 output138 (.A(net138),
    .X(E6BEG[3]));
 sg13g2_buf_1 output139 (.A(net139),
    .X(E6BEG[4]));
 sg13g2_buf_1 output140 (.A(net140),
    .X(E6BEG[5]));
 sg13g2_buf_1 output141 (.A(net141),
    .X(E6BEG[6]));
 sg13g2_buf_1 output142 (.A(net142),
    .X(E6BEG[7]));
 sg13g2_buf_1 output143 (.A(net143),
    .X(E6BEG[8]));
 sg13g2_buf_1 output144 (.A(net144),
    .X(E6BEG[9]));
 sg13g2_buf_1 output145 (.A(net145),
    .X(EE4BEG[0]));
 sg13g2_buf_1 output146 (.A(net146),
    .X(EE4BEG[10]));
 sg13g2_buf_1 output147 (.A(net147),
    .X(EE4BEG[11]));
 sg13g2_buf_1 output148 (.A(net148),
    .X(EE4BEG[12]));
 sg13g2_buf_1 output149 (.A(net149),
    .X(EE4BEG[13]));
 sg13g2_buf_1 output150 (.A(\Inst_LUT4AB_switch_matrix.EE4BEG2 ),
    .X(EE4BEG[14]));
 sg13g2_buf_1 output151 (.A(\Inst_LUT4AB_switch_matrix.EE4BEG3 ),
    .X(EE4BEG[15]));
 sg13g2_buf_1 output152 (.A(net152),
    .X(EE4BEG[1]));
 sg13g2_buf_1 output153 (.A(net153),
    .X(EE4BEG[2]));
 sg13g2_buf_1 output154 (.A(net154),
    .X(EE4BEG[3]));
 sg13g2_buf_1 output155 (.A(net155),
    .X(EE4BEG[4]));
 sg13g2_buf_1 output156 (.A(net156),
    .X(EE4BEG[5]));
 sg13g2_buf_1 output157 (.A(net157),
    .X(EE4BEG[6]));
 sg13g2_buf_1 output158 (.A(net158),
    .X(EE4BEG[7]));
 sg13g2_buf_1 output159 (.A(net159),
    .X(EE4BEG[8]));
 sg13g2_buf_1 output160 (.A(net160),
    .X(EE4BEG[9]));
 sg13g2_buf_1 output161 (.A(net161),
    .X(FrameData_O[0]));
 sg13g2_buf_1 output162 (.A(net162),
    .X(FrameData_O[10]));
 sg13g2_buf_1 output163 (.A(net163),
    .X(FrameData_O[11]));
 sg13g2_buf_1 output164 (.A(net164),
    .X(FrameData_O[12]));
 sg13g2_buf_1 output165 (.A(net165),
    .X(FrameData_O[13]));
 sg13g2_buf_1 output166 (.A(net166),
    .X(FrameData_O[14]));
 sg13g2_buf_1 output167 (.A(net167),
    .X(FrameData_O[15]));
 sg13g2_buf_1 output168 (.A(net168),
    .X(FrameData_O[16]));
 sg13g2_buf_1 output169 (.A(net169),
    .X(FrameData_O[17]));
 sg13g2_buf_1 output170 (.A(net170),
    .X(FrameData_O[18]));
 sg13g2_buf_1 output171 (.A(net171),
    .X(FrameData_O[19]));
 sg13g2_buf_1 output172 (.A(net172),
    .X(FrameData_O[1]));
 sg13g2_buf_1 output173 (.A(net173),
    .X(FrameData_O[20]));
 sg13g2_buf_1 output174 (.A(net174),
    .X(FrameData_O[21]));
 sg13g2_buf_1 output175 (.A(net175),
    .X(FrameData_O[22]));
 sg13g2_buf_1 output176 (.A(net176),
    .X(FrameData_O[23]));
 sg13g2_buf_1 output177 (.A(net177),
    .X(FrameData_O[24]));
 sg13g2_buf_1 output178 (.A(net178),
    .X(FrameData_O[25]));
 sg13g2_buf_1 output179 (.A(net179),
    .X(FrameData_O[26]));
 sg13g2_buf_1 output180 (.A(net180),
    .X(FrameData_O[27]));
 sg13g2_buf_1 output181 (.A(net181),
    .X(FrameData_O[28]));
 sg13g2_buf_1 output182 (.A(net182),
    .X(FrameData_O[29]));
 sg13g2_buf_1 output183 (.A(net183),
    .X(FrameData_O[2]));
 sg13g2_buf_1 output184 (.A(net184),
    .X(FrameData_O[30]));
 sg13g2_buf_1 output185 (.A(net185),
    .X(FrameData_O[31]));
 sg13g2_buf_1 output186 (.A(net186),
    .X(FrameData_O[3]));
 sg13g2_buf_1 output187 (.A(net187),
    .X(FrameData_O[4]));
 sg13g2_buf_1 output188 (.A(net188),
    .X(FrameData_O[5]));
 sg13g2_buf_1 output189 (.A(net189),
    .X(FrameData_O[6]));
 sg13g2_buf_1 output190 (.A(net190),
    .X(FrameData_O[7]));
 sg13g2_buf_1 output191 (.A(net191),
    .X(FrameData_O[8]));
 sg13g2_buf_1 output192 (.A(net192),
    .X(FrameData_O[9]));
 sg13g2_buf_1 output193 (.A(net193),
    .X(FrameStrobe_O[0]));
 sg13g2_buf_1 output194 (.A(net194),
    .X(FrameStrobe_O[10]));
 sg13g2_buf_1 output195 (.A(net195),
    .X(FrameStrobe_O[11]));
 sg13g2_buf_1 output196 (.A(net196),
    .X(FrameStrobe_O[12]));
 sg13g2_buf_1 output197 (.A(net197),
    .X(FrameStrobe_O[13]));
 sg13g2_buf_1 output198 (.A(net198),
    .X(FrameStrobe_O[14]));
 sg13g2_buf_1 output199 (.A(net199),
    .X(FrameStrobe_O[15]));
 sg13g2_buf_1 output200 (.A(net200),
    .X(FrameStrobe_O[16]));
 sg13g2_buf_1 output201 (.A(net201),
    .X(FrameStrobe_O[17]));
 sg13g2_buf_1 output202 (.A(net202),
    .X(FrameStrobe_O[18]));
 sg13g2_buf_1 output203 (.A(net203),
    .X(FrameStrobe_O[19]));
 sg13g2_buf_1 output204 (.A(net204),
    .X(FrameStrobe_O[1]));
 sg13g2_buf_1 output205 (.A(net205),
    .X(FrameStrobe_O[2]));
 sg13g2_buf_1 output206 (.A(net206),
    .X(FrameStrobe_O[3]));
 sg13g2_buf_1 output207 (.A(net207),
    .X(FrameStrobe_O[4]));
 sg13g2_buf_1 output208 (.A(net208),
    .X(FrameStrobe_O[5]));
 sg13g2_buf_1 output209 (.A(net209),
    .X(FrameStrobe_O[6]));
 sg13g2_buf_1 output210 (.A(net210),
    .X(FrameStrobe_O[7]));
 sg13g2_buf_1 output211 (.A(net211),
    .X(FrameStrobe_O[8]));
 sg13g2_buf_1 output212 (.A(net212),
    .X(FrameStrobe_O[9]));
 sg13g2_buf_1 output213 (.A(\Inst_LUT4AB_switch_matrix.N1BEG0 ),
    .X(N1BEG[0]));
 sg13g2_buf_1 output214 (.A(net214),
    .X(N1BEG[1]));
 sg13g2_buf_1 output215 (.A(\Inst_LUT4AB_switch_matrix.N1BEG2 ),
    .X(N1BEG[2]));
 sg13g2_buf_1 output216 (.A(\Inst_LUT4AB_switch_matrix.N1BEG3 ),
    .X(N1BEG[3]));
 sg13g2_buf_1 output217 (.A(net217),
    .X(N2BEG[0]));
 sg13g2_buf_8 output218 (.A(net218),
    .X(N2BEG[1]));
 sg13g2_buf_8 output219 (.A(net219),
    .X(N2BEG[2]));
 sg13g2_buf_1 output220 (.A(net220),
    .X(N2BEG[3]));
 sg13g2_buf_1 output221 (.A(net221),
    .X(N2BEG[4]));
 sg13g2_buf_1 output222 (.A(\Inst_LUT4AB_switch_matrix.JN2BEG5 ),
    .X(N2BEG[5]));
 sg13g2_buf_1 output223 (.A(net223),
    .X(N2BEG[6]));
 sg13g2_buf_1 output224 (.A(net224),
    .X(N2BEG[7]));
 sg13g2_buf_1 output225 (.A(net225),
    .X(N2BEGb[0]));
 sg13g2_buf_1 output226 (.A(net226),
    .X(N2BEGb[1]));
 sg13g2_buf_1 output227 (.A(net227),
    .X(N2BEGb[2]));
 sg13g2_buf_1 output228 (.A(net228),
    .X(N2BEGb[3]));
 sg13g2_buf_1 output229 (.A(net229),
    .X(N2BEGb[4]));
 sg13g2_buf_1 output230 (.A(net230),
    .X(N2BEGb[5]));
 sg13g2_buf_1 output231 (.A(net231),
    .X(N2BEGb[6]));
 sg13g2_buf_1 output232 (.A(net232),
    .X(N2BEGb[7]));
 sg13g2_buf_1 output233 (.A(net233),
    .X(N4BEG[0]));
 sg13g2_buf_1 output234 (.A(net234),
    .X(N4BEG[10]));
 sg13g2_buf_1 output235 (.A(net235),
    .X(N4BEG[11]));
 sg13g2_buf_1 output236 (.A(net236),
    .X(N4BEG[12]));
 sg13g2_buf_1 output237 (.A(net237),
    .X(N4BEG[13]));
 sg13g2_buf_1 output238 (.A(net238),
    .X(N4BEG[14]));
 sg13g2_buf_1 output239 (.A(\Inst_LUT4AB_switch_matrix.N4BEG3 ),
    .X(N4BEG[15]));
 sg13g2_buf_1 output240 (.A(net240),
    .X(N4BEG[1]));
 sg13g2_buf_1 output241 (.A(net241),
    .X(N4BEG[2]));
 sg13g2_buf_1 output242 (.A(net242),
    .X(N4BEG[3]));
 sg13g2_buf_1 output243 (.A(net243),
    .X(N4BEG[4]));
 sg13g2_buf_1 output244 (.A(net244),
    .X(N4BEG[5]));
 sg13g2_buf_1 output245 (.A(net245),
    .X(N4BEG[6]));
 sg13g2_buf_1 output246 (.A(net246),
    .X(N4BEG[7]));
 sg13g2_buf_1 output247 (.A(net247),
    .X(N4BEG[8]));
 sg13g2_buf_1 output248 (.A(net248),
    .X(N4BEG[9]));
 sg13g2_buf_1 output249 (.A(net249),
    .X(NN4BEG[0]));
 sg13g2_buf_1 output250 (.A(net250),
    .X(NN4BEG[10]));
 sg13g2_buf_1 output251 (.A(net251),
    .X(NN4BEG[11]));
 sg13g2_buf_1 output252 (.A(net252),
    .X(NN4BEG[12]));
 sg13g2_buf_1 output253 (.A(net253),
    .X(NN4BEG[13]));
 sg13g2_buf_1 output254 (.A(\Inst_LUT4AB_switch_matrix.NN4BEG2 ),
    .X(NN4BEG[14]));
 sg13g2_buf_1 output255 (.A(\Inst_LUT4AB_switch_matrix.NN4BEG3 ),
    .X(NN4BEG[15]));
 sg13g2_buf_1 output256 (.A(net256),
    .X(NN4BEG[1]));
 sg13g2_buf_1 output257 (.A(net257),
    .X(NN4BEG[2]));
 sg13g2_buf_1 output258 (.A(net258),
    .X(NN4BEG[3]));
 sg13g2_buf_1 output259 (.A(net259),
    .X(NN4BEG[4]));
 sg13g2_buf_1 output260 (.A(net260),
    .X(NN4BEG[5]));
 sg13g2_buf_1 output261 (.A(net261),
    .X(NN4BEG[6]));
 sg13g2_buf_1 output262 (.A(net262),
    .X(NN4BEG[7]));
 sg13g2_buf_1 output263 (.A(net263),
    .X(NN4BEG[8]));
 sg13g2_buf_1 output264 (.A(net264),
    .X(NN4BEG[9]));
 sg13g2_buf_1 output265 (.A(net265),
    .X(S1BEG[0]));
 sg13g2_buf_1 output266 (.A(net266),
    .X(S1BEG[1]));
 sg13g2_buf_1 output267 (.A(\Inst_LUT4AB_switch_matrix.S1BEG2 ),
    .X(S1BEG[2]));
 sg13g2_buf_1 output268 (.A(\Inst_LUT4AB_switch_matrix.S1BEG3 ),
    .X(S1BEG[3]));
 sg13g2_buf_1 output269 (.A(net269),
    .X(S2BEG[0]));
 sg13g2_buf_1 output270 (.A(net270),
    .X(S2BEG[1]));
 sg13g2_buf_1 output271 (.A(net271),
    .X(S2BEG[2]));
 sg13g2_buf_1 output272 (.A(net272),
    .X(S2BEG[3]));
 sg13g2_buf_1 output273 (.A(net273),
    .X(S2BEG[4]));
 sg13g2_buf_1 output274 (.A(\Inst_LUT4AB_switch_matrix.JS2BEG5 ),
    .X(S2BEG[5]));
 sg13g2_buf_1 output275 (.A(net275),
    .X(S2BEG[6]));
 sg13g2_buf_1 output276 (.A(net276),
    .X(S2BEG[7]));
 sg13g2_buf_1 output277 (.A(net277),
    .X(S2BEGb[0]));
 sg13g2_buf_1 output278 (.A(net278),
    .X(S2BEGb[1]));
 sg13g2_buf_1 output279 (.A(net279),
    .X(S2BEGb[2]));
 sg13g2_buf_1 output280 (.A(net280),
    .X(S2BEGb[3]));
 sg13g2_buf_1 output281 (.A(net281),
    .X(S2BEGb[4]));
 sg13g2_buf_1 output282 (.A(net282),
    .X(S2BEGb[5]));
 sg13g2_buf_1 output283 (.A(net283),
    .X(S2BEGb[6]));
 sg13g2_buf_1 output284 (.A(net284),
    .X(S2BEGb[7]));
 sg13g2_buf_1 output285 (.A(net285),
    .X(S4BEG[0]));
 sg13g2_buf_1 output286 (.A(net286),
    .X(S4BEG[10]));
 sg13g2_buf_1 output287 (.A(net287),
    .X(S4BEG[11]));
 sg13g2_buf_1 output288 (.A(net288),
    .X(S4BEG[12]));
 sg13g2_buf_1 output289 (.A(net289),
    .X(S4BEG[13]));
 sg13g2_buf_1 output290 (.A(net290),
    .X(S4BEG[14]));
 sg13g2_buf_1 output291 (.A(net291),
    .X(S4BEG[15]));
 sg13g2_buf_1 output292 (.A(net292),
    .X(S4BEG[1]));
 sg13g2_buf_1 output293 (.A(net293),
    .X(S4BEG[2]));
 sg13g2_buf_1 output294 (.A(net294),
    .X(S4BEG[3]));
 sg13g2_buf_1 output295 (.A(net295),
    .X(S4BEG[4]));
 sg13g2_buf_1 output296 (.A(net296),
    .X(S4BEG[5]));
 sg13g2_buf_1 output297 (.A(net297),
    .X(S4BEG[6]));
 sg13g2_buf_1 output298 (.A(net298),
    .X(S4BEG[7]));
 sg13g2_buf_1 output299 (.A(net299),
    .X(S4BEG[8]));
 sg13g2_buf_1 output300 (.A(net300),
    .X(S4BEG[9]));
 sg13g2_buf_1 output301 (.A(net301),
    .X(SS4BEG[0]));
 sg13g2_buf_1 output302 (.A(net302),
    .X(SS4BEG[10]));
 sg13g2_buf_1 output303 (.A(net303),
    .X(SS4BEG[11]));
 sg13g2_buf_1 output304 (.A(\Inst_LUT4AB_switch_matrix.SS4BEG0 ),
    .X(SS4BEG[12]));
 sg13g2_buf_1 output305 (.A(net305),
    .X(SS4BEG[13]));
 sg13g2_buf_1 output306 (.A(net306),
    .X(SS4BEG[14]));
 sg13g2_buf_1 output307 (.A(\Inst_LUT4AB_switch_matrix.SS4BEG3 ),
    .X(SS4BEG[15]));
 sg13g2_buf_1 output308 (.A(net308),
    .X(SS4BEG[1]));
 sg13g2_buf_1 output309 (.A(net309),
    .X(SS4BEG[2]));
 sg13g2_buf_1 output310 (.A(net310),
    .X(SS4BEG[3]));
 sg13g2_buf_1 output311 (.A(net311),
    .X(SS4BEG[4]));
 sg13g2_buf_1 output312 (.A(net312),
    .X(SS4BEG[5]));
 sg13g2_buf_1 output313 (.A(net313),
    .X(SS4BEG[6]));
 sg13g2_buf_1 output314 (.A(net314),
    .X(SS4BEG[7]));
 sg13g2_buf_1 output315 (.A(net315),
    .X(SS4BEG[8]));
 sg13g2_buf_1 output316 (.A(net316),
    .X(SS4BEG[9]));
 sg13g2_buf_1 output317 (.A(net317),
    .X(UserCLKo));
 sg13g2_buf_1 output318 (.A(net318),
    .X(W1BEG[0]));
 sg13g2_buf_1 output319 (.A(net319),
    .X(W1BEG[1]));
 sg13g2_buf_1 output320 (.A(net320),
    .X(W1BEG[2]));
 sg13g2_buf_1 output321 (.A(\Inst_LUT4AB_switch_matrix.W1BEG3 ),
    .X(W1BEG[3]));
 sg13g2_buf_1 output322 (.A(net322),
    .X(W2BEG[0]));
 sg13g2_buf_1 output323 (.A(net323),
    .X(W2BEG[1]));
 sg13g2_buf_1 output324 (.A(net324),
    .X(W2BEG[2]));
 sg13g2_buf_1 output325 (.A(net325),
    .X(W2BEG[3]));
 sg13g2_buf_1 output326 (.A(net326),
    .X(W2BEG[4]));
 sg13g2_buf_1 output327 (.A(net327),
    .X(W2BEG[5]));
 sg13g2_buf_1 output328 (.A(net328),
    .X(W2BEG[6]));
 sg13g2_buf_1 output329 (.A(net329),
    .X(W2BEG[7]));
 sg13g2_buf_1 output330 (.A(net330),
    .X(W2BEGb[0]));
 sg13g2_buf_1 output331 (.A(net331),
    .X(W2BEGb[1]));
 sg13g2_buf_1 output332 (.A(net332),
    .X(W2BEGb[2]));
 sg13g2_buf_1 output333 (.A(net333),
    .X(W2BEGb[3]));
 sg13g2_buf_1 output334 (.A(net334),
    .X(W2BEGb[4]));
 sg13g2_buf_1 output335 (.A(net335),
    .X(W2BEGb[5]));
 sg13g2_buf_1 output336 (.A(net336),
    .X(W2BEGb[6]));
 sg13g2_buf_1 output337 (.A(net337),
    .X(W2BEGb[7]));
 sg13g2_buf_1 output338 (.A(net338),
    .X(W6BEG[0]));
 sg13g2_buf_1 output339 (.A(\Inst_LUT4AB_switch_matrix.W6BEG0 ),
    .X(W6BEG[10]));
 sg13g2_buf_1 output340 (.A(\Inst_LUT4AB_switch_matrix.W6BEG1 ),
    .X(W6BEG[11]));
 sg13g2_buf_1 output341 (.A(net341),
    .X(W6BEG[1]));
 sg13g2_buf_1 output342 (.A(net342),
    .X(W6BEG[2]));
 sg13g2_buf_1 output343 (.A(net343),
    .X(W6BEG[3]));
 sg13g2_buf_1 output344 (.A(net344),
    .X(W6BEG[4]));
 sg13g2_buf_1 output345 (.A(net345),
    .X(W6BEG[5]));
 sg13g2_buf_1 output346 (.A(net346),
    .X(W6BEG[6]));
 sg13g2_buf_1 output347 (.A(net347),
    .X(W6BEG[7]));
 sg13g2_buf_1 output348 (.A(net348),
    .X(W6BEG[8]));
 sg13g2_buf_1 output349 (.A(net349),
    .X(W6BEG[9]));
 sg13g2_buf_1 output350 (.A(net350),
    .X(WW4BEG[0]));
 sg13g2_buf_1 output351 (.A(net351),
    .X(WW4BEG[10]));
 sg13g2_buf_1 output352 (.A(net352),
    .X(WW4BEG[11]));
 sg13g2_buf_1 output353 (.A(net353),
    .X(WW4BEG[12]));
 sg13g2_buf_1 output354 (.A(net354),
    .X(WW4BEG[13]));
 sg13g2_buf_1 output355 (.A(net355),
    .X(WW4BEG[14]));
 sg13g2_buf_1 output356 (.A(\Inst_LUT4AB_switch_matrix.WW4BEG3 ),
    .X(WW4BEG[15]));
 sg13g2_buf_1 output357 (.A(net357),
    .X(WW4BEG[1]));
 sg13g2_buf_1 output358 (.A(net358),
    .X(WW4BEG[2]));
 sg13g2_buf_1 output359 (.A(net359),
    .X(WW4BEG[3]));
 sg13g2_buf_1 output360 (.A(net360),
    .X(WW4BEG[4]));
 sg13g2_buf_1 output361 (.A(net361),
    .X(WW4BEG[5]));
 sg13g2_buf_1 output362 (.A(net362),
    .X(WW4BEG[6]));
 sg13g2_buf_1 output363 (.A(net363),
    .X(WW4BEG[7]));
 sg13g2_buf_1 output364 (.A(net364),
    .X(WW4BEG[8]));
 sg13g2_buf_1 output365 (.A(net365),
    .X(WW4BEG[9]));
 sg13g2_tiehi _3052__366 (.L_HI(net366));
 sg13g2_dlygate4sd1_1 rebuffer2 (.A(_0248_),
    .X(net375));
 sg13g2_dlygate4sd1_1 rebuffer3 (.A(_0248_),
    .X(net376));
 sg13g2_dlygate4sd1_1 rebuffer4 (.A(\Inst_LUT4AB_switch_matrix.JW2BEG5 ),
    .X(net377));
 sg13g2_buf_2 rebuffer5 (.A(_0590_),
    .X(net378));
 sg13g2_buf_2 rebuffer6 (.A(_0649_),
    .X(net379));
 sg13g2_buf_2 rebuffer8 (.A(_0640_),
    .X(net381));
 sg13g2_dlygate4sd1_1 rebuffer9 (.A(\Inst_LUT4AB_switch_matrix.E2BEG1 ),
    .X(net382));
 sg13g2_dlygate4sd1_1 rebuffer10 (.A(\Inst_LUT4AB_switch_matrix.E2BEG1 ),
    .X(net383));
 sg13g2_dlygate4sd1_1 rebuffer11 (.A(\Inst_LUT4AB_switch_matrix.JW2BEG2 ),
    .X(net384));
 sg13g2_dlygate4sd1_1 rebuffer12 (.A(_0520_),
    .X(net385));
 sg13g2_dlygate4sd1_1 rebuffer14 (.A(_0638_),
    .X(net387));
 sg13g2_buf_2 rebuffer15 (.A(_0640_),
    .X(net388));
 sg13g2_dlygate4sd1_1 rebuffer16 (.A(_0348_),
    .X(net389));
 sg13g2_fill_1 FILLER_0_334 ();
 sg13g2_fill_2 FILLER_0_361 ();
 sg13g2_fill_2 FILLER_0_421 ();
 sg13g2_fill_1 FILLER_0_423 ();
 sg13g2_fill_2 FILLER_0_457 ();
 sg13g2_fill_2 FILLER_1_8 ();
 sg13g2_fill_1 FILLER_1_27 ();
 sg13g2_fill_1 FILLER_1_49 ();
 sg13g2_fill_2 FILLER_1_232 ();
 sg13g2_fill_1 FILLER_1_234 ();
 sg13g2_fill_2 FILLER_1_252 ();
 sg13g2_fill_1 FILLER_1_315 ();
 sg13g2_fill_1 FILLER_1_333 ();
 sg13g2_fill_1 FILLER_1_362 ();
 sg13g2_fill_2 FILLER_2_0 ();
 sg13g2_fill_1 FILLER_2_2 ();
 sg13g2_fill_2 FILLER_2_20 ();
 sg13g2_fill_2 FILLER_2_39 ();
 sg13g2_fill_1 FILLER_2_84 ();
 sg13g2_fill_2 FILLER_2_167 ();
 sg13g2_fill_2 FILLER_2_174 ();
 sg13g2_fill_1 FILLER_2_176 ();
 sg13g2_fill_1 FILLER_2_198 ();
 sg13g2_fill_1 FILLER_2_220 ();
 sg13g2_fill_1 FILLER_2_225 ();
 sg13g2_fill_2 FILLER_2_247 ();
 sg13g2_fill_2 FILLER_2_270 ();
 sg13g2_fill_2 FILLER_2_276 ();
 sg13g2_fill_2 FILLER_2_307 ();
 sg13g2_fill_1 FILLER_2_309 ();
 sg13g2_fill_1 FILLER_2_359 ();
 sg13g2_fill_2 FILLER_2_398 ();
 sg13g2_fill_1 FILLER_2_400 ();
 sg13g2_fill_1 FILLER_2_422 ();
 sg13g2_fill_1 FILLER_2_454 ();
 sg13g2_fill_2 FILLER_3_0 ();
 sg13g2_fill_2 FILLER_3_19 ();
 sg13g2_fill_2 FILLER_3_49 ();
 sg13g2_fill_1 FILLER_3_51 ();
 sg13g2_fill_2 FILLER_3_140 ();
 sg13g2_fill_1 FILLER_3_142 ();
 sg13g2_fill_2 FILLER_3_153 ();
 sg13g2_fill_2 FILLER_3_235 ();
 sg13g2_fill_1 FILLER_3_237 ();
 sg13g2_fill_1 FILLER_3_276 ();
 sg13g2_fill_2 FILLER_3_335 ();
 sg13g2_fill_1 FILLER_3_337 ();
 sg13g2_fill_1 FILLER_3_400 ();
 sg13g2_fill_2 FILLER_3_452 ();
 sg13g2_fill_1 FILLER_3_454 ();
 sg13g2_fill_2 FILLER_4_0 ();
 sg13g2_fill_1 FILLER_4_19 ();
 sg13g2_fill_2 FILLER_4_78 ();
 sg13g2_fill_2 FILLER_4_118 ();
 sg13g2_fill_1 FILLER_4_120 ();
 sg13g2_fill_2 FILLER_4_172 ();
 sg13g2_fill_2 FILLER_4_302 ();
 sg13g2_fill_1 FILLER_4_312 ();
 sg13g2_fill_2 FILLER_4_360 ();
 sg13g2_fill_1 FILLER_4_362 ();
 sg13g2_fill_1 FILLER_4_384 ();
 sg13g2_fill_1 FILLER_4_403 ();
 sg13g2_fill_2 FILLER_4_452 ();
 sg13g2_fill_1 FILLER_4_454 ();
 sg13g2_fill_1 FILLER_5_0 ();
 sg13g2_fill_1 FILLER_5_114 ();
 sg13g2_fill_1 FILLER_5_174 ();
 sg13g2_fill_1 FILLER_5_215 ();
 sg13g2_fill_2 FILLER_5_249 ();
 sg13g2_fill_2 FILLER_5_256 ();
 sg13g2_fill_1 FILLER_5_258 ();
 sg13g2_fill_2 FILLER_5_284 ();
 sg13g2_fill_1 FILLER_5_286 ();
 sg13g2_fill_2 FILLER_5_360 ();
 sg13g2_fill_1 FILLER_5_362 ();
 sg13g2_fill_2 FILLER_5_380 ();
 sg13g2_fill_1 FILLER_5_382 ();
 sg13g2_fill_1 FILLER_6_20 ();
 sg13g2_fill_2 FILLER_6_60 ();
 sg13g2_fill_1 FILLER_6_62 ();
 sg13g2_fill_1 FILLER_6_82 ();
 sg13g2_fill_2 FILLER_6_158 ();
 sg13g2_fill_1 FILLER_6_160 ();
 sg13g2_fill_1 FILLER_6_189 ();
 sg13g2_fill_1 FILLER_6_248 ();
 sg13g2_fill_2 FILLER_6_254 ();
 sg13g2_fill_2 FILLER_6_295 ();
 sg13g2_fill_1 FILLER_6_297 ();
 sg13g2_fill_1 FILLER_6_320 ();
 sg13g2_fill_1 FILLER_6_342 ();
 sg13g2_fill_1 FILLER_6_377 ();
 sg13g2_fill_2 FILLER_6_457 ();
 sg13g2_fill_2 FILLER_7_0 ();
 sg13g2_fill_1 FILLER_7_2 ();
 sg13g2_fill_1 FILLER_7_20 ();
 sg13g2_fill_2 FILLER_7_54 ();
 sg13g2_fill_2 FILLER_7_60 ();
 sg13g2_fill_1 FILLER_7_70 ();
 sg13g2_fill_2 FILLER_7_96 ();
 sg13g2_fill_1 FILLER_7_182 ();
 sg13g2_fill_1 FILLER_7_242 ();
 sg13g2_fill_1 FILLER_7_269 ();
 sg13g2_fill_2 FILLER_7_287 ();
 sg13g2_fill_2 FILLER_7_352 ();
 sg13g2_fill_2 FILLER_7_371 ();
 sg13g2_fill_1 FILLER_7_373 ();
 sg13g2_fill_2 FILLER_7_389 ();
 sg13g2_fill_1 FILLER_7_391 ();
 sg13g2_fill_2 FILLER_7_398 ();
 sg13g2_fill_1 FILLER_7_400 ();
 sg13g2_fill_2 FILLER_7_418 ();
 sg13g2_fill_1 FILLER_7_454 ();
 sg13g2_fill_1 FILLER_8_0 ();
 sg13g2_fill_1 FILLER_8_63 ();
 sg13g2_fill_1 FILLER_8_68 ();
 sg13g2_fill_2 FILLER_8_111 ();
 sg13g2_fill_1 FILLER_8_113 ();
 sg13g2_fill_1 FILLER_8_189 ();
 sg13g2_fill_1 FILLER_8_266 ();
 sg13g2_fill_2 FILLER_8_296 ();
 sg13g2_fill_1 FILLER_8_298 ();
 sg13g2_fill_1 FILLER_8_304 ();
 sg13g2_fill_2 FILLER_8_326 ();
 sg13g2_fill_1 FILLER_8_328 ();
 sg13g2_fill_2 FILLER_8_367 ();
 sg13g2_fill_1 FILLER_8_369 ();
 sg13g2_fill_2 FILLER_8_424 ();
 sg13g2_fill_1 FILLER_8_426 ();
 sg13g2_fill_2 FILLER_8_435 ();
 sg13g2_fill_1 FILLER_8_437 ();
 sg13g2_fill_2 FILLER_8_456 ();
 sg13g2_fill_1 FILLER_8_458 ();
 sg13g2_fill_1 FILLER_9_109 ();
 sg13g2_fill_1 FILLER_9_152 ();
 sg13g2_fill_2 FILLER_9_269 ();
 sg13g2_fill_1 FILLER_9_307 ();
 sg13g2_fill_2 FILLER_9_329 ();
 sg13g2_fill_1 FILLER_9_331 ();
 sg13g2_fill_2 FILLER_9_364 ();
 sg13g2_fill_1 FILLER_9_424 ();
 sg13g2_fill_2 FILLER_9_456 ();
 sg13g2_fill_1 FILLER_9_458 ();
 sg13g2_fill_2 FILLER_10_21 ();
 sg13g2_fill_1 FILLER_10_46 ();
 sg13g2_fill_2 FILLER_10_67 ();
 sg13g2_fill_1 FILLER_10_69 ();
 sg13g2_fill_2 FILLER_10_87 ();
 sg13g2_fill_1 FILLER_10_143 ();
 sg13g2_fill_2 FILLER_10_268 ();
 sg13g2_fill_2 FILLER_10_274 ();
 sg13g2_fill_2 FILLER_10_329 ();
 sg13g2_fill_1 FILLER_10_331 ();
 sg13g2_fill_1 FILLER_10_364 ();
 sg13g2_fill_2 FILLER_10_388 ();
 sg13g2_fill_2 FILLER_10_416 ();
 sg13g2_fill_1 FILLER_10_418 ();
 sg13g2_fill_2 FILLER_11_0 ();
 sg13g2_fill_1 FILLER_11_38 ();
 sg13g2_fill_2 FILLER_11_67 ();
 sg13g2_fill_1 FILLER_11_128 ();
 sg13g2_fill_2 FILLER_11_182 ();
 sg13g2_fill_1 FILLER_11_184 ();
 sg13g2_fill_1 FILLER_11_193 ();
 sg13g2_decap_4 FILLER_11_247 ();
 sg13g2_fill_2 FILLER_11_251 ();
 sg13g2_fill_2 FILLER_11_302 ();
 sg13g2_fill_1 FILLER_11_304 ();
 sg13g2_fill_2 FILLER_11_330 ();
 sg13g2_fill_1 FILLER_11_332 ();
 sg13g2_fill_2 FILLER_11_379 ();
 sg13g2_fill_1 FILLER_11_438 ();
 sg13g2_fill_2 FILLER_11_456 ();
 sg13g2_fill_1 FILLER_11_458 ();
 sg13g2_fill_2 FILLER_12_0 ();
 sg13g2_fill_2 FILLER_12_163 ();
 sg13g2_fill_2 FILLER_12_215 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_4 FILLER_12_245 ();
 sg13g2_fill_1 FILLER_12_249 ();
 sg13g2_fill_1 FILLER_12_377 ();
 sg13g2_fill_2 FILLER_12_395 ();
 sg13g2_fill_2 FILLER_12_439 ();
 sg13g2_fill_1 FILLER_13_4 ();
 sg13g2_fill_1 FILLER_13_98 ();
 sg13g2_fill_2 FILLER_13_107 ();
 sg13g2_fill_1 FILLER_13_109 ();
 sg13g2_fill_1 FILLER_13_148 ();
 sg13g2_fill_1 FILLER_13_201 ();
 sg13g2_fill_2 FILLER_13_247 ();
 sg13g2_decap_8 FILLER_13_253 ();
 sg13g2_decap_4 FILLER_13_260 ();
 sg13g2_fill_1 FILLER_13_268 ();
 sg13g2_fill_1 FILLER_13_373 ();
 sg13g2_fill_2 FILLER_13_410 ();
 sg13g2_fill_1 FILLER_13_430 ();
 sg13g2_fill_2 FILLER_13_452 ();
 sg13g2_fill_2 FILLER_14_0 ();
 sg13g2_fill_1 FILLER_14_19 ();
 sg13g2_fill_2 FILLER_14_92 ();
 sg13g2_fill_1 FILLER_14_135 ();
 sg13g2_fill_2 FILLER_14_173 ();
 sg13g2_fill_2 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_219 ();
 sg13g2_decap_8 FILLER_14_226 ();
 sg13g2_fill_1 FILLER_14_233 ();
 sg13g2_fill_1 FILLER_14_255 ();
 sg13g2_fill_1 FILLER_14_397 ();
 sg13g2_fill_2 FILLER_14_436 ();
 sg13g2_fill_1 FILLER_15_0 ();
 sg13g2_fill_2 FILLER_15_22 ();
 sg13g2_fill_2 FILLER_15_49 ();
 sg13g2_fill_1 FILLER_15_70 ();
 sg13g2_fill_2 FILLER_15_113 ();
 sg13g2_fill_1 FILLER_15_123 ();
 sg13g2_fill_1 FILLER_15_162 ();
 sg13g2_fill_1 FILLER_15_223 ();
 sg13g2_decap_4 FILLER_15_312 ();
 sg13g2_fill_2 FILLER_15_320 ();
 sg13g2_fill_1 FILLER_15_354 ();
 sg13g2_fill_2 FILLER_16_0 ();
 sg13g2_fill_1 FILLER_16_2 ();
 sg13g2_fill_2 FILLER_16_47 ();
 sg13g2_fill_1 FILLER_16_64 ();
 sg13g2_fill_2 FILLER_16_86 ();
 sg13g2_fill_1 FILLER_16_162 ();
 sg13g2_decap_8 FILLER_16_260 ();
 sg13g2_decap_8 FILLER_16_267 ();
 sg13g2_decap_8 FILLER_16_274 ();
 sg13g2_decap_8 FILLER_16_281 ();
 sg13g2_decap_8 FILLER_16_288 ();
 sg13g2_fill_1 FILLER_16_295 ();
 sg13g2_decap_8 FILLER_16_304 ();
 sg13g2_decap_4 FILLER_16_311 ();
 sg13g2_fill_2 FILLER_16_315 ();
 sg13g2_fill_2 FILLER_16_355 ();
 sg13g2_fill_1 FILLER_16_357 ();
 sg13g2_fill_1 FILLER_16_402 ();
 sg13g2_fill_1 FILLER_17_38 ();
 sg13g2_fill_1 FILLER_17_44 ();
 sg13g2_fill_1 FILLER_17_66 ();
 sg13g2_fill_2 FILLER_17_138 ();
 sg13g2_fill_1 FILLER_17_140 ();
 sg13g2_fill_2 FILLER_17_253 ();
 sg13g2_fill_1 FILLER_17_255 ();
 sg13g2_fill_1 FILLER_17_277 ();
 sg13g2_fill_1 FILLER_17_304 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_4 FILLER_17_329 ();
 sg13g2_fill_1 FILLER_17_333 ();
 sg13g2_fill_1 FILLER_17_432 ();
 sg13g2_fill_2 FILLER_18_0 ();
 sg13g2_fill_2 FILLER_18_38 ();
 sg13g2_fill_1 FILLER_18_45 ();
 sg13g2_fill_2 FILLER_18_61 ();
 sg13g2_fill_1 FILLER_18_103 ();
 sg13g2_fill_2 FILLER_18_133 ();
 sg13g2_fill_1 FILLER_18_135 ();
 sg13g2_fill_1 FILLER_18_181 ();
 sg13g2_decap_8 FILLER_18_263 ();
 sg13g2_fill_2 FILLER_18_270 ();
 sg13g2_fill_2 FILLER_18_358 ();
 sg13g2_fill_1 FILLER_18_360 ();
 sg13g2_fill_2 FILLER_18_412 ();
 sg13g2_fill_1 FILLER_18_430 ();
 sg13g2_fill_2 FILLER_18_445 ();
 sg13g2_fill_2 FILLER_18_456 ();
 sg13g2_fill_1 FILLER_18_458 ();
 sg13g2_fill_2 FILLER_19_0 ();
 sg13g2_fill_1 FILLER_19_2 ();
 sg13g2_fill_1 FILLER_19_37 ();
 sg13g2_fill_2 FILLER_19_43 ();
 sg13g2_fill_2 FILLER_19_60 ();
 sg13g2_fill_1 FILLER_19_62 ();
 sg13g2_fill_1 FILLER_19_73 ();
 sg13g2_fill_1 FILLER_19_95 ();
 sg13g2_fill_2 FILLER_19_106 ();
 sg13g2_fill_2 FILLER_19_175 ();
 sg13g2_fill_1 FILLER_19_235 ();
 sg13g2_fill_1 FILLER_19_253 ();
 sg13g2_decap_8 FILLER_19_279 ();
 sg13g2_decap_4 FILLER_19_286 ();
 sg13g2_fill_1 FILLER_19_300 ();
 sg13g2_decap_8 FILLER_19_318 ();
 sg13g2_decap_4 FILLER_19_325 ();
 sg13g2_fill_2 FILLER_19_329 ();
 sg13g2_decap_4 FILLER_19_348 ();
 sg13g2_fill_1 FILLER_19_352 ();
 sg13g2_fill_2 FILLER_19_452 ();
 sg13g2_fill_1 FILLER_19_454 ();
 sg13g2_fill_2 FILLER_20_4 ();
 sg13g2_fill_1 FILLER_20_6 ();
 sg13g2_fill_2 FILLER_20_41 ();
 sg13g2_fill_2 FILLER_20_122 ();
 sg13g2_fill_1 FILLER_20_162 ();
 sg13g2_fill_1 FILLER_20_202 ();
 sg13g2_decap_8 FILLER_20_224 ();
 sg13g2_decap_4 FILLER_20_231 ();
 sg13g2_fill_2 FILLER_20_249 ();
 sg13g2_fill_2 FILLER_20_256 ();
 sg13g2_fill_1 FILLER_20_285 ();
 sg13g2_fill_1 FILLER_20_290 ();
 sg13g2_fill_1 FILLER_20_296 ();
 sg13g2_decap_8 FILLER_20_301 ();
 sg13g2_fill_1 FILLER_20_308 ();
 sg13g2_decap_4 FILLER_20_334 ();
 sg13g2_fill_1 FILLER_20_338 ();
 sg13g2_fill_2 FILLER_20_364 ();
 sg13g2_fill_2 FILLER_20_383 ();
 sg13g2_fill_1 FILLER_20_385 ();
 sg13g2_fill_1 FILLER_20_424 ();
 sg13g2_fill_2 FILLER_21_4 ();
 sg13g2_fill_1 FILLER_21_6 ();
 sg13g2_fill_2 FILLER_21_41 ();
 sg13g2_fill_1 FILLER_21_48 ();
 sg13g2_fill_1 FILLER_21_83 ();
 sg13g2_fill_1 FILLER_21_88 ();
 sg13g2_fill_2 FILLER_21_165 ();
 sg13g2_decap_4 FILLER_21_188 ();
 sg13g2_decap_4 FILLER_21_200 ();
 sg13g2_fill_1 FILLER_21_204 ();
 sg13g2_decap_8 FILLER_21_222 ();
 sg13g2_fill_1 FILLER_21_229 ();
 sg13g2_fill_2 FILLER_21_272 ();
 sg13g2_fill_1 FILLER_21_274 ();
 sg13g2_fill_2 FILLER_21_300 ();
 sg13g2_decap_4 FILLER_21_306 ();
 sg13g2_fill_1 FILLER_21_310 ();
 sg13g2_decap_4 FILLER_21_328 ();
 sg13g2_decap_4 FILLER_21_335 ();
 sg13g2_fill_2 FILLER_21_339 ();
 sg13g2_fill_2 FILLER_21_379 ();
 sg13g2_fill_2 FILLER_21_424 ();
 sg13g2_fill_1 FILLER_21_426 ();
 sg13g2_fill_2 FILLER_21_431 ();
 sg13g2_fill_2 FILLER_21_457 ();
 sg13g2_fill_1 FILLER_22_29 ();
 sg13g2_fill_1 FILLER_22_51 ();
 sg13g2_fill_1 FILLER_22_87 ();
 sg13g2_decap_8 FILLER_22_143 ();
 sg13g2_decap_8 FILLER_22_167 ();
 sg13g2_fill_1 FILLER_22_174 ();
 sg13g2_fill_1 FILLER_22_179 ();
 sg13g2_fill_2 FILLER_22_207 ();
 sg13g2_fill_2 FILLER_22_247 ();
 sg13g2_decap_4 FILLER_22_305 ();
 sg13g2_fill_1 FILLER_22_309 ();
 sg13g2_fill_1 FILLER_22_365 ();
 sg13g2_fill_1 FILLER_22_434 ();
 sg13g2_fill_2 FILLER_22_452 ();
 sg13g2_fill_1 FILLER_22_454 ();
 sg13g2_fill_2 FILLER_23_12 ();
 sg13g2_fill_2 FILLER_23_31 ();
 sg13g2_fill_1 FILLER_23_42 ();
 sg13g2_fill_1 FILLER_23_125 ();
 sg13g2_decap_8 FILLER_23_143 ();
 sg13g2_fill_2 FILLER_23_150 ();
 sg13g2_fill_2 FILLER_23_177 ();
 sg13g2_decap_4 FILLER_23_200 ();
 sg13g2_decap_8 FILLER_23_225 ();
 sg13g2_fill_1 FILLER_23_232 ();
 sg13g2_decap_8 FILLER_23_245 ();
 sg13g2_decap_8 FILLER_23_269 ();
 sg13g2_fill_1 FILLER_23_310 ();
 sg13g2_fill_2 FILLER_23_353 ();
 sg13g2_fill_1 FILLER_23_355 ();
 sg13g2_decap_4 FILLER_23_360 ();
 sg13g2_fill_1 FILLER_23_364 ();
 sg13g2_fill_2 FILLER_23_430 ();
 sg13g2_fill_1 FILLER_23_432 ();
 sg13g2_fill_2 FILLER_24_0 ();
 sg13g2_fill_2 FILLER_24_23 ();
 sg13g2_fill_1 FILLER_24_82 ();
 sg13g2_fill_2 FILLER_24_125 ();
 sg13g2_decap_4 FILLER_24_130 ();
 sg13g2_fill_2 FILLER_24_172 ();
 sg13g2_fill_2 FILLER_24_195 ();
 sg13g2_fill_1 FILLER_24_197 ();
 sg13g2_fill_2 FILLER_24_208 ();
 sg13g2_fill_2 FILLER_24_227 ();
 sg13g2_decap_8 FILLER_24_277 ();
 sg13g2_decap_4 FILLER_24_305 ();
 sg13g2_fill_1 FILLER_24_309 ();
 sg13g2_decap_4 FILLER_24_330 ();
 sg13g2_fill_1 FILLER_24_334 ();
 sg13g2_fill_2 FILLER_25_0 ();
 sg13g2_fill_1 FILLER_25_19 ();
 sg13g2_fill_1 FILLER_25_39 ();
 sg13g2_fill_2 FILLER_25_57 ();
 sg13g2_fill_1 FILLER_25_69 ();
 sg13g2_fill_1 FILLER_25_75 ();
 sg13g2_fill_1 FILLER_25_89 ();
 sg13g2_decap_4 FILLER_25_116 ();
 sg13g2_fill_1 FILLER_25_120 ();
 sg13g2_fill_2 FILLER_25_138 ();
 sg13g2_fill_1 FILLER_25_181 ();
 sg13g2_fill_2 FILLER_25_238 ();
 sg13g2_fill_2 FILLER_25_282 ();
 sg13g2_decap_8 FILLER_25_318 ();
 sg13g2_fill_1 FILLER_25_325 ();
 sg13g2_decap_8 FILLER_25_364 ();
 sg13g2_decap_8 FILLER_25_371 ();
 sg13g2_decap_8 FILLER_25_378 ();
 sg13g2_fill_2 FILLER_25_385 ();
 sg13g2_fill_2 FILLER_25_415 ();
 sg13g2_fill_2 FILLER_26_0 ();
 sg13g2_fill_1 FILLER_26_19 ();
 sg13g2_fill_1 FILLER_26_35 ();
 sg13g2_fill_2 FILLER_26_57 ();
 sg13g2_fill_1 FILLER_26_98 ();
 sg13g2_decap_4 FILLER_26_122 ();
 sg13g2_fill_1 FILLER_26_126 ();
 sg13g2_decap_8 FILLER_26_137 ();
 sg13g2_fill_2 FILLER_26_144 ();
 sg13g2_fill_1 FILLER_26_146 ();
 sg13g2_fill_2 FILLER_26_172 ();
 sg13g2_decap_4 FILLER_26_195 ();
 sg13g2_fill_1 FILLER_26_208 ();
 sg13g2_fill_2 FILLER_26_214 ();
 sg13g2_fill_2 FILLER_26_237 ();
 sg13g2_decap_8 FILLER_26_249 ();
 sg13g2_fill_2 FILLER_26_277 ();
 sg13g2_fill_1 FILLER_26_279 ();
 sg13g2_decap_8 FILLER_26_297 ();
 sg13g2_decap_4 FILLER_26_304 ();
 sg13g2_fill_1 FILLER_26_325 ();
 sg13g2_fill_2 FILLER_26_355 ();
 sg13g2_decap_8 FILLER_26_378 ();
 sg13g2_decap_4 FILLER_26_385 ();
 sg13g2_fill_1 FILLER_26_411 ();
 sg13g2_fill_1 FILLER_26_454 ();
 sg13g2_fill_2 FILLER_27_0 ();
 sg13g2_fill_1 FILLER_27_19 ();
 sg13g2_fill_1 FILLER_27_64 ();
 sg13g2_fill_2 FILLER_27_82 ();
 sg13g2_decap_4 FILLER_27_146 ();
 sg13g2_decap_8 FILLER_27_193 ();
 sg13g2_decap_8 FILLER_27_200 ();
 sg13g2_fill_1 FILLER_27_207 ();
 sg13g2_decap_8 FILLER_27_225 ();
 sg13g2_fill_1 FILLER_27_236 ();
 sg13g2_decap_8 FILLER_27_258 ();
 sg13g2_decap_8 FILLER_27_265 ();
 sg13g2_decap_8 FILLER_27_272 ();
 sg13g2_decap_8 FILLER_27_279 ();
 sg13g2_fill_1 FILLER_27_286 ();
 sg13g2_fill_1 FILLER_27_325 ();
 sg13g2_fill_2 FILLER_27_331 ();
 sg13g2_fill_1 FILLER_27_333 ();
 sg13g2_fill_2 FILLER_27_355 ();
 sg13g2_fill_1 FILLER_27_357 ();
 sg13g2_fill_1 FILLER_27_425 ();
 sg13g2_fill_2 FILLER_28_8 ();
 sg13g2_fill_2 FILLER_28_22 ();
 sg13g2_fill_2 FILLER_28_47 ();
 sg13g2_fill_2 FILLER_28_104 ();
 sg13g2_decap_4 FILLER_28_118 ();
 sg13g2_fill_1 FILLER_28_122 ();
 sg13g2_fill_2 FILLER_28_131 ();
 sg13g2_decap_4 FILLER_28_143 ();
 sg13g2_decap_8 FILLER_28_164 ();
 sg13g2_decap_8 FILLER_28_171 ();
 sg13g2_fill_2 FILLER_28_178 ();
 sg13g2_fill_2 FILLER_28_197 ();
 sg13g2_fill_1 FILLER_28_241 ();
 sg13g2_decap_8 FILLER_28_268 ();
 sg13g2_decap_4 FILLER_28_275 ();
 sg13g2_fill_1 FILLER_28_279 ();
 sg13g2_fill_2 FILLER_28_303 ();
 sg13g2_fill_2 FILLER_28_322 ();
 sg13g2_fill_2 FILLER_28_345 ();
 sg13g2_fill_1 FILLER_28_347 ();
 sg13g2_fill_2 FILLER_28_426 ();
 sg13g2_fill_1 FILLER_28_428 ();
 sg13g2_fill_2 FILLER_28_433 ();
 sg13g2_fill_2 FILLER_28_452 ();
 sg13g2_fill_1 FILLER_28_454 ();
 sg13g2_fill_2 FILLER_29_4 ();
 sg13g2_fill_1 FILLER_29_40 ();
 sg13g2_fill_2 FILLER_29_105 ();
 sg13g2_fill_2 FILLER_29_154 ();
 sg13g2_fill_2 FILLER_29_173 ();
 sg13g2_fill_1 FILLER_29_175 ();
 sg13g2_decap_4 FILLER_29_193 ();
 sg13g2_decap_4 FILLER_29_218 ();
 sg13g2_fill_2 FILLER_29_222 ();
 sg13g2_fill_2 FILLER_29_228 ();
 sg13g2_fill_2 FILLER_29_255 ();
 sg13g2_fill_2 FILLER_29_268 ();
 sg13g2_fill_2 FILLER_29_331 ();
 sg13g2_decap_8 FILLER_29_358 ();
 sg13g2_fill_2 FILLER_29_365 ();
 sg13g2_fill_1 FILLER_29_367 ();
 sg13g2_fill_1 FILLER_29_385 ();
 sg13g2_fill_2 FILLER_29_401 ();
 sg13g2_fill_1 FILLER_29_403 ();
 sg13g2_fill_1 FILLER_29_447 ();
 sg13g2_fill_1 FILLER_29_458 ();
 sg13g2_fill_2 FILLER_30_61 ();
 sg13g2_fill_2 FILLER_30_80 ();
 sg13g2_fill_1 FILLER_30_82 ();
 sg13g2_decap_8 FILLER_30_117 ();
 sg13g2_decap_4 FILLER_30_128 ();
 sg13g2_fill_2 FILLER_30_132 ();
 sg13g2_decap_4 FILLER_30_173 ();
 sg13g2_fill_1 FILLER_30_186 ();
 sg13g2_decap_4 FILLER_30_199 ();
 sg13g2_fill_2 FILLER_30_229 ();
 sg13g2_fill_1 FILLER_30_231 ();
 sg13g2_decap_4 FILLER_30_249 ();
 sg13g2_fill_1 FILLER_30_258 ();
 sg13g2_decap_4 FILLER_30_292 ();
 sg13g2_fill_2 FILLER_30_362 ();
 sg13g2_fill_1 FILLER_30_364 ();
 sg13g2_fill_1 FILLER_30_386 ();
 sg13g2_decap_8 FILLER_30_407 ();
 sg13g2_fill_2 FILLER_30_435 ();
 sg13g2_fill_1 FILLER_30_437 ();
 sg13g2_fill_2 FILLER_31_66 ();
 sg13g2_fill_1 FILLER_31_68 ();
 sg13g2_fill_2 FILLER_31_122 ();
 sg13g2_fill_1 FILLER_31_124 ();
 sg13g2_decap_8 FILLER_31_161 ();
 sg13g2_fill_1 FILLER_31_168 ();
 sg13g2_fill_2 FILLER_31_173 ();
 sg13g2_fill_2 FILLER_31_190 ();
 sg13g2_fill_1 FILLER_31_192 ();
 sg13g2_fill_1 FILLER_31_210 ();
 sg13g2_decap_8 FILLER_31_232 ();
 sg13g2_fill_1 FILLER_31_256 ();
 sg13g2_fill_2 FILLER_31_282 ();
 sg13g2_fill_1 FILLER_31_284 ();
 sg13g2_decap_4 FILLER_31_297 ();
 sg13g2_decap_8 FILLER_31_309 ();
 sg13g2_decap_8 FILLER_31_316 ();
 sg13g2_decap_4 FILLER_31_323 ();
 sg13g2_fill_2 FILLER_31_365 ();
 sg13g2_fill_1 FILLER_31_367 ();
 sg13g2_decap_8 FILLER_31_372 ();
 sg13g2_decap_8 FILLER_31_379 ();
 sg13g2_fill_1 FILLER_31_448 ();
 sg13g2_fill_1 FILLER_31_458 ();
 sg13g2_fill_2 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_23 ();
 sg13g2_decap_8 FILLER_32_30 ();
 sg13g2_decap_4 FILLER_32_37 ();
 sg13g2_decap_4 FILLER_32_66 ();
 sg13g2_decap_4 FILLER_32_91 ();
 sg13g2_fill_1 FILLER_32_95 ();
 sg13g2_decap_4 FILLER_32_106 ();
 sg13g2_fill_2 FILLER_32_110 ();
 sg13g2_fill_2 FILLER_32_133 ();
 sg13g2_fill_1 FILLER_32_135 ();
 sg13g2_fill_1 FILLER_32_147 ();
 sg13g2_fill_1 FILLER_32_153 ();
 sg13g2_decap_4 FILLER_32_159 ();
 sg13g2_fill_1 FILLER_32_163 ();
 sg13g2_fill_1 FILLER_32_217 ();
 sg13g2_fill_1 FILLER_32_268 ();
 sg13g2_decap_8 FILLER_32_307 ();
 sg13g2_fill_1 FILLER_32_314 ();
 sg13g2_fill_1 FILLER_32_319 ();
 sg13g2_decap_4 FILLER_32_324 ();
 sg13g2_fill_2 FILLER_32_328 ();
 sg13g2_fill_2 FILLER_32_431 ();
 sg13g2_fill_1 FILLER_32_458 ();
 sg13g2_fill_2 FILLER_33_4 ();
 sg13g2_fill_1 FILLER_33_6 ();
 sg13g2_decap_4 FILLER_33_93 ();
 sg13g2_fill_1 FILLER_33_97 ();
 sg13g2_decap_4 FILLER_33_123 ();
 sg13g2_fill_2 FILLER_33_148 ();
 sg13g2_fill_1 FILLER_33_150 ();
 sg13g2_fill_2 FILLER_33_171 ();
 sg13g2_decap_8 FILLER_33_191 ();
 sg13g2_decap_8 FILLER_33_198 ();
 sg13g2_decap_8 FILLER_33_205 ();
 sg13g2_fill_2 FILLER_33_212 ();
 sg13g2_fill_1 FILLER_33_214 ();
 sg13g2_fill_2 FILLER_33_236 ();
 sg13g2_fill_2 FILLER_33_257 ();
 sg13g2_fill_2 FILLER_33_284 ();
 sg13g2_fill_2 FILLER_33_290 ();
 sg13g2_decap_8 FILLER_33_338 ();
 sg13g2_fill_2 FILLER_33_345 ();
 sg13g2_fill_2 FILLER_33_377 ();
 sg13g2_fill_1 FILLER_33_438 ();
 sg13g2_fill_1 FILLER_34_39 ();
 sg13g2_fill_1 FILLER_34_108 ();
 sg13g2_fill_2 FILLER_34_113 ();
 sg13g2_decap_8 FILLER_34_120 ();
 sg13g2_fill_1 FILLER_34_127 ();
 sg13g2_fill_1 FILLER_34_149 ();
 sg13g2_fill_2 FILLER_34_179 ();
 sg13g2_fill_1 FILLER_34_215 ();
 sg13g2_fill_2 FILLER_34_243 ();
 sg13g2_fill_2 FILLER_34_253 ();
 sg13g2_fill_2 FILLER_34_261 ();
 sg13g2_fill_1 FILLER_34_284 ();
 sg13g2_fill_2 FILLER_34_350 ();
 sg13g2_fill_2 FILLER_34_386 ();
 sg13g2_fill_2 FILLER_34_440 ();
 sg13g2_fill_2 FILLER_35_0 ();
 sg13g2_fill_1 FILLER_35_2 ();
 sg13g2_fill_2 FILLER_35_20 ();
 sg13g2_fill_1 FILLER_35_22 ();
 sg13g2_fill_2 FILLER_35_37 ();
 sg13g2_fill_1 FILLER_35_39 ();
 sg13g2_decap_8 FILLER_35_114 ();
 sg13g2_fill_1 FILLER_35_121 ();
 sg13g2_fill_1 FILLER_35_139 ();
 sg13g2_fill_1 FILLER_35_216 ();
 sg13g2_fill_2 FILLER_35_238 ();
 sg13g2_fill_1 FILLER_35_240 ();
 sg13g2_decap_8 FILLER_35_300 ();
 sg13g2_fill_1 FILLER_35_307 ();
 sg13g2_fill_2 FILLER_35_367 ();
 sg13g2_fill_1 FILLER_35_399 ();
 sg13g2_fill_2 FILLER_35_417 ();
 sg13g2_fill_2 FILLER_36_0 ();
 sg13g2_fill_2 FILLER_36_31 ();
 sg13g2_fill_1 FILLER_36_33 ();
 sg13g2_decap_8 FILLER_36_43 ();
 sg13g2_decap_4 FILLER_36_50 ();
 sg13g2_fill_1 FILLER_36_54 ();
 sg13g2_fill_1 FILLER_36_60 ();
 sg13g2_fill_2 FILLER_36_82 ();
 sg13g2_fill_1 FILLER_36_84 ();
 sg13g2_decap_4 FILLER_36_110 ();
 sg13g2_decap_8 FILLER_36_131 ();
 sg13g2_decap_4 FILLER_36_143 ();
 sg13g2_decap_8 FILLER_36_173 ();
 sg13g2_decap_4 FILLER_36_180 ();
 sg13g2_fill_2 FILLER_36_192 ();
 sg13g2_decap_8 FILLER_36_221 ();
 sg13g2_decap_8 FILLER_36_228 ();
 sg13g2_decap_8 FILLER_36_281 ();
 sg13g2_fill_2 FILLER_36_309 ();
 sg13g2_fill_1 FILLER_36_311 ();
 sg13g2_decap_4 FILLER_36_324 ();
 sg13g2_fill_2 FILLER_36_328 ();
 sg13g2_fill_2 FILLER_36_362 ();
 sg13g2_fill_1 FILLER_36_364 ();
 sg13g2_fill_2 FILLER_36_390 ();
 sg13g2_fill_1 FILLER_36_392 ();
 sg13g2_fill_2 FILLER_36_457 ();
 sg13g2_decap_8 FILLER_37_55 ();
 sg13g2_fill_1 FILLER_37_62 ();
 sg13g2_decap_8 FILLER_37_80 ();
 sg13g2_decap_8 FILLER_37_87 ();
 sg13g2_fill_2 FILLER_37_94 ();
 sg13g2_decap_4 FILLER_37_134 ();
 sg13g2_fill_1 FILLER_37_138 ();
 sg13g2_decap_8 FILLER_37_187 ();
 sg13g2_decap_8 FILLER_37_194 ();
 sg13g2_decap_4 FILLER_37_201 ();
 sg13g2_fill_2 FILLER_37_218 ();
 sg13g2_fill_1 FILLER_37_220 ();
 sg13g2_decap_4 FILLER_37_263 ();
 sg13g2_fill_1 FILLER_37_267 ();
 sg13g2_decap_4 FILLER_37_276 ();
 sg13g2_fill_1 FILLER_37_280 ();
 sg13g2_decap_8 FILLER_37_331 ();
 sg13g2_decap_4 FILLER_37_342 ();
 sg13g2_fill_1 FILLER_37_355 ();
 sg13g2_fill_2 FILLER_37_412 ();
 sg13g2_fill_1 FILLER_37_431 ();
 sg13g2_fill_2 FILLER_37_437 ();
 sg13g2_fill_1 FILLER_37_439 ();
 sg13g2_fill_2 FILLER_37_457 ();
 sg13g2_fill_2 FILLER_38_0 ();
 sg13g2_fill_1 FILLER_38_2 ();
 sg13g2_decap_4 FILLER_38_62 ();
 sg13g2_fill_1 FILLER_38_66 ();
 sg13g2_decap_8 FILLER_38_98 ();
 sg13g2_decap_8 FILLER_38_105 ();
 sg13g2_fill_2 FILLER_38_112 ();
 sg13g2_fill_1 FILLER_38_140 ();
 sg13g2_fill_1 FILLER_38_179 ();
 sg13g2_fill_2 FILLER_38_197 ();
 sg13g2_fill_1 FILLER_38_199 ();
 sg13g2_decap_8 FILLER_38_244 ();
 sg13g2_decap_8 FILLER_38_251 ();
 sg13g2_fill_2 FILLER_38_258 ();
 sg13g2_fill_2 FILLER_38_268 ();
 sg13g2_fill_1 FILLER_38_270 ();
 sg13g2_fill_2 FILLER_38_307 ();
 sg13g2_fill_1 FILLER_38_309 ();
 sg13g2_fill_2 FILLER_38_337 ();
 sg13g2_fill_1 FILLER_38_408 ();
 sg13g2_fill_2 FILLER_38_434 ();
 sg13g2_fill_2 FILLER_38_453 ();
 sg13g2_fill_2 FILLER_39_21 ();
 sg13g2_fill_1 FILLER_39_23 ();
 sg13g2_fill_2 FILLER_39_29 ();
 sg13g2_decap_4 FILLER_39_96 ();
 sg13g2_fill_1 FILLER_39_100 ();
 sg13g2_decap_4 FILLER_39_118 ();
 sg13g2_fill_1 FILLER_39_122 ();
 sg13g2_decap_4 FILLER_39_126 ();
 sg13g2_fill_1 FILLER_39_130 ();
 sg13g2_decap_4 FILLER_39_154 ();
 sg13g2_decap_8 FILLER_39_184 ();
 sg13g2_fill_2 FILLER_39_191 ();
 sg13g2_decap_4 FILLER_39_233 ();
 sg13g2_fill_1 FILLER_39_237 ();
 sg13g2_fill_2 FILLER_39_255 ();
 sg13g2_decap_8 FILLER_39_274 ();
 sg13g2_decap_8 FILLER_39_281 ();
 sg13g2_fill_2 FILLER_39_288 ();
 sg13g2_decap_4 FILLER_39_304 ();
 sg13g2_fill_2 FILLER_39_352 ();
 sg13g2_fill_1 FILLER_39_401 ();
 sg13g2_fill_2 FILLER_39_452 ();
 sg13g2_fill_1 FILLER_39_454 ();
 sg13g2_fill_2 FILLER_40_0 ();
 sg13g2_fill_1 FILLER_40_2 ();
 sg13g2_fill_2 FILLER_40_20 ();
 sg13g2_fill_2 FILLER_40_37 ();
 sg13g2_fill_1 FILLER_40_39 ();
 sg13g2_decap_8 FILLER_40_76 ();
 sg13g2_decap_8 FILLER_40_120 ();
 sg13g2_fill_2 FILLER_40_127 ();
 sg13g2_fill_1 FILLER_40_129 ();
 sg13g2_decap_8 FILLER_40_160 ();
 sg13g2_fill_1 FILLER_40_167 ();
 sg13g2_fill_2 FILLER_40_189 ();
 sg13g2_fill_1 FILLER_40_223 ();
 sg13g2_decap_8 FILLER_40_253 ();
 sg13g2_decap_8 FILLER_40_260 ();
 sg13g2_fill_1 FILLER_40_267 ();
 sg13g2_decap_8 FILLER_40_293 ();
 sg13g2_fill_2 FILLER_40_300 ();
 sg13g2_fill_1 FILLER_40_314 ();
 sg13g2_fill_2 FILLER_40_350 ();
 sg13g2_fill_2 FILLER_40_419 ();
 sg13g2_fill_1 FILLER_41_0 ();
 sg13g2_fill_1 FILLER_41_22 ();
 sg13g2_fill_1 FILLER_41_53 ();
 sg13g2_fill_1 FILLER_41_111 ();
 sg13g2_fill_2 FILLER_41_120 ();
 sg13g2_decap_8 FILLER_41_167 ();
 sg13g2_decap_4 FILLER_41_174 ();
 sg13g2_fill_2 FILLER_41_199 ();
 sg13g2_fill_2 FILLER_41_223 ();
 sg13g2_decap_8 FILLER_41_242 ();
 sg13g2_decap_4 FILLER_41_249 ();
 sg13g2_fill_1 FILLER_41_253 ();
 sg13g2_fill_1 FILLER_41_275 ();
 sg13g2_decap_4 FILLER_41_300 ();
 sg13g2_fill_2 FILLER_41_304 ();
 sg13g2_fill_1 FILLER_41_355 ();
 sg13g2_fill_1 FILLER_41_361 ();
 sg13g2_fill_2 FILLER_41_367 ();
 sg13g2_fill_1 FILLER_41_369 ();
 sg13g2_fill_1 FILLER_41_381 ();
 sg13g2_fill_2 FILLER_41_448 ();
 sg13g2_fill_1 FILLER_41_450 ();
 sg13g2_fill_2 FILLER_42_0 ();
 sg13g2_fill_2 FILLER_42_19 ();
 sg13g2_fill_1 FILLER_42_21 ();
 sg13g2_fill_2 FILLER_42_38 ();
 sg13g2_fill_1 FILLER_42_63 ();
 sg13g2_fill_1 FILLER_42_131 ();
 sg13g2_fill_2 FILLER_42_136 ();
 sg13g2_fill_1 FILLER_42_160 ();
 sg13g2_decap_4 FILLER_42_202 ();
 sg13g2_decap_8 FILLER_42_244 ();
 sg13g2_decap_8 FILLER_42_276 ();
 sg13g2_fill_2 FILLER_42_283 ();
 sg13g2_fill_2 FILLER_42_297 ();
 sg13g2_fill_2 FILLER_42_311 ();
 sg13g2_fill_1 FILLER_42_418 ();
 sg13g2_fill_1 FILLER_42_429 ();
 sg13g2_fill_2 FILLER_43_0 ();
 sg13g2_fill_2 FILLER_43_21 ();
 sg13g2_fill_1 FILLER_43_23 ();
 sg13g2_fill_2 FILLER_43_114 ();
 sg13g2_fill_1 FILLER_43_116 ();
 sg13g2_fill_2 FILLER_43_123 ();
 sg13g2_fill_1 FILLER_43_125 ();
 sg13g2_decap_4 FILLER_43_143 ();
 sg13g2_decap_4 FILLER_43_154 ();
 sg13g2_fill_2 FILLER_43_158 ();
 sg13g2_fill_2 FILLER_43_181 ();
 sg13g2_fill_2 FILLER_43_188 ();
 sg13g2_fill_1 FILLER_43_190 ();
 sg13g2_fill_2 FILLER_43_223 ();
 sg13g2_fill_2 FILLER_43_259 ();
 sg13g2_decap_4 FILLER_43_285 ();
 sg13g2_fill_1 FILLER_43_289 ();
 sg13g2_fill_1 FILLER_43_322 ();
 sg13g2_fill_2 FILLER_43_327 ();
 sg13g2_fill_2 FILLER_43_337 ();
 sg13g2_fill_2 FILLER_43_351 ();
 sg13g2_fill_1 FILLER_43_357 ();
 sg13g2_fill_2 FILLER_43_370 ();
 sg13g2_fill_1 FILLER_43_372 ();
 sg13g2_fill_2 FILLER_43_395 ();
 sg13g2_fill_1 FILLER_43_397 ();
 sg13g2_fill_1 FILLER_43_429 ();
 sg13g2_fill_2 FILLER_44_0 ();
 sg13g2_fill_2 FILLER_44_47 ();
 sg13g2_fill_1 FILLER_44_49 ();
 sg13g2_fill_2 FILLER_44_90 ();
 sg13g2_decap_4 FILLER_44_139 ();
 sg13g2_fill_1 FILLER_44_143 ();
 sg13g2_fill_1 FILLER_44_205 ();
 sg13g2_fill_2 FILLER_44_217 ();
 sg13g2_fill_1 FILLER_44_219 ();
 sg13g2_fill_1 FILLER_44_237 ();
 sg13g2_fill_1 FILLER_44_255 ();
 sg13g2_fill_1 FILLER_44_278 ();
 sg13g2_fill_2 FILLER_44_368 ();
 sg13g2_fill_1 FILLER_44_374 ();
 sg13g2_fill_1 FILLER_44_388 ();
 sg13g2_fill_2 FILLER_44_406 ();
 sg13g2_fill_2 FILLER_44_452 ();
 sg13g2_fill_1 FILLER_44_454 ();
 sg13g2_fill_2 FILLER_45_0 ();
 sg13g2_fill_2 FILLER_45_39 ();
 sg13g2_fill_1 FILLER_45_41 ();
 sg13g2_fill_2 FILLER_45_50 ();
 sg13g2_fill_1 FILLER_45_52 ();
 sg13g2_fill_2 FILLER_45_62 ();
 sg13g2_fill_1 FILLER_45_64 ();
 sg13g2_fill_1 FILLER_45_80 ();
 sg13g2_fill_1 FILLER_45_99 ();
 sg13g2_decap_4 FILLER_45_163 ();
 sg13g2_fill_1 FILLER_45_167 ();
 sg13g2_decap_4 FILLER_45_185 ();
 sg13g2_fill_1 FILLER_45_219 ();
 sg13g2_fill_1 FILLER_45_237 ();
 sg13g2_fill_1 FILLER_45_283 ();
 sg13g2_fill_2 FILLER_45_402 ();
 sg13g2_fill_1 FILLER_45_404 ();
 sg13g2_fill_1 FILLER_45_458 ();
 sg13g2_fill_2 FILLER_46_0 ();
 sg13g2_fill_2 FILLER_46_19 ();
 sg13g2_fill_2 FILLER_46_49 ();
 sg13g2_fill_1 FILLER_46_51 ();
 sg13g2_fill_2 FILLER_46_99 ();
 sg13g2_fill_1 FILLER_46_101 ();
 sg13g2_fill_2 FILLER_46_113 ();
 sg13g2_fill_1 FILLER_46_143 ();
 sg13g2_fill_2 FILLER_46_165 ();
 sg13g2_fill_1 FILLER_46_167 ();
 sg13g2_decap_8 FILLER_46_193 ();
 sg13g2_fill_2 FILLER_46_200 ();
 sg13g2_decap_8 FILLER_46_221 ();
 sg13g2_fill_2 FILLER_46_245 ();
 sg13g2_fill_1 FILLER_46_247 ();
 sg13g2_fill_2 FILLER_46_346 ();
 sg13g2_fill_1 FILLER_46_348 ();
 sg13g2_fill_2 FILLER_46_407 ();
 sg13g2_fill_1 FILLER_47_0 ();
 sg13g2_fill_2 FILLER_47_56 ();
 sg13g2_fill_1 FILLER_47_58 ();
 sg13g2_fill_2 FILLER_47_162 ();
 sg13g2_fill_1 FILLER_47_185 ();
 sg13g2_decap_4 FILLER_47_226 ();
 sg13g2_fill_1 FILLER_47_280 ();
 sg13g2_fill_1 FILLER_47_289 ();
 sg13g2_fill_2 FILLER_47_302 ();
 sg13g2_fill_1 FILLER_47_304 ();
 sg13g2_fill_1 FILLER_47_327 ();
 sg13g2_fill_2 FILLER_47_399 ();
 sg13g2_fill_1 FILLER_47_401 ();
 sg13g2_fill_1 FILLER_47_432 ();
 sg13g2_fill_1 FILLER_47_458 ();
 sg13g2_fill_2 FILLER_48_82 ();
 sg13g2_fill_2 FILLER_48_133 ();
 sg13g2_fill_1 FILLER_48_135 ();
 sg13g2_decap_8 FILLER_48_186 ();
 sg13g2_fill_2 FILLER_48_193 ();
 sg13g2_fill_2 FILLER_48_223 ();
 sg13g2_fill_2 FILLER_48_268 ();
 sg13g2_fill_1 FILLER_48_330 ();
 sg13g2_fill_2 FILLER_48_352 ();
 sg13g2_fill_1 FILLER_48_354 ();
 sg13g2_fill_2 FILLER_48_380 ();
 sg13g2_fill_2 FILLER_48_396 ();
 sg13g2_fill_1 FILLER_48_398 ();
 sg13g2_fill_2 FILLER_49_0 ();
 sg13g2_fill_1 FILLER_49_19 ();
 sg13g2_fill_1 FILLER_49_43 ();
 sg13g2_fill_2 FILLER_49_49 ();
 sg13g2_fill_1 FILLER_49_51 ();
 sg13g2_fill_2 FILLER_49_79 ();
 sg13g2_fill_2 FILLER_49_158 ();
 sg13g2_fill_2 FILLER_49_193 ();
 sg13g2_fill_1 FILLER_49_221 ();
 sg13g2_fill_2 FILLER_49_247 ();
 sg13g2_fill_1 FILLER_49_249 ();
 sg13g2_fill_2 FILLER_49_271 ();
 sg13g2_fill_1 FILLER_49_273 ();
 sg13g2_fill_1 FILLER_49_387 ();
 sg13g2_fill_2 FILLER_49_417 ();
 sg13g2_fill_2 FILLER_49_457 ();
 sg13g2_fill_2 FILLER_50_0 ();
 sg13g2_fill_1 FILLER_50_2 ();
 sg13g2_fill_1 FILLER_50_24 ();
 sg13g2_fill_2 FILLER_50_35 ();
 sg13g2_fill_2 FILLER_50_96 ();
 sg13g2_fill_1 FILLER_50_98 ();
 sg13g2_fill_2 FILLER_50_149 ();
 sg13g2_fill_2 FILLER_50_168 ();
 sg13g2_fill_2 FILLER_50_188 ();
 sg13g2_fill_1 FILLER_50_211 ();
 sg13g2_fill_2 FILLER_50_222 ();
 sg13g2_fill_1 FILLER_50_234 ();
 sg13g2_fill_1 FILLER_50_272 ();
 sg13g2_fill_2 FILLER_50_307 ();
 sg13g2_fill_2 FILLER_50_407 ();
 sg13g2_fill_1 FILLER_50_409 ();
 sg13g2_fill_2 FILLER_50_418 ();
 sg13g2_fill_1 FILLER_50_420 ();
 sg13g2_fill_2 FILLER_51_0 ();
 sg13g2_fill_2 FILLER_51_19 ();
 sg13g2_fill_1 FILLER_51_21 ();
 sg13g2_fill_2 FILLER_51_47 ();
 sg13g2_fill_2 FILLER_51_75 ();
 sg13g2_fill_1 FILLER_51_77 ();
 sg13g2_fill_2 FILLER_51_103 ();
 sg13g2_fill_1 FILLER_51_105 ();
 sg13g2_fill_2 FILLER_51_136 ();
 sg13g2_fill_1 FILLER_51_138 ();
 sg13g2_fill_2 FILLER_51_144 ();
 sg13g2_fill_1 FILLER_51_146 ();
 sg13g2_fill_2 FILLER_51_164 ();
 sg13g2_fill_1 FILLER_51_166 ();
 sg13g2_fill_2 FILLER_51_209 ();
 sg13g2_fill_2 FILLER_51_258 ();
 sg13g2_fill_2 FILLER_51_276 ();
 sg13g2_fill_2 FILLER_51_302 ();
 sg13g2_fill_1 FILLER_51_304 ();
 sg13g2_fill_2 FILLER_51_327 ();
 sg13g2_fill_1 FILLER_51_329 ();
 sg13g2_fill_2 FILLER_51_432 ();
 sg13g2_fill_1 FILLER_51_434 ();
 sg13g2_fill_2 FILLER_51_456 ();
 sg13g2_fill_1 FILLER_51_458 ();
 sg13g2_fill_2 FILLER_52_0 ();
 sg13g2_fill_1 FILLER_52_2 ();
 sg13g2_fill_2 FILLER_52_41 ();
 sg13g2_fill_1 FILLER_52_43 ();
 sg13g2_fill_1 FILLER_52_82 ();
 sg13g2_fill_1 FILLER_52_119 ();
 sg13g2_fill_2 FILLER_52_179 ();
 sg13g2_fill_2 FILLER_52_249 ();
 sg13g2_fill_1 FILLER_52_251 ();
 sg13g2_fill_2 FILLER_52_294 ();
 sg13g2_fill_1 FILLER_52_296 ();
 sg13g2_fill_2 FILLER_52_321 ();
 sg13g2_fill_1 FILLER_52_369 ();
 sg13g2_fill_2 FILLER_52_388 ();
 sg13g2_fill_2 FILLER_52_415 ();
 sg13g2_fill_2 FILLER_52_434 ();
 sg13g2_fill_2 FILLER_52_457 ();
 sg13g2_fill_2 FILLER_53_0 ();
 sg13g2_fill_2 FILLER_53_19 ();
 sg13g2_fill_1 FILLER_53_36 ();
 sg13g2_fill_2 FILLER_53_71 ();
 sg13g2_fill_1 FILLER_53_73 ();
 sg13g2_fill_2 FILLER_53_101 ();
 sg13g2_fill_2 FILLER_53_130 ();
 sg13g2_fill_2 FILLER_53_137 ();
 sg13g2_fill_2 FILLER_53_178 ();
 sg13g2_fill_1 FILLER_53_180 ();
 sg13g2_fill_2 FILLER_53_191 ();
 sg13g2_fill_1 FILLER_53_193 ();
 sg13g2_fill_2 FILLER_53_258 ();
 sg13g2_fill_1 FILLER_53_260 ();
 sg13g2_fill_2 FILLER_53_303 ();
 sg13g2_fill_1 FILLER_53_305 ();
 sg13g2_fill_2 FILLER_53_340 ();
 sg13g2_fill_1 FILLER_53_342 ();
 sg13g2_fill_2 FILLER_53_350 ();
 sg13g2_fill_1 FILLER_53_382 ();
 sg13g2_fill_1 FILLER_53_417 ();
 sg13g2_fill_2 FILLER_54_0 ();
 sg13g2_fill_2 FILLER_54_44 ();
 sg13g2_fill_2 FILLER_54_128 ();
 sg13g2_fill_1 FILLER_54_148 ();
 sg13g2_fill_2 FILLER_54_159 ();
 sg13g2_fill_1 FILLER_54_167 ();
 sg13g2_fill_1 FILLER_54_200 ();
 sg13g2_fill_2 FILLER_54_209 ();
 sg13g2_fill_1 FILLER_54_211 ();
 sg13g2_fill_2 FILLER_54_237 ();
 sg13g2_fill_1 FILLER_54_251 ();
 sg13g2_fill_2 FILLER_54_273 ();
 sg13g2_fill_1 FILLER_54_275 ();
 sg13g2_fill_1 FILLER_54_305 ();
 sg13g2_fill_1 FILLER_54_327 ();
 sg13g2_fill_2 FILLER_54_375 ();
 sg13g2_fill_1 FILLER_54_377 ();
 sg13g2_fill_1 FILLER_54_412 ();
 sg13g2_fill_1 FILLER_54_458 ();
 sg13g2_fill_2 FILLER_55_0 ();
 sg13g2_fill_2 FILLER_55_31 ();
 sg13g2_fill_1 FILLER_55_33 ();
 sg13g2_fill_2 FILLER_55_111 ();
 sg13g2_fill_2 FILLER_55_164 ();
 sg13g2_fill_1 FILLER_55_166 ();
 sg13g2_fill_1 FILLER_55_207 ();
 sg13g2_fill_2 FILLER_55_237 ();
 sg13g2_fill_1 FILLER_55_239 ();
 sg13g2_fill_2 FILLER_55_244 ();
 sg13g2_fill_1 FILLER_55_246 ();
 sg13g2_fill_2 FILLER_55_281 ();
 sg13g2_fill_1 FILLER_55_283 ();
 sg13g2_fill_2 FILLER_55_301 ();
 sg13g2_fill_1 FILLER_55_303 ();
 sg13g2_fill_1 FILLER_55_325 ();
 sg13g2_fill_1 FILLER_55_352 ();
 sg13g2_fill_2 FILLER_55_367 ();
 sg13g2_fill_1 FILLER_55_376 ();
 sg13g2_fill_1 FILLER_55_403 ();
 sg13g2_fill_2 FILLER_55_421 ();
 sg13g2_fill_2 FILLER_56_0 ();
 sg13g2_fill_2 FILLER_56_41 ();
 sg13g2_fill_1 FILLER_56_43 ();
 sg13g2_fill_2 FILLER_56_59 ();
 sg13g2_fill_2 FILLER_56_87 ();
 sg13g2_fill_1 FILLER_56_104 ();
 sg13g2_fill_2 FILLER_56_120 ();
 sg13g2_fill_2 FILLER_56_126 ();
 sg13g2_fill_2 FILLER_56_159 ();
 sg13g2_fill_2 FILLER_56_198 ();
 sg13g2_fill_1 FILLER_56_200 ();
 sg13g2_fill_2 FILLER_56_222 ();
 sg13g2_fill_1 FILLER_56_278 ();
 sg13g2_fill_2 FILLER_56_287 ();
 sg13g2_fill_2 FILLER_56_297 ();
 sg13g2_fill_1 FILLER_56_299 ();
 sg13g2_fill_2 FILLER_56_333 ();
 sg13g2_fill_1 FILLER_56_335 ();
 sg13g2_fill_1 FILLER_56_371 ();
 sg13g2_fill_1 FILLER_56_435 ();
 sg13g2_fill_1 FILLER_56_454 ();
 sg13g2_fill_2 FILLER_57_0 ();
 sg13g2_fill_2 FILLER_57_10 ();
 sg13g2_fill_1 FILLER_57_12 ();
 sg13g2_fill_2 FILLER_57_67 ();
 sg13g2_fill_1 FILLER_57_69 ();
 sg13g2_fill_2 FILLER_57_87 ();
 sg13g2_fill_1 FILLER_57_140 ();
 sg13g2_fill_2 FILLER_57_158 ();
 sg13g2_fill_2 FILLER_57_214 ();
 sg13g2_fill_1 FILLER_57_216 ();
 sg13g2_fill_2 FILLER_57_262 ();
 sg13g2_fill_1 FILLER_57_338 ();
 sg13g2_fill_1 FILLER_57_377 ();
 sg13g2_fill_2 FILLER_57_407 ();
 sg13g2_fill_1 FILLER_57_409 ();
 sg13g2_fill_2 FILLER_58_0 ();
 sg13g2_fill_1 FILLER_58_2 ();
 sg13g2_fill_2 FILLER_58_36 ();
 sg13g2_fill_1 FILLER_58_38 ();
 sg13g2_fill_1 FILLER_58_64 ();
 sg13g2_fill_2 FILLER_58_121 ();
 sg13g2_fill_2 FILLER_58_284 ();
 sg13g2_fill_1 FILLER_58_324 ();
 sg13g2_fill_2 FILLER_58_379 ();
 sg13g2_fill_1 FILLER_58_381 ();
 sg13g2_fill_2 FILLER_59_0 ();
 sg13g2_fill_1 FILLER_59_2 ();
 sg13g2_fill_2 FILLER_59_28 ();
 sg13g2_fill_1 FILLER_59_30 ();
 sg13g2_fill_1 FILLER_59_69 ();
 sg13g2_fill_2 FILLER_59_87 ();
 sg13g2_fill_2 FILLER_59_108 ();
 sg13g2_fill_1 FILLER_59_110 ();
 sg13g2_fill_2 FILLER_59_140 ();
 sg13g2_fill_1 FILLER_59_150 ();
 sg13g2_fill_2 FILLER_59_196 ();
 sg13g2_fill_1 FILLER_59_198 ();
 sg13g2_fill_2 FILLER_59_239 ();
 sg13g2_fill_2 FILLER_59_289 ();
 sg13g2_fill_1 FILLER_59_291 ();
 sg13g2_fill_2 FILLER_59_317 ();
 sg13g2_fill_1 FILLER_59_319 ();
 sg13g2_fill_1 FILLER_59_357 ();
 sg13g2_fill_2 FILLER_59_379 ();
 sg13g2_fill_1 FILLER_59_381 ();
endmodule
