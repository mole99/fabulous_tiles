* NGSPICE file created from N_term_single.ext - technology: ihp-sg13g2

* Black-box entry subcircuit for sg13g2_decap_8 abstract view
.subckt sg13g2_decap_8 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_1 abstract view
.subckt sg13g2_fill_1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_decap_4 abstract view
.subckt sg13g2_decap_4 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_2 abstract view
.subckt sg13g2_fill_2 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_1 abstract view
.subckt sg13g2_buf_1 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_antennanp abstract view
.subckt sg13g2_antennanp VDD VSS A
.ends

.subckt N_term_single Ci FrameData[0] FrameData[10] FrameData[11] FrameData[12] FrameData[13]
+ FrameData[14] FrameData[15] FrameData[16] FrameData[17] FrameData[18] FrameData[19]
+ FrameData[1] FrameData[20] FrameData[21] FrameData[22] FrameData[23] FrameData[24]
+ FrameData[25] FrameData[26] FrameData[27] FrameData[28] FrameData[29] FrameData[2]
+ FrameData[30] FrameData[31] FrameData[3] FrameData[4] FrameData[5] FrameData[6]
+ FrameData[7] FrameData[8] FrameData[9] FrameData_O[0] FrameData_O[10] FrameData_O[11]
+ FrameData_O[12] FrameData_O[13] FrameData_O[14] FrameData_O[15] FrameData_O[16]
+ FrameData_O[17] FrameData_O[18] FrameData_O[19] FrameData_O[1] FrameData_O[20] FrameData_O[21]
+ FrameData_O[22] FrameData_O[23] FrameData_O[24] FrameData_O[25] FrameData_O[26]
+ FrameData_O[27] FrameData_O[28] FrameData_O[29] FrameData_O[2] FrameData_O[30] FrameData_O[31]
+ FrameData_O[3] FrameData_O[4] FrameData_O[5] FrameData_O[6] FrameData_O[7] FrameData_O[8]
+ FrameData_O[9] FrameStrobe[0] FrameStrobe[10] FrameStrobe[11] FrameStrobe[12] FrameStrobe[13]
+ FrameStrobe[14] FrameStrobe[15] FrameStrobe[16] FrameStrobe[17] FrameStrobe[18]
+ FrameStrobe[19] FrameStrobe[1] FrameStrobe[2] FrameStrobe[3] FrameStrobe[4] FrameStrobe[5]
+ FrameStrobe[6] FrameStrobe[7] FrameStrobe[8] FrameStrobe[9] FrameStrobe_O[0] FrameStrobe_O[10]
+ FrameStrobe_O[11] FrameStrobe_O[12] FrameStrobe_O[13] FrameStrobe_O[14] FrameStrobe_O[15]
+ FrameStrobe_O[16] FrameStrobe_O[17] FrameStrobe_O[18] FrameStrobe_O[19] FrameStrobe_O[1]
+ FrameStrobe_O[2] FrameStrobe_O[3] FrameStrobe_O[4] FrameStrobe_O[5] FrameStrobe_O[6]
+ FrameStrobe_O[7] FrameStrobe_O[8] FrameStrobe_O[9] N1END[0] N1END[1] N1END[2] N1END[3]
+ N2END[0] N2END[1] N2END[2] N2END[3] N2END[4] N2END[5] N2END[6] N2END[7] N2MID[0]
+ N2MID[1] N2MID[2] N2MID[3] N2MID[4] N2MID[5] N2MID[6] N2MID[7] N4END[0] N4END[10]
+ N4END[11] N4END[12] N4END[13] N4END[14] N4END[15] N4END[1] N4END[2] N4END[3] N4END[4]
+ N4END[5] N4END[6] N4END[7] N4END[8] N4END[9] NN4END[0] NN4END[10] NN4END[11] NN4END[12]
+ NN4END[13] NN4END[14] NN4END[15] NN4END[1] NN4END[2] NN4END[3] NN4END[4] NN4END[5]
+ NN4END[6] NN4END[7] NN4END[8] NN4END[9] S1BEG[0] S1BEG[1] S1BEG[2] S1BEG[3] S2BEG[0]
+ S2BEG[1] S2BEG[2] S2BEG[3] S2BEG[4] S2BEG[5] S2BEG[6] S2BEG[7] S2BEGb[0] S2BEGb[1]
+ S2BEGb[2] S2BEGb[3] S2BEGb[4] S2BEGb[5] S2BEGb[6] S2BEGb[7] S4BEG[0] S4BEG[10] S4BEG[11]
+ S4BEG[12] S4BEG[13] S4BEG[14] S4BEG[15] S4BEG[1] S4BEG[2] S4BEG[3] S4BEG[4] S4BEG[5]
+ S4BEG[6] S4BEG[7] S4BEG[8] S4BEG[9] SS4BEG[0] SS4BEG[10] SS4BEG[11] SS4BEG[12] SS4BEG[13]
+ SS4BEG[14] SS4BEG[15] SS4BEG[1] SS4BEG[2] SS4BEG[3] SS4BEG[4] SS4BEG[5] SS4BEG[6]
+ SS4BEG[7] SS4BEG[8] SS4BEG[9] UserCLK UserCLKo VGND VPWR
XFILLER_7_7 VPWR VGND sg13g2_decap_8
XFILLER_5_376 VPWR VGND sg13g2_fill_1
XFILLER_5_354 VPWR VGND sg13g2_decap_8
XFILLER_3_56 VPWR VGND sg13g2_decap_4
XFILLER_10_147 VPWR VGND sg13g2_decap_8
XFILLER_6_118 VPWR VGND sg13g2_decap_8
XFILLER_2_346 VPWR VGND sg13g2_decap_4
XFILLER_2_379 VPWR VGND sg13g2_fill_2
XFILLER_5_195 VPWR VGND sg13g2_decap_8
XFILLER_11_423 VPWR VGND sg13g2_decap_4
XFILLER_11_401 VPWR VGND sg13g2_decap_4
X_062_ N2MID[1] net63 VPWR VGND sg13g2_buf_1
XFILLER_9_88 VPWR VGND sg13g2_decap_8
XFILLER_0_35 VPWR VGND sg13g2_decap_8
XFILLER_2_154 VPWR VGND sg13g2_decap_8
XFILLER_4_408 VPWR VGND sg13g2_fill_1
X_045_ FrameStrobe[13] net37 VPWR VGND sg13g2_buf_1
XFILLER_7_268 VPWR VGND sg13g2_decap_8
XFILLER_0_433 VPWR VGND sg13g2_decap_8
XFILLER_4_249 VPWR VGND sg13g2_decap_8
X_028_ FrameData[28] net21 VPWR VGND sg13g2_buf_1
XFILLER_6_56 VPWR VGND sg13g2_decap_8
XANTENNA_5 VPWR VGND FrameData[5] sg13g2_antennanp
XFILLER_3_271 VPWR VGND sg13g2_decap_4
XFILLER_3_293 VPWR VGND sg13g2_decap_8
Xoutput20 net20 FrameData_O[27] VPWR VGND sg13g2_buf_1
Xoutput42 net42 FrameStrobe_O[18] VPWR VGND sg13g2_buf_1
XFILLER_8_352 VPWR VGND sg13g2_decap_8
Xoutput7 net7 FrameData_O[15] VPWR VGND sg13g2_buf_1
Xoutput75 net75 S4BEG[11] VPWR VGND sg13g2_buf_1
Xoutput86 net86 S4BEG[7] VPWR VGND sg13g2_buf_1
Xoutput64 net64 S2BEG[7] VPWR VGND sg13g2_buf_1
Xoutput53 net53 S1BEG[0] VPWR VGND sg13g2_buf_1
Xoutput97 net97 SS4BEG[2] VPWR VGND sg13g2_buf_1
Xoutput31 net31 FrameData_O[8] VPWR VGND sg13g2_buf_1
XFILLER_11_0 VPWR VGND sg13g2_decap_8
XFILLER_10_329 VPWR VGND sg13g2_decap_8
XFILLER_9_149 VPWR VGND sg13g2_decap_8
XFILLER_9_116 VPWR VGND sg13g2_decap_8
XFILLER_5_399 VPWR VGND sg13g2_decap_8
XFILLER_3_35 VPWR VGND sg13g2_decap_8
XFILLER_3_79 VPWR VGND sg13g2_decap_8
XFILLER_10_126 VPWR VGND sg13g2_decap_8
XFILLER_2_325 VPWR VGND sg13g2_decap_8
XFILLER_5_174 VPWR VGND sg13g2_decap_8
XFILLER_1_391 VPWR VGND sg13g2_decap_8
XFILLER_11_435 VPWR VGND sg13g2_fill_2
XFILLER_9_56 VPWR VGND sg13g2_fill_1
X_061_ N2MID[2] net62 VPWR VGND sg13g2_buf_1
XFILLER_0_14 VPWR VGND sg13g2_decap_8
XFILLER_2_133 VPWR VGND sg13g2_decap_8
X_044_ FrameStrobe[12] net36 VPWR VGND sg13g2_buf_1
XFILLER_7_247 VPWR VGND sg13g2_decap_8
XFILLER_6_291 VPWR VGND sg13g2_decap_8
XFILLER_0_412 VPWR VGND sg13g2_decap_8
X_027_ FrameData[27] net20 VPWR VGND sg13g2_buf_1
XFILLER_6_35 VPWR VGND sg13g2_decap_8
XFILLER_3_250 VPWR VGND sg13g2_fill_1
XANTENNA_6 VPWR VGND FrameData[5] sg13g2_antennanp
Xoutput43 net43 FrameStrobe_O[19] VPWR VGND sg13g2_buf_1
Xoutput21 net21 FrameData_O[28] VPWR VGND sg13g2_buf_1
XFILLER_9_309 VPWR VGND sg13g2_decap_4
Xoutput10 net10 FrameData_O[18] VPWR VGND sg13g2_buf_1
Xoutput8 net8 FrameData_O[16] VPWR VGND sg13g2_buf_1
Xoutput87 net87 S4BEG[8] VPWR VGND sg13g2_buf_1
Xoutput65 net65 S2BEGb[0] VPWR VGND sg13g2_buf_1
Xoutput54 net54 S1BEG[1] VPWR VGND sg13g2_buf_1
Xoutput76 net76 S4BEG[12] VPWR VGND sg13g2_buf_1
Xoutput98 net98 SS4BEG[3] VPWR VGND sg13g2_buf_1
Xoutput32 net32 FrameData_O[9] VPWR VGND sg13g2_buf_1
XFILLER_10_308 VPWR VGND sg13g2_decap_8
XFILLER_8_331 VPWR VGND sg13g2_decap_8
XFILLER_9_128 VPWR VGND sg13g2_decap_8
XFILLER_5_323 VPWR VGND sg13g2_decap_8
XFILLER_8_194 VPWR VGND sg13g2_decap_8
XFILLER_3_14 VPWR VGND sg13g2_decap_8
XFILLER_10_105 VPWR VGND sg13g2_decap_8
XFILLER_2_304 VPWR VGND sg13g2_fill_2
XFILLER_5_153 VPWR VGND sg13g2_decap_8
XFILLER_1_370 VPWR VGND sg13g2_decap_8
XFILLER_9_35 VPWR VGND sg13g2_decap_8
XFILLER_7_429 VPWR VGND sg13g2_decap_8
X_060_ N2MID[3] net61 VPWR VGND sg13g2_buf_1
XFILLER_2_112 VPWR VGND sg13g2_decap_8
XFILLER_2_189 VPWR VGND sg13g2_decap_8
XFILLER_11_299 VPWR VGND sg13g2_decap_8
XFILLER_11_277 VPWR VGND sg13g2_decap_8
XFILLER_11_255 VPWR VGND sg13g2_decap_8
XFILLER_11_233 VPWR VGND sg13g2_decap_8
XFILLER_11_211 VPWR VGND sg13g2_decap_8
X_043_ FrameStrobe[11] net35 VPWR VGND sg13g2_buf_1
XFILLER_7_226 VPWR VGND sg13g2_decap_8
XFILLER_1_0 VPWR VGND sg13g2_decap_8
XFILLER_3_443 VPWR VGND sg13g2_decap_4
XFILLER_1_91 VPWR VGND sg13g2_decap_8
X_026_ FrameData[26] net19 VPWR VGND sg13g2_buf_1
XFILLER_6_14 VPWR VGND sg13g2_decap_8
XANTENNA_7 VPWR VGND FrameData[6] sg13g2_antennanp
Xoutput44 net44 FrameStrobe_O[1] VPWR VGND sg13g2_buf_1
Xoutput33 net33 FrameStrobe_O[0] VPWR VGND sg13g2_buf_1
Xoutput22 net22 FrameData_O[29] VPWR VGND sg13g2_buf_1
Xoutput11 net11 FrameData_O[19] VPWR VGND sg13g2_buf_1
Xoutput9 net9 FrameData_O[17] VPWR VGND sg13g2_buf_1
Xoutput77 net77 S4BEG[13] VPWR VGND sg13g2_buf_1
Xoutput88 net88 S4BEG[9] VPWR VGND sg13g2_buf_1
Xoutput66 net66 S2BEGb[1] VPWR VGND sg13g2_buf_1
Xoutput55 net55 S1BEG[2] VPWR VGND sg13g2_buf_1
Xoutput99 net99 SS4BEG[4] VPWR VGND sg13g2_buf_1
XFILLER_8_387 VPWR VGND sg13g2_decap_8
XFILLER_8_310 VPWR VGND sg13g2_decap_8
X_009_ FrameData[9] net32 VPWR VGND sg13g2_buf_1
XFILLER_8_140 VPWR VGND sg13g2_decap_8
XFILLER_5_368 VPWR VGND sg13g2_decap_4
XFILLER_5_302 VPWR VGND sg13g2_decap_8
XFILLER_5_7 VPWR VGND sg13g2_decap_8
XFILLER_5_132 VPWR VGND sg13g2_decap_8
XFILLER_7_408 VPWR VGND sg13g2_decap_8
XFILLER_0_49 VPWR VGND sg13g2_decap_8
XFILLER_2_168 VPWR VGND sg13g2_decap_8
XFILLER_9_69 VPWR VGND sg13g2_decap_8
XFILLER_9_14 VPWR VGND sg13g2_decap_8
XFILLER_9_290 VPWR VGND sg13g2_fill_1
X_042_ FrameStrobe[10] net34 VPWR VGND sg13g2_buf_1
XFILLER_3_400 VPWR VGND sg13g2_decap_4
XFILLER_6_260 VPWR VGND sg13g2_decap_8
XFILLER_1_70 VPWR VGND sg13g2_decap_8
X_025_ FrameData[25] net18 VPWR VGND sg13g2_buf_1
XFILLER_3_241 VPWR VGND sg13g2_fill_1
XANTENNA_8 VPWR VGND FrameData[6] sg13g2_antennanp
Xoutput34 net34 FrameStrobe_O[10] VPWR VGND sg13g2_buf_1
Xoutput45 net45 FrameStrobe_O[2] VPWR VGND sg13g2_buf_1
Xoutput67 net67 S2BEGb[2] VPWR VGND sg13g2_buf_1
Xoutput56 net56 S1BEG[3] VPWR VGND sg13g2_buf_1
Xoutput78 net78 S4BEG[14] VPWR VGND sg13g2_buf_1
Xoutput89 net89 SS4BEG[0] VPWR VGND sg13g2_buf_1
Xoutput12 net12 FrameData_O[1] VPWR VGND sg13g2_buf_1
Xoutput23 net23 FrameData_O[2] VPWR VGND sg13g2_buf_1
XFILLER_8_366 VPWR VGND sg13g2_decap_8
X_008_ FrameData[8] net31 VPWR VGND sg13g2_buf_1
XFILLER_7_91 VPWR VGND sg13g2_decap_8
XFILLER_5_347 VPWR VGND sg13g2_decap_8
XFILLER_3_49 VPWR VGND sg13g2_decap_8
XFILLER_5_111 VPWR VGND sg13g2_decap_4
XFILLER_2_306 VPWR VGND sg13g2_fill_1
XFILLER_2_339 VPWR VGND sg13g2_decap_8
XFILLER_5_188 VPWR VGND sg13g2_decap_8
XFILLER_11_416 VPWR VGND sg13g2_decap_8
XFILLER_2_147 VPWR VGND sg13g2_decap_8
XFILLER_4_70 VPWR VGND sg13g2_decap_4
XFILLER_4_92 VPWR VGND sg13g2_decap_8
XFILLER_6_442 VPWR VGND sg13g2_decap_8
XFILLER_0_28 VPWR VGND sg13g2_decap_8
X_041_ FrameStrobe[9] net52 VPWR VGND sg13g2_buf_1
XFILLER_0_426 VPWR VGND sg13g2_decap_8
X_024_ FrameData[24] net17 VPWR VGND sg13g2_buf_1
XFILLER_10_91 VPWR VGND sg13g2_decap_8
XFILLER_6_49 VPWR VGND sg13g2_decap_8
XANTENNA_9 VPWR VGND FrameData[8] sg13g2_antennanp
XFILLER_3_264 VPWR VGND sg13g2_decap_8
XFILLER_3_286 VPWR VGND sg13g2_decap_8
Xoutput24 net24 FrameData_O[30] VPWR VGND sg13g2_buf_1
Xoutput35 net35 FrameStrobe_O[11] VPWR VGND sg13g2_buf_1
Xoutput46 net46 FrameStrobe_O[3] VPWR VGND sg13g2_buf_1
Xoutput13 net13 FrameData_O[20] VPWR VGND sg13g2_buf_1
Xoutput57 net57 S2BEG[0] VPWR VGND sg13g2_buf_1
XFILLER_8_345 VPWR VGND sg13g2_decap_8
X_007_ FrameData[7] net30 VPWR VGND sg13g2_buf_1
Xoutput68 net68 S2BEGb[3] VPWR VGND sg13g2_buf_1
Xoutput79 net79 S4BEG[15] VPWR VGND sg13g2_buf_1
XFILLER_7_70 VPWR VGND sg13g2_decap_8
XFILLER_9_109 VPWR VGND sg13g2_decap_8
XFILLER_5_337 VPWR VGND sg13g2_decap_4
XFILLER_3_28 VPWR VGND sg13g2_decap_8
XFILLER_4_370 VPWR VGND sg13g2_decap_8
XFILLER_10_119 VPWR VGND sg13g2_decap_8
XFILLER_2_318 VPWR VGND sg13g2_decap_8
XFILLER_9_440 VPWR VGND sg13g2_decap_8
XFILLER_5_167 VPWR VGND sg13g2_decap_8
XFILLER_1_384 VPWR VGND sg13g2_decap_8
XFILLER_4_60 VPWR VGND sg13g2_fill_2
XFILLER_9_49 VPWR VGND sg13g2_fill_2
XFILLER_6_421 VPWR VGND sg13g2_decap_8
XFILLER_2_126 VPWR VGND sg13g2_decap_8
XFILLER_11_269 VPWR VGND sg13g2_decap_4
XFILLER_11_247 VPWR VGND sg13g2_decap_4
XFILLER_11_225 VPWR VGND sg13g2_decap_4
XFILLER_11_203 VPWR VGND sg13g2_decap_4
X_040_ FrameStrobe[8] net51 VPWR VGND sg13g2_buf_1
XFILLER_10_280 VPWR VGND sg13g2_decap_8
XFILLER_6_284 VPWR VGND sg13g2_decap_8
XFILLER_0_405 VPWR VGND sg13g2_decap_8
X_023_ FrameData[23] net16 VPWR VGND sg13g2_buf_1
XFILLER_10_70 VPWR VGND sg13g2_decap_8
XFILLER_6_28 VPWR VGND sg13g2_decap_8
Xoutput36 net36 FrameStrobe_O[12] VPWR VGND sg13g2_buf_1
Xoutput47 net47 FrameStrobe_O[4] VPWR VGND sg13g2_buf_1
Xoutput25 net25 FrameData_O[31] VPWR VGND sg13g2_buf_1
Xoutput14 net14 FrameData_O[21] VPWR VGND sg13g2_buf_1
XFILLER_8_324 VPWR VGND sg13g2_decap_8
X_006_ FrameData[6] net29 VPWR VGND sg13g2_buf_1
Xoutput69 net69 S2BEGb[4] VPWR VGND sg13g2_buf_1
Xoutput58 net58 S2BEG[1] VPWR VGND sg13g2_buf_1
XFILLER_5_316 VPWR VGND sg13g2_decap_8
XFILLER_8_187 VPWR VGND sg13g2_decap_8
XFILLER_8_176 VPWR VGND sg13g2_fill_2
XFILLER_8_154 VPWR VGND sg13g2_fill_2
XFILLER_5_146 VPWR VGND sg13g2_decap_8
XFILLER_1_363 VPWR VGND sg13g2_decap_8
XFILLER_4_190 VPWR VGND sg13g2_decap_8
XFILLER_9_28 VPWR VGND sg13g2_decap_8
XFILLER_6_400 VPWR VGND sg13g2_decap_8
XFILLER_2_105 VPWR VGND sg13g2_decap_8
XFILLER_3_7 VPWR VGND sg13g2_decap_8
XFILLER_1_182 VPWR VGND sg13g2_decap_8
XFILLER_7_219 VPWR VGND sg13g2_decap_8
XFILLER_3_436 VPWR VGND sg13g2_decap_8
XFILLER_6_274 VPWR VGND sg13g2_decap_4
X_099_ NN4END[4] net91 VPWR VGND sg13g2_buf_1
XFILLER_1_84 VPWR VGND sg13g2_decap_8
X_022_ FrameData[22] net15 VPWR VGND sg13g2_buf_1
XFILLER_3_233 VPWR VGND sg13g2_decap_4
XFILLER_3_255 VPWR VGND sg13g2_decap_4
Xoutput37 net37 FrameStrobe_O[13] VPWR VGND sg13g2_buf_1
Xoutput48 net48 FrameStrobe_O[5] VPWR VGND sg13g2_buf_1
Xoutput15 net15 FrameData_O[22] VPWR VGND sg13g2_buf_1
XFILLER_8_303 VPWR VGND sg13g2_decap_8
Xoutput59 net59 S2BEG[2] VPWR VGND sg13g2_buf_1
XFILLER_0_203 VPWR VGND sg13g2_fill_2
Xoutput26 net26 FrameData_O[3] VPWR VGND sg13g2_buf_1
X_005_ FrameData[5] net28 VPWR VGND sg13g2_buf_1
XFILLER_7_380 VPWR VGND sg13g2_decap_8
XFILLER_8_133 VPWR VGND sg13g2_decap_8
XFILLER_4_383 VPWR VGND sg13g2_decap_4
XFILLER_10_441 VPWR VGND sg13g2_fill_2
XFILLER_9_261 VPWR VGND sg13g2_decap_8
XFILLER_9_250 VPWR VGND sg13g2_decap_8
XFILLER_1_161 VPWR VGND sg13g2_decap_8
XFILLER_6_253 VPWR VGND sg13g2_decap_8
X_098_ NN4END[5] net90 VPWR VGND sg13g2_buf_1
XFILLER_1_63 VPWR VGND sg13g2_decap_8
X_021_ FrameData[21] net14 VPWR VGND sg13g2_buf_1
XFILLER_3_212 VPWR VGND sg13g2_decap_8
Xoutput38 net38 FrameStrobe_O[14] VPWR VGND sg13g2_buf_1
Xoutput49 net49 FrameStrobe_O[6] VPWR VGND sg13g2_buf_1
Xoutput16 net16 FrameData_O[23] VPWR VGND sg13g2_buf_1
Xoutput27 net27 FrameData_O[4] VPWR VGND sg13g2_buf_1
XFILLER_11_7 VPWR VGND sg13g2_fill_2
XFILLER_8_359 VPWR VGND sg13g2_decap_8
X_004_ FrameData[4] net27 VPWR VGND sg13g2_buf_1
XFILLER_7_84 VPWR VGND sg13g2_decap_8
XFILLER_8_178 VPWR VGND sg13g2_fill_1
XFILLER_8_112 VPWR VGND sg13g2_decap_8
XFILLER_5_126 VPWR VGND sg13g2_fill_2
XFILLER_5_104 VPWR VGND sg13g2_fill_2
XFILLER_1_343 VPWR VGND sg13g2_decap_8
XFILLER_1_398 VPWR VGND sg13g2_decap_8
XFILLER_4_85 VPWR VGND sg13g2_decap_8
XFILLER_11_409 VPWR VGND sg13g2_decap_8
XFILLER_10_420 VPWR VGND sg13g2_decap_8
XFILLER_6_435 VPWR VGND sg13g2_decap_8
XFILLER_1_140 VPWR VGND sg13g2_decap_8
XFILLER_9_295 VPWR VGND sg13g2_decap_8
XFILLER_10_294 VPWR VGND sg13g2_decap_8
XFILLER_6_298 VPWR VGND sg13g2_decap_8
XFILLER_6_232 VPWR VGND sg13g2_decap_8
XFILLER_1_42 VPWR VGND sg13g2_decap_8
X_097_ NN4END[6] net104 VPWR VGND sg13g2_buf_1
X_020_ FrameData[20] net13 VPWR VGND sg13g2_buf_1
XFILLER_0_419 VPWR VGND sg13g2_decap_8
XFILLER_3_246 VPWR VGND sg13g2_decap_4
XFILLER_10_84 VPWR VGND sg13g2_decap_8
XFILLER_3_279 VPWR VGND sg13g2_decap_8
Xoutput39 net39 FrameStrobe_O[15] VPWR VGND sg13g2_buf_1
Xoutput17 net17 FrameData_O[24] VPWR VGND sg13g2_buf_1
Xoutput28 net28 FrameData_O[5] VPWR VGND sg13g2_buf_1
XFILLER_8_338 VPWR VGND sg13g2_decap_8
X_003_ FrameData[3] net26 VPWR VGND sg13g2_buf_1
XFILLER_7_63 VPWR VGND sg13g2_decap_8
XFILLER_4_363 VPWR VGND sg13g2_decap_8
XFILLER_4_341 VPWR VGND sg13g2_fill_2
XFILLER_4_330 VPWR VGND sg13g2_decap_8
XFILLER_9_433 VPWR VGND sg13g2_decap_8
XFILLER_1_322 VPWR VGND sg13g2_decap_8
XFILLER_1_377 VPWR VGND sg13g2_decap_8
XFILLER_4_42 VPWR VGND sg13g2_decap_8
XFILLER_2_119 VPWR VGND sg13g2_decap_8
XFILLER_8_0 VPWR VGND sg13g2_decap_8
XFILLER_6_414 VPWR VGND sg13g2_decap_8
XFILLER_1_196 VPWR VGND sg13g2_decap_8
XFILLER_11_218 VPWR VGND sg13g2_decap_8
XFILLER_1_7 VPWR VGND sg13g2_decap_8
XFILLER_10_273 VPWR VGND sg13g2_decap_8
XFILLER_6_211 VPWR VGND sg13g2_decap_8
XFILLER_1_98 VPWR VGND sg13g2_decap_8
XFILLER_1_21 VPWR VGND sg13g2_decap_8
X_096_ NN4END[7] net103 VPWR VGND sg13g2_buf_1
XFILLER_10_63 VPWR VGND sg13g2_decap_8
Xoutput18 net18 FrameData_O[25] VPWR VGND sg13g2_buf_1
X_079_ N4END[8] net86 VPWR VGND sg13g2_buf_1
Xoutput29 net29 FrameData_O[6] VPWR VGND sg13g2_buf_1
XFILLER_8_317 VPWR VGND sg13g2_decap_8
X_002_ FrameData[2] net23 VPWR VGND sg13g2_buf_1
XFILLER_7_394 VPWR VGND sg13g2_decap_8
XFILLER_7_42 VPWR VGND sg13g2_decap_8
XFILLER_5_309 VPWR VGND sg13g2_decap_8
XFILLER_8_147 VPWR VGND sg13g2_decap_8
XFILLER_9_412 VPWR VGND sg13g2_decap_8
XFILLER_5_139 VPWR VGND sg13g2_decap_8
XFILLER_5_106 VPWR VGND sg13g2_fill_1
XFILLER_1_356 VPWR VGND sg13g2_decap_8
XFILLER_4_21 VPWR VGND sg13g2_decap_8
XFILLER_4_183 VPWR VGND sg13g2_decap_8
XFILLER_1_175 VPWR VGND sg13g2_decap_8
XFILLER_3_407 VPWR VGND sg13g2_fill_2
XFILLER_10_252 VPWR VGND sg13g2_decap_8
XFILLER_6_278 VPWR VGND sg13g2_fill_2
XFILLER_6_267 VPWR VGND sg13g2_decap_8
XFILLER_1_77 VPWR VGND sg13g2_decap_8
X_095_ NN4END[8] net102 VPWR VGND sg13g2_buf_1
XFILLER_10_42 VPWR VGND sg13g2_decap_8
XFILLER_3_226 VPWR VGND sg13g2_decap_8
XFILLER_3_259 VPWR VGND sg13g2_fill_1
X_078_ N4END[9] net85 VPWR VGND sg13g2_buf_1
XFILLER_2_292 VPWR VGND sg13g2_decap_8
Xoutput19 net19 FrameData_O[26] VPWR VGND sg13g2_buf_1
X_001_ FrameData[1] net12 VPWR VGND sg13g2_buf_1
XFILLER_7_373 VPWR VGND sg13g2_decap_8
XFILLER_7_98 VPWR VGND sg13g2_decap_8
XFILLER_7_21 VPWR VGND sg13g2_decap_8
XFILLER_8_126 VPWR VGND sg13g2_decap_8
XFILLER_4_99 VPWR VGND sg13g2_decap_8
XFILLER_4_162 VPWR VGND sg13g2_decap_8
XFILLER_10_434 VPWR VGND sg13g2_decap_8
XFILLER_6_449 VPWR VGND sg13g2_fill_2
XFILLER_9_243 VPWR VGND sg13g2_decap_8
XFILLER_1_154 VPWR VGND sg13g2_decap_8
XFILLER_10_231 VPWR VGND sg13g2_decap_8
XFILLER_6_246 VPWR VGND sg13g2_decap_8
X_094_ NN4END[9] net101 VPWR VGND sg13g2_buf_1
XFILLER_1_56 VPWR VGND sg13g2_decap_8
XFILLER_10_98 VPWR VGND sg13g2_decap_8
XFILLER_10_21 VPWR VGND sg13g2_decap_8
XFILLER_3_205 VPWR VGND sg13g2_decap_8
X_077_ N4END[10] net84 VPWR VGND sg13g2_buf_1
XFILLER_7_352 VPWR VGND sg13g2_decap_8
XFILLER_7_77 VPWR VGND sg13g2_decap_8
X_000_ FrameData[0] net1 VPWR VGND sg13g2_buf_1
XFILLER_8_105 VPWR VGND sg13g2_decap_8
XFILLER_4_377 VPWR VGND sg13g2_fill_2
XFILLER_5_119 VPWR VGND sg13g2_decap_8
XFILLER_1_336 VPWR VGND sg13g2_decap_8
XFILLER_9_447 VPWR VGND sg13g2_decap_4
XFILLER_0_391 VPWR VGND sg13g2_decap_8
XFILLER_4_56 VPWR VGND sg13g2_decap_4
XFILLER_4_78 VPWR VGND sg13g2_decap_8
XFILLER_4_141 VPWR VGND sg13g2_decap_8
XFILLER_10_413 VPWR VGND sg13g2_decap_8
XFILLER_6_428 VPWR VGND sg13g2_decap_8
XFILLER_1_133 VPWR VGND sg13g2_decap_8
XFILLER_9_288 VPWR VGND sg13g2_fill_2
XFILLER_5_450 VPWR VGND sg13g2_fill_1
XFILLER_10_287 VPWR VGND sg13g2_decap_8
XFILLER_10_210 VPWR VGND sg13g2_decap_8
XFILLER_6_225 VPWR VGND sg13g2_decap_8
XFILLER_6_0 VPWR VGND sg13g2_decap_8
X_093_ NN4END[10] net100 VPWR VGND sg13g2_buf_1
XFILLER_1_35 VPWR VGND sg13g2_decap_8
XFILLER_2_442 VPWR VGND sg13g2_decap_8
XFILLER_10_77 VPWR VGND sg13g2_decap_8
X_076_ N4END[11] net83 VPWR VGND sg13g2_buf_1
XFILLER_7_331 VPWR VGND sg13g2_decap_8
XFILLER_7_56 VPWR VGND sg13g2_decap_8
X_059_ N2MID[4] net60 VPWR VGND sg13g2_buf_1
XFILLER_4_323 VPWR VGND sg13g2_decap_8
XFILLER_4_356 VPWR VGND sg13g2_decap_8
XFILLER_1_315 VPWR VGND sg13g2_decap_8
XFILLER_9_426 VPWR VGND sg13g2_decap_8
XFILLER_0_370 VPWR VGND sg13g2_decap_8
XFILLER_4_35 VPWR VGND sg13g2_decap_8
XFILLER_4_120 VPWR VGND sg13g2_decap_8
XFILLER_4_197 VPWR VGND sg13g2_decap_8
XFILLER_6_407 VPWR VGND sg13g2_decap_8
XFILLER_1_189 VPWR VGND sg13g2_decap_8
XFILLER_1_112 VPWR VGND sg13g2_decap_8
XFILLER_9_201 VPWR VGND sg13g2_decap_8
XFILLER_10_266 VPWR VGND sg13g2_decap_8
XFILLER_6_204 VPWR VGND sg13g2_decap_8
X_092_ NN4END[11] net99 VPWR VGND sg13g2_buf_1
XFILLER_1_14 VPWR VGND sg13g2_decap_8
XFILLER_2_421 VPWR VGND sg13g2_decap_8
XFILLER_10_56 VPWR VGND sg13g2_decap_8
XFILLER_5_281 VPWR VGND sg13g2_decap_8
X_075_ N4END[12] net82 VPWR VGND sg13g2_buf_1
XFILLER_11_394 VPWR VGND sg13g2_decap_8
XFILLER_11_372 VPWR VGND sg13g2_decap_8
XFILLER_11_350 VPWR VGND sg13g2_decap_8
XFILLER_7_387 VPWR VGND sg13g2_decap_8
XFILLER_7_310 VPWR VGND sg13g2_decap_8
XFILLER_7_35 VPWR VGND sg13g2_decap_8
X_058_ N2MID[5] net59 VPWR VGND sg13g2_buf_1
XFILLER_4_379 VPWR VGND sg13g2_fill_1
XFILLER_4_302 VPWR VGND sg13g2_decap_8
XFILLER_9_405 VPWR VGND sg13g2_decap_8
XFILLER_4_14 VPWR VGND sg13g2_decap_8
XFILLER_4_176 VPWR VGND sg13g2_decap_8
XFILLER_1_168 VPWR VGND sg13g2_decap_8
XFILLER_5_441 VPWR VGND sg13g2_decap_8
XFILLER_10_245 VPWR VGND sg13g2_decap_8
X_091_ NN4END[12] net98 VPWR VGND sg13g2_buf_1
XFILLER_2_400 VPWR VGND sg13g2_decap_8
XFILLER_5_260 VPWR VGND sg13g2_decap_8
XFILLER_10_35 VPWR VGND sg13g2_decap_8
X_074_ N4END[13] net81 VPWR VGND sg13g2_buf_1
XFILLER_3_219 VPWR VGND sg13g2_decap_8
XFILLER_2_252 VPWR VGND sg13g2_decap_4
XFILLER_2_285 VPWR VGND sg13g2_decap_8
XFILLER_2_91 VPWR VGND sg13g2_decap_8
XFILLER_7_366 VPWR VGND sg13g2_decap_8
XFILLER_7_14 VPWR VGND sg13g2_decap_8
X_057_ N2MID[6] net58 VPWR VGND sg13g2_buf_1
XFILLER_8_119 VPWR VGND sg13g2_decap_8
XFILLER_11_181 VPWR VGND sg13g2_decap_4
XFILLER_3_380 VPWR VGND sg13g2_decap_8
XFILLER_8_450 VPWR VGND sg13g2_fill_1
XFILLER_4_155 VPWR VGND sg13g2_decap_8
XFILLER_10_427 VPWR VGND sg13g2_decap_8
XFILLER_1_147 VPWR VGND sg13g2_decap_8
XFILLER_5_420 VPWR VGND sg13g2_decap_8
XFILLER_10_224 VPWR VGND sg13g2_decap_8
XFILLER_6_239 VPWR VGND sg13g2_decap_8
X_090_ NN4END[13] net97 VPWR VGND sg13g2_buf_1
XFILLER_1_49 VPWR VGND sg13g2_decap_8
XFILLER_10_14 VPWR VGND sg13g2_decap_8
X_073_ N4END[14] net80 VPWR VGND sg13g2_buf_1
XFILLER_2_231 VPWR VGND sg13g2_decap_8
XFILLER_4_0 VPWR VGND sg13g2_decap_8
XFILLER_2_70 VPWR VGND sg13g2_decap_8
XANTENNA_20 VPWR VGND FrameData[6] sg13g2_antennanp
XFILLER_7_345 VPWR VGND sg13g2_decap_8
X_056_ N2MID[7] net57 VPWR VGND sg13g2_buf_1
XFILLER_4_337 VPWR VGND sg13g2_decap_4
X_039_ FrameStrobe[7] net50 VPWR VGND sg13g2_buf_1
XFILLER_8_91 VPWR VGND sg13g2_decap_8
XFILLER_1_329 VPWR VGND sg13g2_decap_8
XFILLER_0_384 VPWR VGND sg13g2_decap_8
XFILLER_4_49 VPWR VGND sg13g2_decap_8
XFILLER_4_134 VPWR VGND sg13g2_decap_8
XFILLER_10_406 VPWR VGND sg13g2_decap_8
XFILLER_9_237 VPWR VGND sg13g2_fill_2
XFILLER_8_7 VPWR VGND sg13g2_decap_8
XFILLER_1_126 VPWR VGND sg13g2_decap_8
XFILLER_8_281 VPWR VGND sg13g2_decap_4
XFILLER_5_70 VPWR VGND sg13g2_decap_8
XFILLER_10_203 VPWR VGND sg13g2_decap_8
XFILLER_6_218 VPWR VGND sg13g2_decap_8
XFILLER_1_28 VPWR VGND sg13g2_decap_8
XFILLER_2_435 VPWR VGND sg13g2_decap_8
XFILLER_5_295 VPWR VGND sg13g2_decap_8
X_072_ N4END[15] net73 VPWR VGND sg13g2_buf_1
XFILLER_2_210 VPWR VGND sg13g2_decap_8
XANTENNA_10 VPWR VGND FrameData[12] sg13g2_antennanp
XANTENNA_21 VPWR VGND FrameData[6] sg13g2_antennanp
XFILLER_7_324 VPWR VGND sg13g2_decap_8
XFILLER_7_49 VPWR VGND sg13g2_decap_8
X_055_ N1END[0] net56 VPWR VGND sg13g2_buf_1
XFILLER_4_349 VPWR VGND sg13g2_decap_8
XFILLER_4_316 VPWR VGND sg13g2_decap_8
X_038_ FrameStrobe[6] net49 VPWR VGND sg13g2_buf_1
XFILLER_7_154 VPWR VGND sg13g2_fill_1
XFILLER_7_121 VPWR VGND sg13g2_decap_8
XFILLER_8_70 VPWR VGND sg13g2_decap_8
XFILLER_9_419 VPWR VGND sg13g2_decap_8
XFILLER_0_363 VPWR VGND sg13g2_decap_8
XFILLER_4_28 VPWR VGND sg13g2_decap_8
XFILLER_4_113 VPWR VGND sg13g2_decap_8
XFILLER_1_105 VPWR VGND sg13g2_decap_8
XFILLER_8_260 VPWR VGND sg13g2_fill_1
XFILLER_0_182 VPWR VGND sg13g2_decap_8
XFILLER_10_259 VPWR VGND sg13g2_decap_8
XFILLER_5_82 VPWR VGND sg13g2_decap_8
XFILLER_2_414 VPWR VGND sg13g2_decap_8
XFILLER_5_274 VPWR VGND sg13g2_decap_8
XFILLER_10_49 VPWR VGND sg13g2_decap_8
X_071_ N2END[0] net72 VPWR VGND sg13g2_buf_1
XFILLER_2_299 VPWR VGND sg13g2_fill_1
XFILLER_11_321 VPWR VGND sg13g2_decap_8
XANTENNA_11 VPWR VGND FrameData[3] sg13g2_antennanp
XANTENNA_22 VPWR VGND FrameData[6] sg13g2_antennanp
XFILLER_11_387 VPWR VGND sg13g2_decap_8
XFILLER_11_365 VPWR VGND sg13g2_decap_8
XFILLER_11_343 VPWR VGND sg13g2_decap_8
XFILLER_7_303 VPWR VGND sg13g2_decap_8
XFILLER_7_28 VPWR VGND sg13g2_decap_8
X_054_ N1END[1] net55 VPWR VGND sg13g2_buf_1
X_037_ FrameStrobe[5] net48 VPWR VGND sg13g2_buf_1
XFILLER_3_394 VPWR VGND sg13g2_fill_2
XFILLER_0_342 VPWR VGND sg13g2_decap_8
XFILLER_4_169 VPWR VGND sg13g2_decap_8
XFILLER_3_191 VPWR VGND sg13g2_decap_8
XFILLER_5_434 VPWR VGND sg13g2_decap_8
XFILLER_0_161 VPWR VGND sg13g2_decap_8
XFILLER_10_238 VPWR VGND sg13g2_decap_8
XFILLER_8_272 VPWR VGND sg13g2_decap_4
XFILLER_5_94 VPWR VGND sg13g2_decap_4
XFILLER_5_61 VPWR VGND sg13g2_decap_4
XFILLER_5_253 VPWR VGND sg13g2_decap_8
XFILLER_10_28 VPWR VGND sg13g2_decap_8
X_070_ N2END[1] net71 VPWR VGND sg13g2_buf_1
XFILLER_2_245 VPWR VGND sg13g2_decap_8
XFILLER_2_256 VPWR VGND sg13g2_fill_1
XFILLER_2_84 VPWR VGND sg13g2_decap_8
XANTENNA_12 VPWR VGND FrameData[4] sg13g2_antennanp
XANTENNA_23 VPWR VGND FrameData[6] sg13g2_antennanp
XFILLER_11_93 VPWR VGND sg13g2_decap_4
XFILLER_11_71 VPWR VGND sg13g2_decap_4
XFILLER_7_359 VPWR VGND sg13g2_decap_8
XFILLER_2_0 VPWR VGND sg13g2_decap_8
X_053_ N1END[2] net54 VPWR VGND sg13g2_buf_1
XFILLER_11_196 VPWR VGND sg13g2_decap_8
XFILLER_11_174 VPWR VGND sg13g2_decap_8
XFILLER_11_152 VPWR VGND sg13g2_decap_8
XFILLER_11_130 VPWR VGND sg13g2_decap_8
XFILLER_7_112 VPWR VGND sg13g2_decap_4
X_036_ FrameStrobe[4] net47 VPWR VGND sg13g2_buf_1
XFILLER_7_167 VPWR VGND sg13g2_fill_1
XFILLER_3_373 VPWR VGND sg13g2_decap_8
XFILLER_0_321 VPWR VGND sg13g2_decap_8
XFILLER_4_148 VPWR VGND sg13g2_decap_8
XFILLER_8_443 VPWR VGND sg13g2_decap_8
XFILLER_0_398 VPWR VGND sg13g2_decap_8
XFILLER_3_170 VPWR VGND sg13g2_decap_8
X_019_ FrameData[19] net11 VPWR VGND sg13g2_buf_1
XFILLER_5_413 VPWR VGND sg13g2_decap_8
XFILLER_0_140 VPWR VGND sg13g2_decap_8
XFILLER_8_251 VPWR VGND sg13g2_fill_1
XFILLER_10_217 VPWR VGND sg13g2_decap_8
XFILLER_6_7 VPWR VGND sg13g2_decap_8
XFILLER_2_449 VPWR VGND sg13g2_fill_2
XFILLER_5_232 VPWR VGND sg13g2_decap_8
XFILLER_2_224 VPWR VGND sg13g2_decap_8
XANTENNA_13 VPWR VGND FrameData[5] sg13g2_antennanp
XFILLER_2_63 VPWR VGND sg13g2_decap_8
XANTENNA_24 VPWR VGND FrameData[6] sg13g2_antennanp
XFILLER_7_338 VPWR VGND sg13g2_decap_8
X_052_ N1END[3] net53 VPWR VGND sg13g2_buf_1
XFILLER_6_393 VPWR VGND sg13g2_decap_8
X_035_ FrameStrobe[3] net46 VPWR VGND sg13g2_buf_1
X_104_ UserCLK net105 VPWR VGND sg13g2_buf_1
XFILLER_3_352 VPWR VGND sg13g2_decap_8
XFILLER_3_396 VPWR VGND sg13g2_fill_1
XFILLER_8_84 VPWR VGND sg13g2_decap_8
XFILLER_8_422 VPWR VGND sg13g2_decap_8
XFILLER_0_377 VPWR VGND sg13g2_decap_8
X_018_ FrameData[18] net10 VPWR VGND sg13g2_buf_1
XFILLER_4_127 VPWR VGND sg13g2_decap_8
XFILLER_1_119 VPWR VGND sg13g2_decap_8
XFILLER_9_208 VPWR VGND sg13g2_fill_1
XFILLER_0_196 VPWR VGND sg13g2_decap_8
XFILLER_10_0 VPWR VGND sg13g2_decap_8
XFILLER_8_296 VPWR VGND sg13g2_decap_8
XFILLER_2_428 VPWR VGND sg13g2_decap_8
XFILLER_5_288 VPWR VGND sg13g2_decap_8
XFILLER_2_203 VPWR VGND sg13g2_decap_8
XFILLER_9_391 VPWR VGND sg13g2_decap_8
XANTENNA_25 VPWR VGND FrameData[6] sg13g2_antennanp
XFILLER_2_42 VPWR VGND sg13g2_decap_8
XANTENNA_14 VPWR VGND FrameData[5] sg13g2_antennanp
XFILLER_11_379 VPWR VGND sg13g2_decap_4
XFILLER_11_357 VPWR VGND sg13g2_decap_4
XFILLER_11_335 VPWR VGND sg13g2_decap_4
XFILLER_11_313 VPWR VGND sg13g2_decap_4
XFILLER_7_317 VPWR VGND sg13g2_decap_8
X_051_ FrameStrobe[19] net43 VPWR VGND sg13g2_buf_1
XFILLER_6_372 VPWR VGND sg13g2_decap_8
XFILLER_4_309 VPWR VGND sg13g2_decap_8
X_034_ FrameStrobe[2] net45 VPWR VGND sg13g2_buf_1
XFILLER_7_147 VPWR VGND sg13g2_decap_8
XFILLER_7_136 VPWR VGND sg13g2_decap_8
XFILLER_3_331 VPWR VGND sg13g2_decap_8
X_103_ NN4END[0] net95 VPWR VGND sg13g2_buf_1
XFILLER_8_63 VPWR VGND sg13g2_decap_8
XFILLER_8_401 VPWR VGND sg13g2_decap_8
XFILLER_0_356 VPWR VGND sg13g2_decap_8
XFILLER_4_106 VPWR VGND sg13g2_decap_8
X_017_ FrameData[17] net9 VPWR VGND sg13g2_buf_1
XFILLER_5_448 VPWR VGND sg13g2_fill_2
XFILLER_5_42 VPWR VGND sg13g2_decap_8
XFILLER_0_175 VPWR VGND sg13g2_decap_8
XFILLER_2_407 VPWR VGND sg13g2_decap_8
XFILLER_5_267 VPWR VGND sg13g2_decap_8
XFILLER_1_440 VPWR VGND sg13g2_decap_8
XFILLER_9_370 VPWR VGND sg13g2_decap_8
XANTENNA_15 VPWR VGND FrameData[6] sg13g2_antennanp
XFILLER_2_21 VPWR VGND sg13g2_decap_8
XFILLER_2_98 VPWR VGND sg13g2_decap_8
Xoutput100 net100 SS4BEG[5] VPWR VGND sg13g2_buf_1
X_050_ FrameStrobe[18] net42 VPWR VGND sg13g2_buf_1
XFILLER_6_351 VPWR VGND sg13g2_decap_8
X_033_ FrameStrobe[1] net44 VPWR VGND sg13g2_buf_1
XFILLER_7_159 VPWR VGND sg13g2_decap_4
XFILLER_0_0 VPWR VGND sg13g2_decap_8
XFILLER_3_321 VPWR VGND sg13g2_decap_4
XFILLER_3_387 VPWR VGND sg13g2_decap_8
X_102_ NN4END[1] net94 VPWR VGND sg13g2_buf_1
XFILLER_8_42 VPWR VGND sg13g2_decap_8
XFILLER_6_181 VPWR VGND sg13g2_decap_8
XFILLER_0_335 VPWR VGND sg13g2_decap_8
X_016_ FrameData[16] net8 VPWR VGND sg13g2_buf_1
XFILLER_3_184 VPWR VGND sg13g2_decap_8
XFILLER_8_276 VPWR VGND sg13g2_fill_1
XFILLER_8_265 VPWR VGND sg13g2_decap_8
XFILLER_8_243 VPWR VGND sg13g2_fill_2
XFILLER_5_427 VPWR VGND sg13g2_decap_8
XFILLER_5_21 VPWR VGND sg13g2_decap_8
XFILLER_0_154 VPWR VGND sg13g2_decap_8
XFILLER_5_98 VPWR VGND sg13g2_fill_2
XFILLER_5_65 VPWR VGND sg13g2_fill_1
XFILLER_5_246 VPWR VGND sg13g2_decap_8
XFILLER_5_202 VPWR VGND sg13g2_decap_4
XFILLER_2_238 VPWR VGND sg13g2_decap_8
XFILLER_4_7 VPWR VGND sg13g2_decap_8
XFILLER_2_77 VPWR VGND sg13g2_decap_8
Xoutput101 net101 SS4BEG[6] VPWR VGND sg13g2_buf_1
XANTENNA_16 VPWR VGND FrameData[6] sg13g2_antennanp
XFILLER_11_86 VPWR VGND sg13g2_decap_8
XFILLER_11_64 VPWR VGND sg13g2_decap_8
XFILLER_11_42 VPWR VGND sg13g2_decap_8
XFILLER_11_20 VPWR VGND sg13g2_decap_8
XFILLER_10_392 VPWR VGND sg13g2_decap_8
XFILLER_11_189 VPWR VGND sg13g2_decap_8
XFILLER_11_167 VPWR VGND sg13g2_decap_8
XFILLER_11_145 VPWR VGND sg13g2_decap_8
XFILLER_11_123 VPWR VGND sg13g2_decap_8
XFILLER_11_101 VPWR VGND sg13g2_decap_8
X_032_ FrameStrobe[0] net33 VPWR VGND sg13g2_buf_1
XFILLER_7_116 VPWR VGND sg13g2_fill_1
XFILLER_7_105 VPWR VGND sg13g2_decap_8
XFILLER_3_300 VPWR VGND sg13g2_decap_8
XFILLER_3_366 VPWR VGND sg13g2_decap_8
X_101_ NN4END[2] net93 VPWR VGND sg13g2_buf_1
XFILLER_8_98 VPWR VGND sg13g2_decap_8
XFILLER_8_21 VPWR VGND sg13g2_decap_8
XFILLER_6_160 VPWR VGND sg13g2_decap_8
XFILLER_8_436 VPWR VGND sg13g2_decap_8
X_015_ FrameData[15] net7 VPWR VGND sg13g2_buf_1
XFILLER_3_163 VPWR VGND sg13g2_decap_8
XFILLER_5_406 VPWR VGND sg13g2_decap_8
XFILLER_0_133 VPWR VGND sg13g2_decap_8
XFILLER_8_222 VPWR VGND sg13g2_decap_8
XFILLER_5_77 VPWR VGND sg13g2_fill_1
XFILLER_5_225 VPWR VGND sg13g2_decap_8
XFILLER_2_217 VPWR VGND sg13g2_decap_8
XFILLER_2_56 VPWR VGND sg13g2_decap_8
XANTENNA_17 VPWR VGND FrameData[8] sg13g2_antennanp
Xoutput102 net102 SS4BEG[7] VPWR VGND sg13g2_buf_1
XFILLER_10_371 VPWR VGND sg13g2_decap_8
XFILLER_6_386 VPWR VGND sg13g2_decap_8
X_031_ FrameData[31] net25 VPWR VGND sg13g2_buf_1
XFILLER_7_128 VPWR VGND sg13g2_decap_4
X_100_ NN4END[3] net92 VPWR VGND sg13g2_buf_1
XFILLER_8_77 VPWR VGND sg13g2_decap_8
XFILLER_3_345 VPWR VGND sg13g2_decap_8
XFILLER_8_415 VPWR VGND sg13g2_decap_8
X_014_ FrameData[14] net6 VPWR VGND sg13g2_buf_1
XFILLER_3_142 VPWR VGND sg13g2_decap_8
XFILLER_0_189 VPWR VGND sg13g2_decap_8
XFILLER_0_112 VPWR VGND sg13g2_decap_8
XFILLER_8_289 VPWR VGND sg13g2_decap_8
XFILLER_8_256 VPWR VGND sg13g2_decap_4
XFILLER_8_201 VPWR VGND sg13g2_decap_8
XFILLER_5_89 VPWR VGND sg13g2_fill_1
XFILLER_5_56 VPWR VGND sg13g2_fill_1
XFILLER_4_440 VPWR VGND sg13g2_decap_8
XFILLER_9_384 VPWR VGND sg13g2_decap_8
XANTENNA_18 VPWR VGND FrameData[5] sg13g2_antennanp
Xoutput103 net103 SS4BEG[8] VPWR VGND sg13g2_buf_1
XFILLER_2_35 VPWR VGND sg13g2_decap_8
XFILLER_11_328 VPWR VGND sg13g2_decap_8
XFILLER_11_306 VPWR VGND sg13g2_decap_8
XFILLER_10_350 VPWR VGND sg13g2_decap_8
XFILLER_6_365 VPWR VGND sg13g2_decap_8
XFILLER_9_181 VPWR VGND sg13g2_fill_2
XFILLER_9_170 VPWR VGND sg13g2_decap_8
X_030_ FrameData[30] net24 VPWR VGND sg13g2_buf_1
XFILLER_8_56 VPWR VGND sg13g2_decap_8
XFILLER_0_349 VPWR VGND sg13g2_decap_8
X_013_ FrameData[13] net5 VPWR VGND sg13g2_buf_1
XFILLER_3_121 VPWR VGND sg13g2_decap_8
XFILLER_3_198 VPWR VGND sg13g2_decap_8
XFILLER_0_168 VPWR VGND sg13g2_decap_8
XFILLER_5_35 VPWR VGND sg13g2_decap_8
XFILLER_1_433 VPWR VGND sg13g2_decap_8
XFILLER_4_271 VPWR VGND sg13g2_decap_4
XFILLER_9_363 VPWR VGND sg13g2_decap_8
XFILLER_9_0 VPWR VGND sg13g2_decap_8
Xoutput104 net104 SS4BEG[9] VPWR VGND sg13g2_buf_1
XFILLER_2_14 VPWR VGND sg13g2_decap_8
XANTENNA_19 VPWR VGND FrameData[6] sg13g2_antennanp
XFILLER_2_7 VPWR VGND sg13g2_decap_8
XFILLER_6_344 VPWR VGND sg13g2_decap_8
XFILLER_11_159 VPWR VGND sg13g2_decap_4
XFILLER_11_137 VPWR VGND sg13g2_decap_4
XFILLER_11_115 VPWR VGND sg13g2_decap_4
XFILLER_3_314 VPWR VGND sg13g2_decap_8
XFILLER_3_325 VPWR VGND sg13g2_fill_2
XFILLER_8_35 VPWR VGND sg13g2_decap_8
X_089_ NN4END[14] net96 VPWR VGND sg13g2_buf_1
XFILLER_6_174 VPWR VGND sg13g2_decap_8
XFILLER_0_328 VPWR VGND sg13g2_decap_8
XFILLER_7_450 VPWR VGND sg13g2_fill_1
X_012_ FrameData[12] net4 VPWR VGND sg13g2_buf_1
XFILLER_3_100 VPWR VGND sg13g2_decap_8
XFILLER_3_177 VPWR VGND sg13g2_decap_8
XFILLER_0_91 VPWR VGND sg13g2_decap_8
XFILLER_8_236 VPWR VGND sg13g2_decap_8
XFILLER_5_14 VPWR VGND sg13g2_decap_8
XFILLER_0_147 VPWR VGND sg13g2_decap_8
XFILLER_5_239 VPWR VGND sg13g2_decap_8
XFILLER_1_412 VPWR VGND sg13g2_decap_8
XFILLER_9_342 VPWR VGND sg13g2_decap_8
XFILLER_11_57 VPWR VGND sg13g2_decap_8
XFILLER_11_35 VPWR VGND sg13g2_decap_8
Xoutput105 net105 UserCLKo VPWR VGND sg13g2_buf_1
XFILLER_11_13 VPWR VGND sg13g2_decap_8
XFILLER_11_79 VPWR VGND sg13g2_decap_8
XFILLER_10_385 VPWR VGND sg13g2_decap_8
XFILLER_6_312 VPWR VGND sg13g2_decap_8
XFILLER_9_194 VPWR VGND sg13g2_decap_8
XFILLER_3_359 VPWR VGND sg13g2_decap_8
XFILLER_10_182 VPWR VGND sg13g2_decap_8
XFILLER_8_14 VPWR VGND sg13g2_decap_8
X_088_ NN4END[15] net89 VPWR VGND sg13g2_buf_1
XFILLER_6_153 VPWR VGND sg13g2_decap_8
XFILLER_2_381 VPWR VGND sg13g2_fill_1
XFILLER_8_429 VPWR VGND sg13g2_decap_8
X_011_ FrameData[11] net3 VPWR VGND sg13g2_buf_1
XFILLER_3_156 VPWR VGND sg13g2_decap_8
XFILLER_0_70 VPWR VGND sg13g2_decap_8
XFILLER_8_215 VPWR VGND sg13g2_decap_8
XFILLER_0_126 VPWR VGND sg13g2_decap_8
XFILLER_10_7 VPWR VGND sg13g2_decap_8
XFILLER_5_218 VPWR VGND sg13g2_decap_8
XFILLER_4_295 VPWR VGND sg13g2_decap_8
XFILLER_6_91 VPWR VGND sg13g2_decap_8
XFILLER_2_49 VPWR VGND sg13g2_decap_8
XFILLER_9_398 VPWR VGND sg13g2_decap_8
XFILLER_9_321 VPWR VGND sg13g2_decap_8
XFILLER_10_364 VPWR VGND sg13g2_decap_8
XFILLER_6_379 VPWR VGND sg13g2_decap_8
XFILLER_3_338 VPWR VGND sg13g2_decap_8
XFILLER_10_161 VPWR VGND sg13g2_decap_8
X_087_ N4END[0] net79 VPWR VGND sg13g2_buf_1
XFILLER_6_132 VPWR VGND sg13g2_decap_8
XFILLER_2_393 VPWR VGND sg13g2_decap_8
XFILLER_8_408 VPWR VGND sg13g2_decap_8
X_010_ FrameData[10] net2 VPWR VGND sg13g2_buf_1
XFILLER_3_135 VPWR VGND sg13g2_decap_8
XFILLER_0_105 VPWR VGND sg13g2_decap_8
XFILLER_8_249 VPWR VGND sg13g2_fill_2
XFILLER_5_49 VPWR VGND sg13g2_decap_8
XFILLER_4_433 VPWR VGND sg13g2_decap_8
XFILLER_7_282 VPWR VGND sg13g2_decap_8
XFILLER_4_230 VPWR VGND sg13g2_fill_1
XFILLER_4_263 VPWR VGND sg13g2_decap_4
XFILLER_6_70 VPWR VGND sg13g2_decap_8
XFILLER_1_244 VPWR VGND sg13g2_decap_8
XFILLER_2_28 VPWR VGND sg13g2_decap_8
XFILLER_9_377 VPWR VGND sg13g2_decap_8
XFILLER_10_343 VPWR VGND sg13g2_decap_8
XFILLER_7_0 VPWR VGND sg13g2_decap_8
XFILLER_6_358 VPWR VGND sg13g2_decap_8
XFILLER_9_163 VPWR VGND sg13g2_decap_8
XFILLER_5_380 VPWR VGND sg13g2_fill_1
XFILLER_3_60 VPWR VGND sg13g2_fill_1
XFILLER_3_93 VPWR VGND sg13g2_decap_8
XFILLER_10_140 VPWR VGND sg13g2_decap_8
X_086_ N4END[1] net78 VPWR VGND sg13g2_buf_1
XFILLER_8_49 VPWR VGND sg13g2_decap_8
XFILLER_6_199 VPWR VGND sg13g2_fill_1
XFILLER_6_188 VPWR VGND sg13g2_decap_8
XFILLER_6_111 VPWR VGND sg13g2_decap_8
XFILLER_0_7 VPWR VGND sg13g2_decap_8
XFILLER_2_361 VPWR VGND sg13g2_decap_8
XFILLER_2_372 VPWR VGND sg13g2_decap_8
XFILLER_3_114 VPWR VGND sg13g2_decap_8
X_069_ N2END[2] net70 VPWR VGND sg13g2_buf_1
XFILLER_9_81 VPWR VGND sg13g2_decap_8
XFILLER_5_28 VPWR VGND sg13g2_decap_8
XFILLER_7_261 VPWR VGND sg13g2_decap_8
XFILLER_1_426 VPWR VGND sg13g2_decap_8
XFILLER_4_242 VPWR VGND sg13g2_decap_8
XFILLER_4_275 VPWR VGND sg13g2_fill_1
XFILLER_9_356 VPWR VGND sg13g2_decap_8
Xoutput90 net90 SS4BEG[10] VPWR VGND sg13g2_buf_1
XFILLER_11_49 VPWR VGND sg13g2_decap_4
XFILLER_11_27 VPWR VGND sg13g2_decap_4
XFILLER_10_399 VPWR VGND sg13g2_decap_8
XFILLER_10_322 VPWR VGND sg13g2_decap_8
XFILLER_6_337 VPWR VGND sg13g2_decap_8
XFILLER_6_326 VPWR VGND sg13g2_decap_8
XFILLER_11_108 VPWR VGND sg13g2_decap_8
XFILLER_9_142 VPWR VGND sg13g2_decap_8
XFILLER_5_392 VPWR VGND sg13g2_decap_8
XFILLER_3_72 VPWR VGND sg13g2_decap_8
XFILLER_8_28 VPWR VGND sg13g2_decap_8
XFILLER_3_307 VPWR VGND sg13g2_decap_8
XFILLER_10_196 VPWR VGND sg13g2_decap_8
X_085_ N4END[2] net77 VPWR VGND sg13g2_buf_1
XFILLER_6_167 VPWR VGND sg13g2_decap_8
XFILLER_7_443 VPWR VGND sg13g2_decap_8
X_068_ N2END[3] net69 VPWR VGND sg13g2_buf_1
XFILLER_0_84 VPWR VGND sg13g2_decap_8
XFILLER_8_229 VPWR VGND sg13g2_decap_8
XFILLER_11_291 VPWR VGND sg13g2_decap_4
XFILLER_7_240 VPWR VGND sg13g2_decap_8
XFILLER_1_405 VPWR VGND sg13g2_decap_8
XFILLER_9_335 VPWR VGND sg13g2_decap_8
XFILLER_9_302 VPWR VGND sg13g2_decap_8
Xoutput1 net1 FrameData_O[0] VPWR VGND sg13g2_buf_1
Xoutput80 net80 S4BEG[1] VPWR VGND sg13g2_buf_1
Xoutput91 net91 SS4BEG[11] VPWR VGND sg13g2_buf_1
XFILLER_10_378 VPWR VGND sg13g2_decap_8
XFILLER_10_301 VPWR VGND sg13g2_decap_8
XFILLER_6_305 VPWR VGND sg13g2_decap_8
XFILLER_9_187 VPWR VGND sg13g2_decap_8
XFILLER_10_175 VPWR VGND sg13g2_decap_8
X_084_ N4END[3] net76 VPWR VGND sg13g2_buf_1
XFILLER_6_146 VPWR VGND sg13g2_decap_8
XFILLER_7_422 VPWR VGND sg13g2_decap_8
XFILLER_3_149 VPWR VGND sg13g2_decap_8
XFILLER_9_61 VPWR VGND sg13g2_decap_4
X_067_ N2END[4] net68 VPWR VGND sg13g2_buf_1
XFILLER_0_63 VPWR VGND sg13g2_decap_8
XFILLER_2_182 VPWR VGND sg13g2_decap_8
XFILLER_8_208 VPWR VGND sg13g2_decap_8
XFILLER_4_447 VPWR VGND sg13g2_decap_4
XFILLER_0_119 VPWR VGND sg13g2_decap_8
XFILLER_7_296 VPWR VGND sg13g2_decap_8
XFILLER_4_211 VPWR VGND sg13g2_decap_4
XFILLER_4_288 VPWR VGND sg13g2_decap_8
XFILLER_6_84 VPWR VGND sg13g2_decap_8
XFILLER_1_203 VPWR VGND sg13g2_decap_4
XFILLER_8_380 VPWR VGND sg13g2_decap_8
Xoutput81 net81 S4BEG[2] VPWR VGND sg13g2_buf_1
Xoutput70 net70 S2BEGb[5] VPWR VGND sg13g2_buf_1
Xoutput92 net92 SS4BEG[12] VPWR VGND sg13g2_buf_1
Xoutput2 net2 FrameData_O[10] VPWR VGND sg13g2_buf_1
XFILLER_10_357 VPWR VGND sg13g2_decap_8
XFILLER_9_177 VPWR VGND sg13g2_decap_4
XFILLER_5_361 VPWR VGND sg13g2_decap_8
XFILLER_10_154 VPWR VGND sg13g2_decap_8
X_083_ N4END[4] net75 VPWR VGND sg13g2_buf_1
XFILLER_6_125 VPWR VGND sg13g2_decap_8
XFILLER_5_0 VPWR VGND sg13g2_decap_8
XFILLER_2_386 VPWR VGND sg13g2_decap_8
XFILLER_3_128 VPWR VGND sg13g2_decap_8
XFILLER_9_95 VPWR VGND sg13g2_decap_8
XFILLER_9_51 VPWR VGND sg13g2_fill_1
XFILLER_7_401 VPWR VGND sg13g2_decap_8
X_066_ N2END[5] net67 VPWR VGND sg13g2_buf_1
XFILLER_0_42 VPWR VGND sg13g2_decap_8
XFILLER_2_161 VPWR VGND sg13g2_decap_8
XFILLER_4_426 VPWR VGND sg13g2_decap_8
XFILLER_4_404 VPWR VGND sg13g2_fill_1
XFILLER_7_275 VPWR VGND sg13g2_decap_8
X_049_ FrameStrobe[17] net41 VPWR VGND sg13g2_buf_1
XFILLER_0_440 VPWR VGND sg13g2_fill_2
XFILLER_4_256 VPWR VGND sg13g2_decap_8
XFILLER_6_63 VPWR VGND sg13g2_decap_8
XANTENNA_1 VPWR VGND FrameData[12] sg13g2_antennanp
XFILLER_9_7 VPWR VGND sg13g2_decap_8
XFILLER_1_237 VPWR VGND sg13g2_decap_8
Xoutput82 net82 S4BEG[3] VPWR VGND sg13g2_buf_1
Xoutput71 net71 S2BEGb[6] VPWR VGND sg13g2_buf_1
Xoutput60 net60 S2BEG[3] VPWR VGND sg13g2_buf_1
Xoutput93 net93 SS4BEG[13] VPWR VGND sg13g2_buf_1
Xoutput3 net3 FrameData_O[11] VPWR VGND sg13g2_buf_1
XFILLER_10_336 VPWR VGND sg13g2_decap_8
XFILLER_9_156 VPWR VGND sg13g2_decap_8
XFILLER_9_123 VPWR VGND sg13g2_fill_1
XFILLER_3_42 VPWR VGND sg13g2_decap_8
XFILLER_3_86 VPWR VGND sg13g2_decap_8
XFILLER_10_133 VPWR VGND sg13g2_decap_8
X_082_ N4END[5] net74 VPWR VGND sg13g2_buf_1
XFILLER_6_104 VPWR VGND sg13g2_decap_8
XFILLER_2_332 VPWR VGND sg13g2_decap_8
XFILLER_2_354 VPWR VGND sg13g2_decap_8
XFILLER_5_181 VPWR VGND sg13g2_decap_8
XFILLER_3_107 VPWR VGND sg13g2_decap_8
XFILLER_11_453 VPWR VGND sg13g2_fill_2
XFILLER_11_431 VPWR VGND sg13g2_decap_4
X_065_ N2END[6] net66 VPWR VGND sg13g2_buf_1
XFILLER_0_98 VPWR VGND sg13g2_decap_8
XFILLER_0_21 VPWR VGND sg13g2_decap_8
XFILLER_2_140 VPWR VGND sg13g2_decap_8
XFILLER_7_254 VPWR VGND sg13g2_decap_8
X_048_ FrameStrobe[16] net40 VPWR VGND sg13g2_buf_1
XFILLER_1_419 VPWR VGND sg13g2_decap_8
XFILLER_4_235 VPWR VGND sg13g2_decap_8
XFILLER_6_42 VPWR VGND sg13g2_decap_8
XANTENNA_2 VPWR VGND FrameData[2] sg13g2_antennanp
Xoutput50 net50 FrameStrobe_O[7] VPWR VGND sg13g2_buf_1
XFILLER_9_349 VPWR VGND sg13g2_decap_8
Xoutput4 net4 FrameData_O[12] VPWR VGND sg13g2_buf_1
Xoutput83 net83 S4BEG[4] VPWR VGND sg13g2_buf_1
Xoutput72 net72 S2BEGb[7] VPWR VGND sg13g2_buf_1
Xoutput61 net61 S2BEG[4] VPWR VGND sg13g2_buf_1
Xoutput94 net94 SS4BEG[14] VPWR VGND sg13g2_buf_1
XFILLER_10_315 VPWR VGND sg13g2_decap_8
XFILLER_9_135 VPWR VGND sg13g2_decap_8
XFILLER_9_102 VPWR VGND sg13g2_decap_8
XFILLER_6_319 VPWR VGND sg13g2_decap_8
XFILLER_5_341 VPWR VGND sg13g2_fill_2
XFILLER_5_330 VPWR VGND sg13g2_decap_8
XFILLER_3_21 VPWR VGND sg13g2_decap_8
XFILLER_3_65 VPWR VGND sg13g2_decap_8
XFILLER_10_189 VPWR VGND sg13g2_decap_8
XFILLER_10_112 VPWR VGND sg13g2_decap_8
X_081_ N4END[6] net88 VPWR VGND sg13g2_buf_1
XFILLER_2_311 VPWR VGND sg13g2_decap_8
XFILLER_5_160 VPWR VGND sg13g2_decap_8
XFILLER_7_436 VPWR VGND sg13g2_decap_8
X_064_ N2END[7] net65 VPWR VGND sg13g2_buf_1
XFILLER_2_196 VPWR VGND sg13g2_decap_8
XFILLER_9_42 VPWR VGND sg13g2_decap_8
XFILLER_0_77 VPWR VGND sg13g2_decap_8
XFILLER_11_284 VPWR VGND sg13g2_decap_8
XFILLER_11_262 VPWR VGND sg13g2_decap_8
XFILLER_11_240 VPWR VGND sg13g2_decap_8
XFILLER_7_233 VPWR VGND sg13g2_decap_8
X_047_ FrameStrobe[15] net39 VPWR VGND sg13g2_buf_1
XFILLER_6_98 VPWR VGND sg13g2_fill_2
XFILLER_6_21 VPWR VGND sg13g2_decap_8
XANTENNA_3 VPWR VGND FrameData[2] sg13g2_antennanp
XFILLER_0_442 VPWR VGND sg13g2_fill_1
XFILLER_4_225 VPWR VGND sg13g2_fill_1
Xoutput40 net40 FrameStrobe_O[16] VPWR VGND sg13g2_buf_1
Xoutput51 net51 FrameStrobe_O[8] VPWR VGND sg13g2_buf_1
XFILLER_9_328 VPWR VGND sg13g2_decap_8
Xoutput5 net5 FrameData_O[13] VPWR VGND sg13g2_buf_1
Xoutput84 net84 S4BEG[5] VPWR VGND sg13g2_buf_1
Xoutput73 net73 S4BEG[0] VPWR VGND sg13g2_buf_1
Xoutput62 net62 S2BEG[5] VPWR VGND sg13g2_buf_1
Xoutput95 net95 SS4BEG[15] VPWR VGND sg13g2_buf_1
XFILLER_8_394 VPWR VGND sg13g2_decap_8
XFILLER_10_168 VPWR VGND sg13g2_decap_8
X_080_ N4END[7] net87 VPWR VGND sg13g2_buf_1
XFILLER_6_139 VPWR VGND sg13g2_decap_8
XFILLER_7_415 VPWR VGND sg13g2_decap_8
X_063_ N2MID[0] net64 VPWR VGND sg13g2_buf_1
XFILLER_2_175 VPWR VGND sg13g2_decap_8
XFILLER_3_0 VPWR VGND sg13g2_decap_8
XFILLER_9_76 VPWR VGND sg13g2_fill_1
XFILLER_9_21 VPWR VGND sg13g2_decap_8
XFILLER_0_56 VPWR VGND sg13g2_decap_8
X_046_ FrameStrobe[14] net38 VPWR VGND sg13g2_buf_1
XFILLER_7_289 VPWR VGND sg13g2_decap_8
XFILLER_7_212 VPWR VGND sg13g2_decap_8
XFILLER_4_204 VPWR VGND sg13g2_decap_8
XFILLER_4_215 VPWR VGND sg13g2_fill_2
X_029_ FrameData[29] net22 VPWR VGND sg13g2_buf_1
XFILLER_6_77 VPWR VGND sg13g2_decap_8
XANTENNA_4 VPWR VGND FrameData[4] sg13g2_antennanp
Xoutput41 net41 FrameStrobe_O[17] VPWR VGND sg13g2_buf_1
Xoutput52 net52 FrameStrobe_O[9] VPWR VGND sg13g2_buf_1
Xoutput6 net6 FrameData_O[14] VPWR VGND sg13g2_buf_1
XFILLER_1_207 VPWR VGND sg13g2_fill_2
Xoutput30 net30 FrameData_O[7] VPWR VGND sg13g2_buf_1
XFILLER_8_373 VPWR VGND sg13g2_decap_8
Xoutput74 net74 S4BEG[10] VPWR VGND sg13g2_buf_1
Xoutput85 net85 S4BEG[6] VPWR VGND sg13g2_buf_1
Xoutput63 net63 S2BEG[6] VPWR VGND sg13g2_buf_1
Xoutput96 net96 SS4BEG[1] VPWR VGND sg13g2_buf_1
.ends

