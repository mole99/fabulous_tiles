magic
tech ihp-sg13g2
magscale 1 2
timestamp 1743692728
<< metal1 >>
rect 1152 9848 45216 9872
rect 1152 9808 3688 9848
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 4056 9808 18808 9848
rect 18848 9808 18890 9848
rect 18930 9808 18972 9848
rect 19012 9808 19054 9848
rect 19094 9808 19136 9848
rect 19176 9808 33928 9848
rect 33968 9808 34010 9848
rect 34050 9808 34092 9848
rect 34132 9808 34174 9848
rect 34214 9808 34256 9848
rect 34296 9808 45216 9848
rect 1152 9784 45216 9808
rect 10971 9680 11013 9689
rect 10971 9640 10972 9680
rect 11012 9640 11013 9680
rect 10971 9631 11013 9640
rect 11355 9680 11397 9689
rect 11355 9640 11356 9680
rect 11396 9640 11397 9680
rect 11355 9631 11397 9640
rect 11739 9680 11781 9689
rect 11739 9640 11740 9680
rect 11780 9640 11781 9680
rect 11739 9631 11781 9640
rect 12123 9680 12165 9689
rect 12123 9640 12124 9680
rect 12164 9640 12165 9680
rect 12123 9631 12165 9640
rect 12507 9680 12549 9689
rect 12507 9640 12508 9680
rect 12548 9640 12549 9680
rect 12507 9631 12549 9640
rect 12891 9680 12933 9689
rect 12891 9640 12892 9680
rect 12932 9640 12933 9680
rect 12891 9631 12933 9640
rect 13275 9680 13317 9689
rect 13275 9640 13276 9680
rect 13316 9640 13317 9680
rect 13275 9631 13317 9640
rect 13659 9680 13701 9689
rect 13659 9640 13660 9680
rect 13700 9640 13701 9680
rect 13659 9631 13701 9640
rect 14043 9680 14085 9689
rect 14043 9640 14044 9680
rect 14084 9640 14085 9680
rect 14043 9631 14085 9640
rect 14427 9680 14469 9689
rect 14427 9640 14428 9680
rect 14468 9640 14469 9680
rect 14427 9631 14469 9640
rect 14811 9680 14853 9689
rect 14811 9640 14812 9680
rect 14852 9640 14853 9680
rect 14811 9631 14853 9640
rect 15195 9680 15237 9689
rect 15195 9640 15196 9680
rect 15236 9640 15237 9680
rect 15195 9631 15237 9640
rect 15579 9680 15621 9689
rect 15579 9640 15580 9680
rect 15620 9640 15621 9680
rect 15579 9631 15621 9640
rect 15963 9680 16005 9689
rect 15963 9640 15964 9680
rect 16004 9640 16005 9680
rect 15963 9631 16005 9640
rect 16347 9680 16389 9689
rect 16347 9640 16348 9680
rect 16388 9640 16389 9680
rect 16347 9631 16389 9640
rect 16731 9680 16773 9689
rect 16731 9640 16732 9680
rect 16772 9640 16773 9680
rect 16731 9631 16773 9640
rect 17115 9680 17157 9689
rect 17115 9640 17116 9680
rect 17156 9640 17157 9680
rect 17115 9631 17157 9640
rect 17499 9680 17541 9689
rect 17499 9640 17500 9680
rect 17540 9640 17541 9680
rect 17499 9631 17541 9640
rect 17883 9680 17925 9689
rect 17883 9640 17884 9680
rect 17924 9640 17925 9680
rect 17883 9631 17925 9640
rect 18267 9680 18309 9689
rect 18267 9640 18268 9680
rect 18308 9640 18309 9680
rect 18267 9631 18309 9640
rect 18651 9680 18693 9689
rect 18651 9640 18652 9680
rect 18692 9640 18693 9680
rect 18651 9631 18693 9640
rect 19035 9680 19077 9689
rect 19035 9640 19036 9680
rect 19076 9640 19077 9680
rect 19035 9631 19077 9640
rect 20187 9680 20229 9689
rect 20187 9640 20188 9680
rect 20228 9640 20229 9680
rect 20187 9631 20229 9640
rect 20667 9680 20709 9689
rect 20667 9640 20668 9680
rect 20708 9640 20709 9680
rect 20667 9631 20709 9640
rect 21435 9680 21477 9689
rect 21435 9640 21436 9680
rect 21476 9640 21477 9680
rect 21435 9631 21477 9640
rect 31227 9680 31269 9689
rect 31227 9640 31228 9680
rect 31268 9640 31269 9680
rect 31227 9631 31269 9640
rect 31995 9680 32037 9689
rect 31995 9640 31996 9680
rect 32036 9640 32037 9680
rect 31995 9631 32037 9640
rect 32763 9680 32805 9689
rect 32763 9640 32764 9680
rect 32804 9640 32805 9680
rect 32763 9631 32805 9640
rect 33147 9680 33189 9689
rect 33147 9640 33148 9680
rect 33188 9640 33189 9680
rect 33147 9631 33189 9640
rect 34683 9680 34725 9689
rect 34683 9640 34684 9680
rect 34724 9640 34725 9680
rect 34683 9631 34725 9640
rect 36219 9680 36261 9689
rect 36219 9640 36220 9680
rect 36260 9640 36261 9680
rect 36219 9631 36261 9640
rect 43227 9680 43269 9689
rect 43227 9640 43228 9680
rect 43268 9640 43269 9680
rect 43227 9631 43269 9640
rect 43611 9680 43653 9689
rect 43611 9640 43612 9680
rect 43652 9640 43653 9680
rect 43611 9631 43653 9640
rect 43995 9680 44037 9689
rect 43995 9640 43996 9680
rect 44036 9640 44037 9680
rect 43995 9631 44037 9640
rect 19419 9596 19461 9605
rect 19419 9556 19420 9596
rect 19460 9556 19461 9596
rect 19419 9547 19461 9556
rect 20283 9596 20325 9605
rect 20283 9556 20284 9596
rect 20324 9556 20325 9596
rect 20283 9547 20325 9556
rect 31611 9596 31653 9605
rect 31611 9556 31612 9596
rect 31652 9556 31653 9596
rect 31611 9547 31653 9556
rect 32379 9596 32421 9605
rect 32379 9556 32380 9596
rect 32420 9556 32421 9596
rect 32379 9547 32421 9556
rect 36603 9596 36645 9605
rect 36603 9556 36604 9596
rect 36644 9556 36645 9596
rect 36603 9547 36645 9556
rect 10731 9512 10773 9521
rect 10731 9472 10732 9512
rect 10772 9472 10773 9512
rect 10731 9463 10773 9472
rect 11115 9512 11157 9521
rect 11115 9472 11116 9512
rect 11156 9472 11157 9512
rect 11115 9463 11157 9472
rect 11499 9512 11541 9521
rect 11499 9472 11500 9512
rect 11540 9472 11541 9512
rect 11499 9463 11541 9472
rect 11883 9512 11925 9521
rect 11883 9472 11884 9512
rect 11924 9472 11925 9512
rect 11883 9463 11925 9472
rect 12267 9512 12309 9521
rect 12267 9472 12268 9512
rect 12308 9472 12309 9512
rect 12267 9463 12309 9472
rect 12651 9512 12693 9521
rect 12651 9472 12652 9512
rect 12692 9472 12693 9512
rect 12651 9463 12693 9472
rect 13035 9512 13077 9521
rect 13035 9472 13036 9512
rect 13076 9472 13077 9512
rect 13035 9463 13077 9472
rect 13419 9512 13461 9521
rect 13419 9472 13420 9512
rect 13460 9472 13461 9512
rect 13419 9463 13461 9472
rect 13803 9512 13845 9521
rect 13803 9472 13804 9512
rect 13844 9472 13845 9512
rect 13803 9463 13845 9472
rect 14187 9512 14229 9521
rect 14187 9472 14188 9512
rect 14228 9472 14229 9512
rect 14187 9463 14229 9472
rect 14571 9512 14613 9521
rect 14571 9472 14572 9512
rect 14612 9472 14613 9512
rect 14571 9463 14613 9472
rect 14955 9512 14997 9521
rect 14955 9472 14956 9512
rect 14996 9472 14997 9512
rect 14955 9463 14997 9472
rect 15339 9512 15381 9521
rect 15339 9472 15340 9512
rect 15380 9472 15381 9512
rect 15339 9463 15381 9472
rect 15723 9512 15765 9521
rect 15723 9472 15724 9512
rect 15764 9472 15765 9512
rect 15723 9463 15765 9472
rect 16107 9512 16149 9521
rect 16107 9472 16108 9512
rect 16148 9472 16149 9512
rect 16107 9463 16149 9472
rect 16491 9512 16533 9521
rect 16491 9472 16492 9512
rect 16532 9472 16533 9512
rect 16491 9463 16533 9472
rect 16875 9512 16917 9521
rect 16875 9472 16876 9512
rect 16916 9472 16917 9512
rect 16875 9463 16917 9472
rect 17259 9512 17301 9521
rect 17259 9472 17260 9512
rect 17300 9472 17301 9512
rect 17259 9463 17301 9472
rect 17643 9512 17685 9521
rect 17643 9472 17644 9512
rect 17684 9472 17685 9512
rect 17643 9463 17685 9472
rect 18027 9512 18069 9521
rect 18027 9472 18028 9512
rect 18068 9472 18069 9512
rect 18027 9463 18069 9472
rect 18411 9512 18453 9521
rect 18411 9472 18412 9512
rect 18452 9472 18453 9512
rect 18411 9463 18453 9472
rect 18795 9512 18837 9521
rect 18795 9472 18796 9512
rect 18836 9472 18837 9512
rect 18795 9463 18837 9472
rect 19179 9512 19221 9521
rect 19179 9472 19180 9512
rect 19220 9472 19221 9512
rect 19179 9463 19221 9472
rect 19563 9512 19605 9521
rect 19563 9472 19564 9512
rect 19604 9472 19605 9512
rect 19563 9463 19605 9472
rect 19947 9512 19989 9521
rect 19947 9472 19948 9512
rect 19988 9472 19989 9512
rect 19947 9463 19989 9472
rect 20523 9512 20565 9521
rect 20523 9472 20524 9512
rect 20564 9472 20565 9512
rect 20523 9463 20565 9472
rect 20907 9512 20949 9521
rect 20907 9472 20908 9512
rect 20948 9472 20949 9512
rect 20907 9463 20949 9472
rect 21675 9512 21717 9521
rect 21675 9472 21676 9512
rect 21716 9472 21717 9512
rect 21675 9463 21717 9472
rect 31467 9512 31509 9521
rect 31467 9472 31468 9512
rect 31508 9472 31509 9512
rect 31467 9463 31509 9472
rect 31851 9512 31893 9521
rect 31851 9472 31852 9512
rect 31892 9472 31893 9512
rect 31851 9463 31893 9472
rect 32235 9512 32277 9521
rect 32235 9472 32236 9512
rect 32276 9472 32277 9512
rect 32235 9463 32277 9472
rect 32619 9512 32661 9521
rect 32619 9472 32620 9512
rect 32660 9472 32661 9512
rect 32619 9463 32661 9472
rect 33003 9512 33045 9521
rect 33003 9472 33004 9512
rect 33044 9472 33045 9512
rect 33003 9463 33045 9472
rect 33387 9512 33429 9521
rect 33387 9472 33388 9512
rect 33428 9472 33429 9512
rect 33387 9463 33429 9472
rect 33531 9512 33573 9521
rect 33531 9472 33532 9512
rect 33572 9472 33573 9512
rect 33531 9463 33573 9472
rect 33771 9512 33813 9521
rect 33771 9472 33772 9512
rect 33812 9472 33813 9512
rect 33771 9463 33813 9472
rect 34155 9512 34197 9521
rect 34155 9472 34156 9512
rect 34196 9472 34197 9512
rect 34155 9463 34197 9472
rect 34539 9512 34581 9521
rect 34539 9472 34540 9512
rect 34580 9472 34581 9512
rect 34539 9463 34581 9472
rect 34923 9512 34965 9521
rect 34923 9472 34924 9512
rect 34964 9472 34965 9512
rect 34923 9463 34965 9472
rect 35307 9512 35349 9521
rect 35307 9472 35308 9512
rect 35348 9472 35349 9512
rect 35307 9463 35349 9472
rect 35691 9512 35733 9521
rect 35691 9472 35692 9512
rect 35732 9472 35733 9512
rect 35691 9463 35733 9472
rect 36075 9512 36117 9521
rect 36075 9472 36076 9512
rect 36116 9472 36117 9512
rect 36075 9463 36117 9472
rect 36459 9512 36501 9521
rect 36459 9472 36460 9512
rect 36500 9472 36501 9512
rect 36459 9463 36501 9472
rect 36843 9512 36885 9521
rect 36843 9472 36844 9512
rect 36884 9472 36885 9512
rect 36843 9463 36885 9472
rect 37131 9512 37173 9521
rect 37131 9472 37132 9512
rect 37172 9472 37173 9512
rect 37131 9463 37173 9472
rect 37707 9512 37749 9521
rect 37707 9472 37708 9512
rect 37748 9472 37749 9512
rect 37707 9463 37749 9472
rect 37899 9512 37941 9521
rect 37899 9472 37900 9512
rect 37940 9472 37941 9512
rect 37899 9463 37941 9472
rect 38475 9512 38517 9521
rect 38475 9472 38476 9512
rect 38516 9472 38517 9512
rect 38475 9463 38517 9472
rect 39051 9512 39093 9521
rect 39051 9472 39052 9512
rect 39092 9472 39093 9512
rect 39051 9463 39093 9472
rect 39627 9512 39669 9521
rect 39627 9472 39628 9512
rect 39668 9472 39669 9512
rect 39627 9463 39669 9472
rect 39915 9512 39957 9521
rect 39915 9472 39916 9512
rect 39956 9472 39957 9512
rect 39915 9463 39957 9472
rect 40491 9512 40533 9521
rect 40491 9472 40492 9512
rect 40532 9472 40533 9512
rect 40491 9463 40533 9472
rect 40779 9512 40821 9521
rect 40779 9472 40780 9512
rect 40820 9472 40821 9512
rect 40779 9463 40821 9472
rect 42987 9512 43029 9521
rect 42987 9472 42988 9512
rect 43028 9472 43029 9512
rect 42987 9463 43029 9472
rect 43371 9512 43413 9521
rect 43371 9472 43372 9512
rect 43412 9472 43413 9512
rect 43371 9463 43413 9472
rect 43755 9512 43797 9521
rect 43755 9472 43756 9512
rect 43796 9472 43797 9512
rect 43755 9463 43797 9472
rect 44139 9512 44181 9521
rect 44139 9472 44140 9512
rect 44180 9472 44181 9512
rect 44139 9463 44181 9472
rect 44523 9512 44565 9521
rect 44523 9472 44524 9512
rect 44564 9472 44565 9512
rect 44523 9463 44565 9472
rect 44907 9512 44949 9521
rect 44907 9472 44908 9512
rect 44948 9472 44949 9512
rect 44907 9463 44949 9472
rect 19803 9344 19845 9353
rect 19803 9304 19804 9344
rect 19844 9304 19845 9344
rect 19803 9295 19845 9304
rect 34299 9344 34341 9353
rect 34299 9304 34300 9344
rect 34340 9304 34341 9344
rect 34299 9295 34341 9304
rect 35835 9344 35877 9353
rect 35835 9304 35836 9344
rect 35876 9304 35877 9344
rect 35835 9295 35877 9304
rect 44379 9344 44421 9353
rect 44379 9304 44380 9344
rect 44420 9304 44421 9344
rect 44379 9295 44421 9304
rect 21099 9260 21141 9269
rect 21099 9220 21100 9260
rect 21140 9220 21141 9260
rect 21099 9211 21141 9220
rect 33915 9260 33957 9269
rect 33915 9220 33916 9260
rect 33956 9220 33957 9260
rect 33915 9211 33957 9220
rect 35067 9260 35109 9269
rect 35067 9220 35068 9260
rect 35108 9220 35109 9260
rect 35067 9211 35109 9220
rect 35451 9260 35493 9269
rect 35451 9220 35452 9260
rect 35492 9220 35493 9260
rect 35451 9211 35493 9220
rect 37035 9260 37077 9269
rect 37035 9220 37036 9260
rect 37076 9220 37077 9260
rect 37035 9211 37077 9220
rect 37306 9260 37364 9261
rect 37306 9220 37315 9260
rect 37355 9220 37364 9260
rect 37306 9219 37364 9220
rect 37882 9260 37940 9261
rect 37882 9220 37891 9260
rect 37931 9220 37940 9260
rect 37882 9219 37940 9220
rect 38187 9260 38229 9269
rect 38187 9220 38188 9260
rect 38228 9220 38229 9260
rect 38187 9211 38229 9220
rect 38763 9260 38805 9269
rect 38763 9220 38764 9260
rect 38804 9220 38805 9260
rect 38763 9211 38805 9220
rect 39322 9260 39380 9261
rect 39322 9220 39331 9260
rect 39371 9220 39380 9260
rect 39322 9219 39380 9220
rect 40203 9260 40245 9269
rect 40203 9220 40204 9260
rect 40244 9220 40245 9260
rect 40203 9211 40245 9220
rect 44763 9260 44805 9269
rect 44763 9220 44764 9260
rect 44804 9220 44805 9260
rect 44763 9211 44805 9220
rect 45147 9260 45189 9269
rect 45147 9220 45148 9260
rect 45188 9220 45189 9260
rect 45147 9211 45189 9220
rect 1152 9092 45216 9116
rect 1152 9052 4928 9092
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 5296 9052 20048 9092
rect 20088 9052 20130 9092
rect 20170 9052 20212 9092
rect 20252 9052 20294 9092
rect 20334 9052 20376 9092
rect 20416 9052 35168 9092
rect 35208 9052 35250 9092
rect 35290 9052 35332 9092
rect 35372 9052 35414 9092
rect 35454 9052 35496 9092
rect 35536 9052 45216 9092
rect 1152 9028 45216 9052
rect 11067 8924 11109 8933
rect 11067 8884 11068 8924
rect 11108 8884 11109 8924
rect 11067 8875 11109 8884
rect 11451 8924 11493 8933
rect 11451 8884 11452 8924
rect 11492 8884 11493 8924
rect 11451 8875 11493 8884
rect 11835 8924 11877 8933
rect 11835 8884 11836 8924
rect 11876 8884 11877 8924
rect 11835 8875 11877 8884
rect 12219 8924 12261 8933
rect 12219 8884 12220 8924
rect 12260 8884 12261 8924
rect 12219 8875 12261 8884
rect 12603 8924 12645 8933
rect 12603 8884 12604 8924
rect 12644 8884 12645 8924
rect 12603 8875 12645 8884
rect 13371 8924 13413 8933
rect 13371 8884 13372 8924
rect 13412 8884 13413 8924
rect 13371 8875 13413 8884
rect 13755 8924 13797 8933
rect 13755 8884 13756 8924
rect 13796 8884 13797 8924
rect 13755 8875 13797 8884
rect 14139 8924 14181 8933
rect 14139 8884 14140 8924
rect 14180 8884 14181 8924
rect 14139 8875 14181 8884
rect 14523 8924 14565 8933
rect 14523 8884 14524 8924
rect 14564 8884 14565 8924
rect 14523 8875 14565 8884
rect 14907 8924 14949 8933
rect 14907 8884 14908 8924
rect 14948 8884 14949 8924
rect 14907 8875 14949 8884
rect 15291 8924 15333 8933
rect 15291 8884 15292 8924
rect 15332 8884 15333 8924
rect 15291 8875 15333 8884
rect 15675 8924 15717 8933
rect 15675 8884 15676 8924
rect 15716 8884 15717 8924
rect 15675 8875 15717 8884
rect 16059 8924 16101 8933
rect 16059 8884 16060 8924
rect 16100 8884 16101 8924
rect 16059 8875 16101 8884
rect 16443 8924 16485 8933
rect 16443 8884 16444 8924
rect 16484 8884 16485 8924
rect 16443 8875 16485 8884
rect 16827 8924 16869 8933
rect 16827 8884 16828 8924
rect 16868 8884 16869 8924
rect 16827 8875 16869 8884
rect 17211 8924 17253 8933
rect 17211 8884 17212 8924
rect 17252 8884 17253 8924
rect 17211 8875 17253 8884
rect 17595 8924 17637 8933
rect 17595 8884 17596 8924
rect 17636 8884 17637 8924
rect 17595 8875 17637 8884
rect 17979 8924 18021 8933
rect 17979 8884 17980 8924
rect 18020 8884 18021 8924
rect 17979 8875 18021 8884
rect 18363 8924 18405 8933
rect 18363 8884 18364 8924
rect 18404 8884 18405 8924
rect 18363 8875 18405 8884
rect 18747 8924 18789 8933
rect 18747 8884 18748 8924
rect 18788 8884 18789 8924
rect 18747 8875 18789 8884
rect 19131 8924 19173 8933
rect 19131 8884 19132 8924
rect 19172 8884 19173 8924
rect 19131 8875 19173 8884
rect 19515 8924 19557 8933
rect 19515 8884 19516 8924
rect 19556 8884 19557 8924
rect 19515 8875 19557 8884
rect 19899 8924 19941 8933
rect 19899 8884 19900 8924
rect 19940 8884 19941 8924
rect 19899 8875 19941 8884
rect 27195 8924 27237 8933
rect 27195 8884 27196 8924
rect 27236 8884 27237 8924
rect 27195 8875 27237 8884
rect 27579 8924 27621 8933
rect 27579 8884 27580 8924
rect 27620 8884 27621 8924
rect 27579 8875 27621 8884
rect 32187 8924 32229 8933
rect 32187 8884 32188 8924
rect 32228 8884 32229 8924
rect 32187 8875 32229 8884
rect 32571 8924 32613 8933
rect 32571 8884 32572 8924
rect 32612 8884 32613 8924
rect 32571 8875 32613 8884
rect 32955 8924 32997 8933
rect 32955 8884 32956 8924
rect 32996 8884 32997 8924
rect 32955 8875 32997 8884
rect 33339 8924 33381 8933
rect 33339 8884 33340 8924
rect 33380 8884 33381 8924
rect 33339 8875 33381 8884
rect 34234 8924 34292 8925
rect 34234 8884 34243 8924
rect 34283 8884 34292 8924
rect 34234 8883 34292 8884
rect 34875 8924 34917 8933
rect 34875 8884 34876 8924
rect 34916 8884 34917 8924
rect 34875 8875 34917 8884
rect 37210 8924 37268 8925
rect 37210 8884 37219 8924
rect 37259 8884 37268 8924
rect 37210 8883 37268 8884
rect 37755 8924 37797 8933
rect 37755 8884 37756 8924
rect 37796 8884 37797 8924
rect 37755 8875 37797 8884
rect 39994 8924 40052 8925
rect 39994 8884 40003 8924
rect 40043 8884 40052 8924
rect 39994 8883 40052 8884
rect 43995 8924 44037 8933
rect 43995 8884 43996 8924
rect 44036 8884 44037 8924
rect 43995 8875 44037 8884
rect 44379 8924 44421 8933
rect 44379 8884 44380 8924
rect 44420 8884 44421 8924
rect 44379 8875 44421 8884
rect 25851 8840 25893 8849
rect 25851 8800 25852 8840
rect 25892 8800 25893 8840
rect 25851 8791 25893 8800
rect 26427 8840 26469 8849
rect 26427 8800 26428 8840
rect 26468 8800 26469 8840
rect 26427 8791 26469 8800
rect 27963 8840 28005 8849
rect 27963 8800 27964 8840
rect 28004 8800 28005 8840
rect 27963 8791 28005 8800
rect 32091 8840 32133 8849
rect 32091 8800 32092 8840
rect 32132 8800 32133 8840
rect 32091 8791 32133 8800
rect 35259 8840 35301 8849
rect 35259 8800 35260 8840
rect 35300 8800 35301 8840
rect 35259 8791 35301 8800
rect 36315 8840 36357 8849
rect 36315 8800 36316 8840
rect 36356 8800 36357 8840
rect 36315 8791 36357 8800
rect 36699 8840 36741 8849
rect 36699 8800 36700 8840
rect 36740 8800 36741 8840
rect 36699 8791 36741 8800
rect 38139 8840 38181 8849
rect 38139 8800 38140 8840
rect 38180 8800 38181 8840
rect 38139 8791 38181 8800
rect 11242 8672 11300 8673
rect 11242 8632 11251 8672
rect 11291 8632 11300 8672
rect 11242 8631 11300 8632
rect 11691 8672 11733 8681
rect 11691 8632 11692 8672
rect 11732 8632 11733 8672
rect 11691 8623 11733 8632
rect 12075 8672 12117 8681
rect 12075 8632 12076 8672
rect 12116 8632 12117 8672
rect 12075 8623 12117 8632
rect 12459 8672 12501 8681
rect 12459 8632 12460 8672
rect 12500 8632 12501 8672
rect 12459 8623 12501 8632
rect 12843 8672 12885 8681
rect 12843 8632 12844 8672
rect 12884 8632 12885 8672
rect 12843 8623 12885 8632
rect 13227 8672 13269 8681
rect 13227 8632 13228 8672
rect 13268 8632 13269 8672
rect 13227 8623 13269 8632
rect 13611 8672 13653 8681
rect 13611 8632 13612 8672
rect 13652 8632 13653 8672
rect 13611 8623 13653 8632
rect 13995 8672 14037 8681
rect 13995 8632 13996 8672
rect 14036 8632 14037 8672
rect 13995 8623 14037 8632
rect 14379 8672 14421 8681
rect 14379 8632 14380 8672
rect 14420 8632 14421 8672
rect 14379 8623 14421 8632
rect 14763 8672 14805 8681
rect 14763 8632 14764 8672
rect 14804 8632 14805 8672
rect 14763 8623 14805 8632
rect 15147 8672 15189 8681
rect 15147 8632 15148 8672
rect 15188 8632 15189 8672
rect 15147 8623 15189 8632
rect 15531 8672 15573 8681
rect 15531 8632 15532 8672
rect 15572 8632 15573 8672
rect 15531 8623 15573 8632
rect 15915 8672 15957 8681
rect 15915 8632 15916 8672
rect 15956 8632 15957 8672
rect 15915 8623 15957 8632
rect 16299 8672 16341 8681
rect 16299 8632 16300 8672
rect 16340 8632 16341 8672
rect 16299 8623 16341 8632
rect 16683 8672 16725 8681
rect 16683 8632 16684 8672
rect 16724 8632 16725 8672
rect 16683 8623 16725 8632
rect 17067 8672 17109 8681
rect 17067 8632 17068 8672
rect 17108 8632 17109 8672
rect 17067 8623 17109 8632
rect 17451 8672 17493 8681
rect 17451 8632 17452 8672
rect 17492 8632 17493 8672
rect 17451 8623 17493 8632
rect 17835 8672 17877 8681
rect 17835 8632 17836 8672
rect 17876 8632 17877 8672
rect 17835 8623 17877 8632
rect 18219 8672 18261 8681
rect 18219 8632 18220 8672
rect 18260 8632 18261 8672
rect 18219 8623 18261 8632
rect 18603 8672 18645 8681
rect 18603 8632 18604 8672
rect 18644 8632 18645 8672
rect 18603 8623 18645 8632
rect 18987 8672 19029 8681
rect 18987 8632 18988 8672
rect 19028 8632 19029 8672
rect 18987 8623 19029 8632
rect 19371 8672 19413 8681
rect 19371 8632 19372 8672
rect 19412 8632 19413 8672
rect 19371 8623 19413 8632
rect 19755 8672 19797 8681
rect 19755 8632 19756 8672
rect 19796 8632 19797 8672
rect 19755 8623 19797 8632
rect 20139 8672 20181 8681
rect 20139 8632 20140 8672
rect 20180 8632 20181 8672
rect 20139 8623 20181 8632
rect 26091 8672 26133 8681
rect 26091 8632 26092 8672
rect 26132 8632 26133 8672
rect 26091 8623 26133 8632
rect 26667 8672 26709 8681
rect 26667 8632 26668 8672
rect 26708 8632 26709 8672
rect 26667 8623 26709 8632
rect 27435 8672 27477 8681
rect 27435 8632 27436 8672
rect 27476 8632 27477 8672
rect 27435 8623 27477 8632
rect 27819 8672 27861 8681
rect 27819 8632 27820 8672
rect 27860 8632 27861 8672
rect 27819 8623 27861 8632
rect 28203 8672 28245 8681
rect 28203 8632 28204 8672
rect 28244 8632 28245 8672
rect 28203 8623 28245 8632
rect 28347 8672 28389 8681
rect 28347 8632 28348 8672
rect 28388 8632 28389 8672
rect 28347 8623 28389 8632
rect 28587 8672 28629 8681
rect 28587 8632 28588 8672
rect 28628 8632 28629 8672
rect 28587 8623 28629 8632
rect 28731 8672 28773 8681
rect 28731 8632 28732 8672
rect 28772 8632 28773 8672
rect 28731 8623 28773 8632
rect 28971 8672 29013 8681
rect 28971 8632 28972 8672
rect 29012 8632 29013 8672
rect 28971 8623 29013 8632
rect 31851 8672 31893 8681
rect 31851 8632 31852 8672
rect 31892 8632 31893 8672
rect 31851 8623 31893 8632
rect 32427 8672 32469 8681
rect 32427 8632 32428 8672
rect 32468 8632 32469 8672
rect 32427 8623 32469 8632
rect 32811 8672 32853 8681
rect 32811 8632 32812 8672
rect 32852 8632 32853 8672
rect 32811 8623 32853 8632
rect 33195 8672 33237 8681
rect 33195 8632 33196 8672
rect 33236 8632 33237 8672
rect 33195 8623 33237 8632
rect 33579 8672 33621 8681
rect 33579 8632 33580 8672
rect 33620 8632 33621 8672
rect 33579 8623 33621 8632
rect 33867 8672 33909 8681
rect 33867 8632 33868 8672
rect 33908 8632 33909 8672
rect 33867 8623 33909 8632
rect 34251 8672 34293 8681
rect 34251 8632 34252 8672
rect 34292 8632 34293 8672
rect 34251 8623 34293 8632
rect 34539 8672 34581 8681
rect 34539 8632 34540 8672
rect 34580 8632 34581 8672
rect 34539 8623 34581 8632
rect 35115 8672 35157 8681
rect 35115 8632 35116 8672
rect 35156 8632 35157 8672
rect 35115 8623 35157 8632
rect 35499 8672 35541 8681
rect 35499 8632 35500 8672
rect 35540 8632 35541 8672
rect 35499 8623 35541 8632
rect 35787 8672 35829 8681
rect 35787 8632 35788 8672
rect 35828 8632 35829 8672
rect 35787 8623 35829 8632
rect 36075 8672 36117 8681
rect 36075 8632 36076 8672
rect 36116 8632 36117 8672
rect 36075 8623 36117 8632
rect 36459 8672 36501 8681
rect 36459 8632 36460 8672
rect 36500 8632 36501 8672
rect 36459 8623 36501 8632
rect 36843 8672 36885 8681
rect 36843 8632 36844 8672
rect 36884 8632 36885 8672
rect 36843 8623 36885 8632
rect 37227 8672 37269 8681
rect 37227 8632 37228 8672
rect 37268 8632 37269 8672
rect 37227 8623 37269 8632
rect 37515 8672 37557 8681
rect 37515 8632 37516 8672
rect 37556 8632 37557 8672
rect 37515 8623 37557 8632
rect 37899 8672 37941 8681
rect 37899 8632 37900 8672
rect 37940 8632 37941 8672
rect 37899 8623 37941 8632
rect 38283 8672 38325 8681
rect 38283 8632 38284 8672
rect 38324 8632 38325 8672
rect 38283 8623 38325 8632
rect 38571 8672 38613 8681
rect 38571 8632 38572 8672
rect 38612 8632 38613 8672
rect 38571 8623 38613 8632
rect 38859 8672 38901 8681
rect 38859 8632 38860 8672
rect 38900 8632 38901 8672
rect 38859 8623 38901 8632
rect 39147 8672 39189 8681
rect 39147 8632 39148 8672
rect 39188 8632 39189 8672
rect 39147 8623 39189 8632
rect 39435 8672 39477 8681
rect 39435 8632 39436 8672
rect 39476 8632 39477 8672
rect 39435 8623 39477 8632
rect 39723 8672 39765 8681
rect 39723 8632 39724 8672
rect 39764 8632 39765 8672
rect 39723 8623 39765 8632
rect 40299 8672 40341 8681
rect 40299 8632 40300 8672
rect 40340 8632 40341 8672
rect 40299 8623 40341 8632
rect 43755 8672 43797 8681
rect 43755 8632 43756 8672
rect 43796 8632 43797 8672
rect 43755 8623 43797 8632
rect 44139 8672 44181 8681
rect 44139 8632 44140 8672
rect 44180 8632 44181 8672
rect 44139 8623 44181 8632
rect 44523 8672 44565 8681
rect 44523 8632 44524 8672
rect 44564 8632 44565 8672
rect 44523 8623 44565 8632
rect 44907 8672 44949 8681
rect 44907 8632 44908 8672
rect 44948 8632 44949 8672
rect 44907 8623 44949 8632
rect 12987 8588 13029 8597
rect 12987 8548 12988 8588
rect 13028 8548 13029 8588
rect 12987 8539 13029 8548
rect 34779 8588 34821 8597
rect 34779 8548 34780 8588
rect 34820 8548 34821 8588
rect 34779 8539 34821 8548
rect 34107 8504 34149 8513
rect 34107 8464 34108 8504
rect 34148 8464 34149 8504
rect 34107 8455 34149 8464
rect 44763 8504 44805 8513
rect 44763 8464 44764 8504
rect 44804 8464 44805 8504
rect 44763 8455 44805 8464
rect 45147 8504 45189 8513
rect 45147 8464 45148 8504
rect 45188 8464 45189 8504
rect 45147 8455 45189 8464
rect 1152 8336 45216 8360
rect 1152 8296 3688 8336
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 4056 8296 18808 8336
rect 18848 8296 18890 8336
rect 18930 8296 18972 8336
rect 19012 8296 19054 8336
rect 19094 8296 19136 8336
rect 19176 8296 33928 8336
rect 33968 8296 34010 8336
rect 34050 8296 34092 8336
rect 34132 8296 34174 8336
rect 34214 8296 34256 8336
rect 34296 8296 45216 8336
rect 1152 8272 45216 8296
rect 25563 8168 25605 8177
rect 25563 8128 25564 8168
rect 25604 8128 25605 8168
rect 25563 8119 25605 8128
rect 25947 8168 25989 8177
rect 25947 8128 25948 8168
rect 25988 8128 25989 8168
rect 25947 8119 25989 8128
rect 26715 8168 26757 8177
rect 26715 8128 26716 8168
rect 26756 8128 26757 8168
rect 26715 8119 26757 8128
rect 27099 8168 27141 8177
rect 27099 8128 27100 8168
rect 27140 8128 27141 8168
rect 27099 8119 27141 8128
rect 32955 8168 32997 8177
rect 32955 8128 32956 8168
rect 32996 8128 32997 8168
rect 32955 8119 32997 8128
rect 39771 8168 39813 8177
rect 39771 8128 39772 8168
rect 39812 8128 39813 8168
rect 39771 8119 39813 8128
rect 43131 8168 43173 8177
rect 43131 8128 43132 8168
rect 43172 8128 43173 8168
rect 43131 8119 43173 8128
rect 26331 8084 26373 8093
rect 26331 8044 26332 8084
rect 26372 8044 26373 8084
rect 26331 8035 26373 8044
rect 25179 8000 25221 8009
rect 25179 7960 25180 8000
rect 25220 7960 25221 8000
rect 25179 7951 25221 7960
rect 25419 8000 25461 8009
rect 25419 7960 25420 8000
rect 25460 7960 25461 8000
rect 25419 7951 25461 7960
rect 25803 8000 25845 8009
rect 25803 7960 25804 8000
rect 25844 7960 25845 8000
rect 25803 7951 25845 7960
rect 26187 8000 26229 8009
rect 26187 7960 26188 8000
rect 26228 7960 26229 8000
rect 26187 7951 26229 7960
rect 26571 8000 26613 8009
rect 26571 7960 26572 8000
rect 26612 7960 26613 8000
rect 26571 7951 26613 7960
rect 26955 8000 26997 8009
rect 26955 7960 26956 8000
rect 26996 7960 26997 8000
rect 26955 7951 26997 7960
rect 27339 8000 27381 8009
rect 27339 7960 27340 8000
rect 27380 7960 27381 8000
rect 27339 7951 27381 7960
rect 27483 8000 27525 8009
rect 27483 7960 27484 8000
rect 27524 7960 27525 8000
rect 27483 7951 27525 7960
rect 27723 8000 27765 8009
rect 27723 7960 27724 8000
rect 27764 7960 27765 8000
rect 27723 7951 27765 7960
rect 28203 8000 28245 8009
rect 28203 7960 28204 8000
rect 28244 7960 28245 8000
rect 28203 7951 28245 7960
rect 32715 8000 32757 8009
rect 32715 7960 32716 8000
rect 32756 7960 32757 8000
rect 32715 7951 32757 7960
rect 34347 8000 34389 8009
rect 34347 7960 34348 8000
rect 34388 7960 34389 8000
rect 34347 7951 34389 7960
rect 34635 8000 34677 8009
rect 34635 7960 34636 8000
rect 34676 7960 34677 8000
rect 34635 7951 34677 7960
rect 34923 8000 34965 8009
rect 34923 7960 34924 8000
rect 34964 7960 34965 8000
rect 34923 7951 34965 7960
rect 35211 8000 35253 8009
rect 35211 7960 35212 8000
rect 35252 7960 35253 8000
rect 35211 7951 35253 7960
rect 35499 8000 35541 8009
rect 35499 7960 35500 8000
rect 35540 7960 35541 8000
rect 35499 7951 35541 7960
rect 35787 8000 35829 8009
rect 35787 7960 35788 8000
rect 35828 7960 35829 8000
rect 35787 7951 35829 7960
rect 36075 8000 36117 8009
rect 36075 7960 36076 8000
rect 36116 7960 36117 8000
rect 36075 7951 36117 7960
rect 36459 8000 36501 8009
rect 36459 7960 36460 8000
rect 36500 7960 36501 8000
rect 36459 7951 36501 7960
rect 36699 8000 36741 8009
rect 36699 7960 36700 8000
rect 36740 7960 36741 8000
rect 36699 7951 36741 7960
rect 38379 8000 38421 8009
rect 38379 7960 38380 8000
rect 38420 7960 38421 8000
rect 38379 7951 38421 7960
rect 38667 8000 38709 8009
rect 38667 7960 38668 8000
rect 38708 7960 38709 8000
rect 38667 7951 38709 7960
rect 39531 8000 39573 8009
rect 39531 7960 39532 8000
rect 39572 7960 39573 8000
rect 39531 7951 39573 7960
rect 43371 8000 43413 8009
rect 43371 7960 43372 8000
rect 43412 7960 43413 8000
rect 43371 7951 43413 7960
rect 44523 8000 44565 8009
rect 44523 7960 44524 8000
rect 44564 7960 44565 8000
rect 44523 7951 44565 7960
rect 44907 8000 44949 8009
rect 44907 7960 44908 8000
rect 44948 7960 44949 8000
rect 44907 7951 44949 7960
rect 36939 7916 36981 7925
rect 36939 7876 36940 7916
rect 36980 7876 36981 7916
rect 36939 7867 36981 7876
rect 37131 7916 37173 7925
rect 37131 7876 37132 7916
rect 37172 7876 37173 7916
rect 37131 7867 37173 7876
rect 27963 7748 28005 7757
rect 27963 7708 27964 7748
rect 28004 7708 28005 7748
rect 27963 7699 28005 7708
rect 37402 7748 37460 7749
rect 37402 7708 37411 7748
rect 37451 7708 37460 7748
rect 37402 7707 37460 7708
rect 37690 7748 37748 7749
rect 37690 7708 37699 7748
rect 37739 7708 37748 7748
rect 37690 7707 37748 7708
rect 37978 7748 38036 7749
rect 37978 7708 37987 7748
rect 38027 7708 38036 7748
rect 37978 7707 38036 7708
rect 44763 7748 44805 7757
rect 44763 7708 44764 7748
rect 44804 7708 44805 7748
rect 44763 7699 44805 7708
rect 45147 7748 45189 7757
rect 45147 7708 45148 7748
rect 45188 7708 45189 7748
rect 45147 7699 45189 7708
rect 1152 7580 45216 7604
rect 1152 7540 4928 7580
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 5296 7540 20048 7580
rect 20088 7540 20130 7580
rect 20170 7540 20212 7580
rect 20252 7540 20294 7580
rect 20334 7540 20376 7580
rect 20416 7540 35168 7580
rect 35208 7540 35250 7580
rect 35290 7540 35332 7580
rect 35372 7540 35414 7580
rect 35454 7540 35496 7580
rect 35536 7540 45216 7580
rect 1152 7516 45216 7540
rect 36075 7412 36117 7421
rect 36075 7372 36076 7412
rect 36116 7372 36117 7412
rect 36075 7363 36117 7372
rect 8331 7160 8373 7169
rect 8331 7120 8332 7160
rect 8372 7120 8373 7160
rect 8331 7111 8373 7120
rect 25899 7160 25941 7169
rect 25899 7120 25900 7160
rect 25940 7120 25941 7160
rect 25899 7111 25941 7120
rect 33291 7160 33333 7169
rect 33291 7120 33292 7160
rect 33332 7120 33333 7160
rect 33291 7111 33333 7120
rect 35691 7160 35733 7169
rect 35691 7120 35692 7160
rect 35732 7120 35733 7160
rect 35691 7111 35733 7120
rect 35931 7160 35973 7169
rect 35931 7120 35932 7160
rect 35972 7120 35973 7160
rect 35931 7111 35973 7120
rect 44523 7160 44565 7169
rect 44523 7120 44524 7160
rect 44564 7120 44565 7160
rect 44523 7111 44565 7120
rect 44907 7160 44949 7169
rect 44907 7120 44908 7160
rect 44948 7120 44949 7160
rect 44907 7111 44949 7120
rect 8571 7076 8613 7085
rect 8571 7036 8572 7076
rect 8612 7036 8613 7076
rect 8571 7027 8613 7036
rect 33531 7076 33573 7085
rect 33531 7036 33532 7076
rect 33572 7036 33573 7076
rect 33531 7027 33573 7036
rect 25659 6992 25701 7001
rect 25659 6952 25660 6992
rect 25700 6952 25701 6992
rect 25659 6943 25701 6952
rect 44763 6992 44805 7001
rect 44763 6952 44764 6992
rect 44804 6952 44805 6992
rect 44763 6943 44805 6952
rect 45147 6992 45189 7001
rect 45147 6952 45148 6992
rect 45188 6952 45189 6992
rect 45147 6943 45189 6952
rect 1152 6824 45216 6848
rect 1152 6784 3688 6824
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 4056 6784 18808 6824
rect 18848 6784 18890 6824
rect 18930 6784 18972 6824
rect 19012 6784 19054 6824
rect 19094 6784 19136 6824
rect 19176 6784 33928 6824
rect 33968 6784 34010 6824
rect 34050 6784 34092 6824
rect 34132 6784 34174 6824
rect 34214 6784 34256 6824
rect 34296 6784 45216 6824
rect 1152 6760 45216 6784
rect 7611 6656 7653 6665
rect 7611 6616 7612 6656
rect 7652 6616 7653 6656
rect 7611 6607 7653 6616
rect 8667 6572 8709 6581
rect 8667 6532 8668 6572
rect 8708 6532 8709 6572
rect 8667 6523 8709 6532
rect 9051 6572 9093 6581
rect 9051 6532 9052 6572
rect 9092 6532 9093 6572
rect 9051 6523 9093 6532
rect 9435 6572 9477 6581
rect 9435 6532 9436 6572
rect 9476 6532 9477 6572
rect 9435 6523 9477 6532
rect 13947 6572 13989 6581
rect 13947 6532 13948 6572
rect 13988 6532 13989 6572
rect 13947 6523 13989 6532
rect 19131 6572 19173 6581
rect 19131 6532 19132 6572
rect 19172 6532 19173 6572
rect 19131 6523 19173 6532
rect 7371 6488 7413 6497
rect 7371 6448 7372 6488
rect 7412 6448 7413 6488
rect 7371 6439 7413 6448
rect 7755 6488 7797 6497
rect 7755 6448 7756 6488
rect 7796 6448 7797 6488
rect 7755 6439 7797 6448
rect 8427 6488 8469 6497
rect 8427 6448 8428 6488
rect 8468 6448 8469 6488
rect 8427 6439 8469 6448
rect 8811 6488 8853 6497
rect 8811 6448 8812 6488
rect 8852 6448 8853 6488
rect 8811 6439 8853 6448
rect 9195 6488 9237 6497
rect 9195 6448 9196 6488
rect 9236 6448 9237 6488
rect 9195 6439 9237 6448
rect 13707 6488 13749 6497
rect 13707 6448 13708 6488
rect 13748 6448 13749 6488
rect 13707 6439 13749 6448
rect 19371 6488 19413 6497
rect 19371 6448 19372 6488
rect 19412 6448 19413 6488
rect 19371 6439 19413 6448
rect 19803 6488 19845 6497
rect 19803 6448 19804 6488
rect 19844 6448 19845 6488
rect 19803 6439 19845 6448
rect 20043 6488 20085 6497
rect 20043 6448 20044 6488
rect 20084 6448 20085 6488
rect 20043 6439 20085 6448
rect 20427 6488 20469 6497
rect 20427 6448 20428 6488
rect 20468 6448 20469 6488
rect 20427 6439 20469 6448
rect 33771 6488 33813 6497
rect 33771 6448 33772 6488
rect 33812 6448 33813 6488
rect 33771 6439 33813 6448
rect 35787 6488 35829 6497
rect 35787 6448 35788 6488
rect 35828 6448 35829 6488
rect 35787 6439 35829 6448
rect 35979 6488 36021 6497
rect 35979 6448 35980 6488
rect 36020 6448 36021 6488
rect 35979 6439 36021 6448
rect 44523 6488 44565 6497
rect 44523 6448 44524 6488
rect 44564 6448 44565 6488
rect 44523 6439 44565 6448
rect 44907 6488 44949 6497
rect 44907 6448 44908 6488
rect 44948 6448 44949 6488
rect 44907 6439 44949 6448
rect 7995 6320 8037 6329
rect 7995 6280 7996 6320
rect 8036 6280 8037 6320
rect 7995 6271 8037 6280
rect 45147 6320 45189 6329
rect 45147 6280 45148 6320
rect 45188 6280 45189 6320
rect 45147 6271 45189 6280
rect 20187 6236 20229 6245
rect 20187 6196 20188 6236
rect 20228 6196 20229 6236
rect 20187 6187 20229 6196
rect 34011 6236 34053 6245
rect 34011 6196 34012 6236
rect 34052 6196 34053 6236
rect 34011 6187 34053 6196
rect 44763 6236 44805 6245
rect 44763 6196 44764 6236
rect 44804 6196 44805 6236
rect 44763 6187 44805 6196
rect 1152 6068 45216 6092
rect 1152 6028 4928 6068
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 5296 6028 20048 6068
rect 20088 6028 20130 6068
rect 20170 6028 20212 6068
rect 20252 6028 20294 6068
rect 20334 6028 20376 6068
rect 20416 6028 35168 6068
rect 35208 6028 35250 6068
rect 35290 6028 35332 6068
rect 35372 6028 35414 6068
rect 35454 6028 35496 6068
rect 35536 6028 45216 6068
rect 1152 6004 45216 6028
rect 18267 5816 18309 5825
rect 18267 5776 18268 5816
rect 18308 5776 18309 5816
rect 18267 5767 18309 5776
rect 18651 5816 18693 5825
rect 18651 5776 18652 5816
rect 18692 5776 18693 5816
rect 18651 5767 18693 5776
rect 19035 5816 19077 5825
rect 19035 5776 19036 5816
rect 19076 5776 19077 5816
rect 19035 5767 19077 5776
rect 9099 5648 9141 5657
rect 9099 5608 9100 5648
rect 9140 5608 9141 5648
rect 9099 5599 9141 5608
rect 9483 5648 9525 5657
rect 9483 5608 9484 5648
rect 9524 5608 9525 5648
rect 9483 5599 9525 5608
rect 9867 5648 9909 5657
rect 9867 5608 9868 5648
rect 9908 5608 9909 5648
rect 9867 5599 9909 5608
rect 10251 5648 10293 5657
rect 10251 5608 10252 5648
rect 10292 5608 10293 5648
rect 10251 5599 10293 5608
rect 10635 5648 10677 5657
rect 10635 5608 10636 5648
rect 10676 5608 10677 5648
rect 10635 5599 10677 5608
rect 11019 5648 11061 5657
rect 11019 5608 11020 5648
rect 11060 5608 11061 5648
rect 11019 5599 11061 5608
rect 11355 5648 11397 5657
rect 11355 5608 11356 5648
rect 11396 5608 11397 5648
rect 11355 5599 11397 5608
rect 11595 5648 11637 5657
rect 11595 5608 11596 5648
rect 11636 5608 11637 5648
rect 11595 5599 11637 5608
rect 11818 5648 11876 5649
rect 11818 5608 11827 5648
rect 11867 5608 11876 5648
rect 11818 5607 11876 5608
rect 13227 5648 13269 5657
rect 13227 5608 13228 5648
rect 13268 5608 13269 5648
rect 13227 5599 13269 5608
rect 13563 5648 13605 5657
rect 13563 5608 13564 5648
rect 13604 5608 13605 5648
rect 13563 5599 13605 5608
rect 13803 5648 13845 5657
rect 13803 5608 13804 5648
rect 13844 5608 13845 5648
rect 13803 5599 13845 5608
rect 13995 5648 14037 5657
rect 13995 5608 13996 5648
rect 14036 5608 14037 5648
rect 13995 5599 14037 5608
rect 14235 5648 14277 5657
rect 14235 5608 14236 5648
rect 14276 5608 14277 5648
rect 14235 5599 14277 5608
rect 14571 5648 14613 5657
rect 14571 5608 14572 5648
rect 14612 5608 14613 5648
rect 14571 5599 14613 5608
rect 14955 5648 14997 5657
rect 14955 5608 14956 5648
rect 14996 5608 14997 5648
rect 14955 5599 14997 5608
rect 15099 5648 15141 5657
rect 15099 5608 15100 5648
rect 15140 5608 15141 5648
rect 15099 5599 15141 5608
rect 15339 5648 15381 5657
rect 15339 5608 15340 5648
rect 15380 5608 15381 5648
rect 15339 5599 15381 5608
rect 17883 5648 17925 5657
rect 17883 5608 17884 5648
rect 17924 5608 17925 5648
rect 17883 5599 17925 5608
rect 18123 5648 18165 5657
rect 18123 5608 18124 5648
rect 18164 5608 18165 5648
rect 18123 5599 18165 5608
rect 18507 5648 18549 5657
rect 18507 5608 18508 5648
rect 18548 5608 18549 5648
rect 18507 5599 18549 5608
rect 18891 5648 18933 5657
rect 18891 5608 18892 5648
rect 18932 5608 18933 5648
rect 18891 5599 18933 5608
rect 19275 5648 19317 5657
rect 19275 5608 19276 5648
rect 19316 5608 19317 5648
rect 19275 5599 19317 5608
rect 19659 5648 19701 5657
rect 19659 5608 19660 5648
rect 19700 5608 19701 5648
rect 19659 5599 19701 5608
rect 20043 5648 20085 5657
rect 20043 5608 20044 5648
rect 20084 5608 20085 5648
rect 20043 5599 20085 5608
rect 20427 5648 20469 5657
rect 20427 5608 20428 5648
rect 20468 5608 20469 5648
rect 20427 5599 20469 5608
rect 20811 5648 20853 5657
rect 20811 5608 20812 5648
rect 20852 5608 20853 5648
rect 20811 5599 20853 5608
rect 21195 5648 21237 5657
rect 21195 5608 21196 5648
rect 21236 5608 21237 5648
rect 21195 5599 21237 5608
rect 21579 5648 21621 5657
rect 21579 5608 21580 5648
rect 21620 5608 21621 5648
rect 21579 5599 21621 5608
rect 27339 5648 27381 5657
rect 27339 5608 27340 5648
rect 27380 5608 27381 5648
rect 27339 5599 27381 5608
rect 29451 5648 29493 5657
rect 29451 5608 29452 5648
rect 29492 5608 29493 5648
rect 29451 5599 29493 5608
rect 29835 5648 29877 5657
rect 29835 5608 29836 5648
rect 29876 5608 29877 5648
rect 29835 5599 29877 5608
rect 30075 5648 30117 5657
rect 30075 5608 30076 5648
rect 30116 5608 30117 5648
rect 30075 5599 30117 5608
rect 30250 5648 30308 5649
rect 30250 5608 30259 5648
rect 30299 5608 30308 5648
rect 30250 5607 30308 5608
rect 30603 5648 30645 5657
rect 30603 5608 30604 5648
rect 30644 5608 30645 5648
rect 30603 5599 30645 5608
rect 32043 5648 32085 5657
rect 32043 5608 32044 5648
rect 32084 5608 32085 5648
rect 32043 5599 32085 5608
rect 32427 5648 32469 5657
rect 32427 5608 32428 5648
rect 32468 5608 32469 5648
rect 32427 5599 32469 5608
rect 33003 5648 33045 5657
rect 33003 5608 33004 5648
rect 33044 5608 33045 5648
rect 33003 5599 33045 5608
rect 33243 5648 33285 5657
rect 33243 5608 33244 5648
rect 33284 5608 33285 5648
rect 33243 5599 33285 5608
rect 33963 5648 34005 5657
rect 33963 5608 33964 5648
rect 34004 5608 34005 5648
rect 33963 5599 34005 5608
rect 34203 5648 34245 5657
rect 34203 5608 34204 5648
rect 34244 5608 34245 5648
rect 34203 5599 34245 5608
rect 34635 5648 34677 5657
rect 34635 5608 34636 5648
rect 34676 5608 34677 5648
rect 34635 5599 34677 5608
rect 34875 5648 34917 5657
rect 34875 5608 34876 5648
rect 34916 5608 34917 5648
rect 34875 5599 34917 5608
rect 44523 5648 44565 5657
rect 44523 5608 44524 5648
rect 44564 5608 44565 5648
rect 44523 5599 44565 5608
rect 44907 5648 44949 5657
rect 44907 5608 44908 5648
rect 44948 5608 44949 5648
rect 44907 5599 44949 5608
rect 45147 5648 45189 5657
rect 45147 5608 45148 5648
rect 45188 5608 45189 5648
rect 45147 5599 45189 5608
rect 9723 5564 9765 5573
rect 9723 5524 9724 5564
rect 9764 5524 9765 5564
rect 9723 5515 9765 5524
rect 10107 5564 10149 5573
rect 10107 5524 10108 5564
rect 10148 5524 10149 5564
rect 10107 5515 10149 5524
rect 10491 5564 10533 5573
rect 10491 5524 10492 5564
rect 10532 5524 10533 5564
rect 10491 5515 10533 5524
rect 11259 5564 11301 5573
rect 11259 5524 11260 5564
rect 11300 5524 11301 5564
rect 11259 5515 11301 5524
rect 12027 5564 12069 5573
rect 12027 5524 12028 5564
rect 12068 5524 12069 5564
rect 12027 5515 12069 5524
rect 13467 5564 13509 5573
rect 13467 5524 13468 5564
rect 13508 5524 13509 5564
rect 13467 5515 13509 5524
rect 14331 5564 14373 5573
rect 14331 5524 14332 5564
rect 14372 5524 14373 5564
rect 14331 5515 14373 5524
rect 20187 5564 20229 5573
rect 20187 5524 20188 5564
rect 20228 5524 20229 5564
rect 20187 5515 20229 5524
rect 32283 5564 32325 5573
rect 32283 5524 32284 5564
rect 32324 5524 32325 5564
rect 32283 5515 32325 5524
rect 9339 5480 9381 5489
rect 9339 5440 9340 5480
rect 9380 5440 9381 5480
rect 9339 5431 9381 5440
rect 10875 5480 10917 5489
rect 10875 5440 10876 5480
rect 10916 5440 10917 5480
rect 10875 5431 10917 5440
rect 14715 5480 14757 5489
rect 14715 5440 14716 5480
rect 14756 5440 14757 5480
rect 14715 5431 14757 5440
rect 19419 5480 19461 5489
rect 19419 5440 19420 5480
rect 19460 5440 19461 5480
rect 19419 5431 19461 5440
rect 19803 5480 19845 5489
rect 19803 5440 19804 5480
rect 19844 5440 19845 5480
rect 19803 5431 19845 5440
rect 20571 5480 20613 5489
rect 20571 5440 20572 5480
rect 20612 5440 20613 5480
rect 20571 5431 20613 5440
rect 20955 5480 20997 5489
rect 20955 5440 20956 5480
rect 20996 5440 20997 5480
rect 20955 5431 20997 5440
rect 21339 5480 21381 5489
rect 21339 5440 21340 5480
rect 21380 5440 21381 5480
rect 21339 5431 21381 5440
rect 27579 5480 27621 5489
rect 27579 5440 27580 5480
rect 27620 5440 27621 5480
rect 27579 5431 27621 5440
rect 29691 5480 29733 5489
rect 29691 5440 29692 5480
rect 29732 5440 29733 5480
rect 29691 5431 29733 5440
rect 30459 5480 30501 5489
rect 30459 5440 30460 5480
rect 30500 5440 30501 5480
rect 30459 5431 30501 5440
rect 30843 5480 30885 5489
rect 30843 5440 30844 5480
rect 30884 5440 30885 5480
rect 30843 5431 30885 5440
rect 32667 5480 32709 5489
rect 32667 5440 32668 5480
rect 32708 5440 32709 5480
rect 32667 5431 32709 5440
rect 44763 5480 44805 5489
rect 44763 5440 44764 5480
rect 44804 5440 44805 5480
rect 44763 5431 44805 5440
rect 1152 5312 45216 5336
rect 1152 5272 3688 5312
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 4056 5272 18808 5312
rect 18848 5272 18890 5312
rect 18930 5272 18972 5312
rect 19012 5272 19054 5312
rect 19094 5272 19136 5312
rect 19176 5272 33928 5312
rect 33968 5272 34010 5312
rect 34050 5272 34092 5312
rect 34132 5272 34174 5312
rect 34214 5272 34256 5312
rect 34296 5272 45216 5312
rect 1152 5248 45216 5272
rect 10107 5144 10149 5153
rect 10107 5104 10108 5144
rect 10148 5104 10149 5144
rect 10107 5095 10149 5104
rect 13947 5144 13989 5153
rect 13947 5104 13948 5144
rect 13988 5104 13989 5144
rect 13947 5095 13989 5104
rect 20187 5144 20229 5153
rect 20187 5104 20188 5144
rect 20228 5104 20229 5144
rect 20187 5095 20229 5104
rect 32283 5144 32325 5153
rect 32283 5104 32284 5144
rect 32324 5104 32325 5144
rect 32283 5095 32325 5104
rect 19803 5060 19845 5069
rect 19803 5020 19804 5060
rect 19844 5020 19845 5060
rect 19803 5011 19845 5020
rect 8523 4976 8565 4985
rect 8523 4936 8524 4976
rect 8564 4936 8565 4976
rect 8523 4927 8565 4936
rect 9867 4976 9909 4985
rect 9867 4936 9868 4976
rect 9908 4936 9909 4976
rect 9867 4927 9909 4936
rect 14187 4976 14229 4985
rect 14187 4936 14188 4976
rect 14228 4936 14229 4976
rect 14187 4927 14229 4936
rect 19563 4976 19605 4985
rect 19563 4936 19564 4976
rect 19604 4936 19605 4976
rect 19563 4927 19605 4936
rect 20043 4976 20085 4985
rect 20043 4936 20044 4976
rect 20084 4936 20085 4976
rect 20043 4927 20085 4936
rect 20427 4976 20469 4985
rect 20427 4936 20428 4976
rect 20468 4936 20469 4976
rect 20427 4927 20469 4936
rect 26091 4976 26133 4985
rect 26091 4936 26092 4976
rect 26132 4936 26133 4976
rect 26091 4927 26133 4936
rect 31659 4976 31701 4985
rect 31659 4936 31660 4976
rect 31700 4936 31701 4976
rect 31659 4927 31701 4936
rect 32043 4976 32085 4985
rect 32043 4936 32044 4976
rect 32084 4936 32085 4976
rect 32043 4927 32085 4936
rect 44523 4976 44565 4985
rect 44523 4936 44524 4976
rect 44564 4936 44565 4976
rect 44523 4927 44565 4936
rect 44907 4976 44949 4985
rect 44907 4936 44908 4976
rect 44948 4936 44949 4976
rect 44907 4927 44949 4936
rect 45147 4976 45189 4985
rect 45147 4936 45148 4976
rect 45188 4936 45189 4976
rect 45147 4927 45189 4936
rect 19323 4808 19365 4817
rect 19323 4768 19324 4808
rect 19364 4768 19365 4808
rect 19323 4759 19365 4768
rect 26331 4808 26373 4817
rect 26331 4768 26332 4808
rect 26372 4768 26373 4808
rect 26331 4759 26373 4768
rect 8763 4724 8805 4733
rect 8763 4684 8764 4724
rect 8804 4684 8805 4724
rect 8763 4675 8805 4684
rect 31899 4724 31941 4733
rect 31899 4684 31900 4724
rect 31940 4684 31941 4724
rect 31899 4675 31941 4684
rect 44763 4724 44805 4733
rect 44763 4684 44764 4724
rect 44804 4684 44805 4724
rect 44763 4675 44805 4684
rect 1152 4556 45216 4580
rect 1152 4516 4928 4556
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 5296 4516 20048 4556
rect 20088 4516 20130 4556
rect 20170 4516 20212 4556
rect 20252 4516 20294 4556
rect 20334 4516 20376 4556
rect 20416 4516 35168 4556
rect 35208 4516 35250 4556
rect 35290 4516 35332 4556
rect 35372 4516 35414 4556
rect 35454 4516 35496 4556
rect 35536 4516 45216 4556
rect 1152 4492 45216 4516
rect 24027 4304 24069 4313
rect 24027 4264 24028 4304
rect 24068 4264 24069 4304
rect 24027 4255 24069 4264
rect 26043 4304 26085 4313
rect 26043 4264 26044 4304
rect 26084 4264 26085 4304
rect 26043 4255 26085 4264
rect 34683 4304 34725 4313
rect 34683 4264 34684 4304
rect 34724 4264 34725 4304
rect 34683 4255 34725 4264
rect 45147 4304 45189 4313
rect 45147 4264 45148 4304
rect 45188 4264 45189 4304
rect 45147 4255 45189 4264
rect 23787 4136 23829 4145
rect 23787 4096 23788 4136
rect 23828 4096 23829 4136
rect 23787 4087 23829 4096
rect 25803 4136 25845 4145
rect 25803 4096 25804 4136
rect 25844 4096 25845 4136
rect 25803 4087 25845 4096
rect 34443 4136 34485 4145
rect 34443 4096 34444 4136
rect 34484 4096 34485 4136
rect 34443 4087 34485 4096
rect 44523 4136 44565 4145
rect 44523 4096 44524 4136
rect 44564 4096 44565 4136
rect 44523 4087 44565 4096
rect 44907 4136 44949 4145
rect 44907 4096 44908 4136
rect 44948 4096 44949 4136
rect 44907 4087 44949 4096
rect 44763 4052 44805 4061
rect 44763 4012 44764 4052
rect 44804 4012 44805 4052
rect 44763 4003 44805 4012
rect 1152 3800 45216 3824
rect 1152 3760 3688 3800
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 4056 3760 18808 3800
rect 18848 3760 18890 3800
rect 18930 3760 18972 3800
rect 19012 3760 19054 3800
rect 19094 3760 19136 3800
rect 19176 3760 33928 3800
rect 33968 3760 34010 3800
rect 34050 3760 34092 3800
rect 34132 3760 34174 3800
rect 34214 3760 34256 3800
rect 34296 3760 45216 3800
rect 1152 3736 45216 3760
rect 27003 3632 27045 3641
rect 27003 3592 27004 3632
rect 27044 3592 27045 3632
rect 27003 3583 27045 3592
rect 32091 3632 32133 3641
rect 32091 3592 32092 3632
rect 32132 3592 32133 3632
rect 32091 3583 32133 3592
rect 45147 3632 45189 3641
rect 45147 3592 45148 3632
rect 45188 3592 45189 3632
rect 45147 3583 45189 3592
rect 26139 3548 26181 3557
rect 26139 3508 26140 3548
rect 26180 3508 26181 3548
rect 26139 3499 26181 3508
rect 18987 3464 19029 3473
rect 18987 3424 18988 3464
rect 19028 3424 19029 3464
rect 18987 3415 19029 3424
rect 19755 3464 19797 3473
rect 19755 3424 19756 3464
rect 19796 3424 19797 3464
rect 19755 3415 19797 3424
rect 21003 3464 21045 3473
rect 21003 3424 21004 3464
rect 21044 3424 21045 3464
rect 21003 3415 21045 3424
rect 21387 3464 21429 3473
rect 21387 3424 21388 3464
rect 21428 3424 21429 3464
rect 21387 3415 21429 3424
rect 21771 3464 21813 3473
rect 21771 3424 21772 3464
rect 21812 3424 21813 3464
rect 21771 3415 21813 3424
rect 22635 3464 22677 3473
rect 22635 3424 22636 3464
rect 22676 3424 22677 3464
rect 22635 3415 22677 3424
rect 23019 3464 23061 3473
rect 23019 3424 23020 3464
rect 23060 3424 23061 3464
rect 23019 3415 23061 3424
rect 23403 3464 23445 3473
rect 23403 3424 23404 3464
rect 23444 3424 23445 3464
rect 23403 3415 23445 3424
rect 24075 3464 24117 3473
rect 24075 3424 24076 3464
rect 24116 3424 24117 3464
rect 24075 3415 24117 3424
rect 24459 3464 24501 3473
rect 24459 3424 24460 3464
rect 24500 3424 24501 3464
rect 24459 3415 24501 3424
rect 24843 3464 24885 3473
rect 24843 3424 24844 3464
rect 24884 3424 24885 3464
rect 24843 3415 24885 3424
rect 25899 3464 25941 3473
rect 25899 3424 25900 3464
rect 25940 3424 25941 3464
rect 25899 3415 25941 3424
rect 26763 3464 26805 3473
rect 26763 3424 26764 3464
rect 26804 3424 26805 3464
rect 26763 3415 26805 3424
rect 27627 3464 27669 3473
rect 27627 3424 27628 3464
rect 27668 3424 27669 3464
rect 27627 3415 27669 3424
rect 27867 3464 27909 3473
rect 27867 3424 27868 3464
rect 27908 3424 27909 3464
rect 27867 3415 27909 3424
rect 31851 3464 31893 3473
rect 31851 3424 31852 3464
rect 31892 3424 31893 3464
rect 31851 3415 31893 3424
rect 44523 3464 44565 3473
rect 44523 3424 44524 3464
rect 44564 3424 44565 3464
rect 44523 3415 44565 3424
rect 44907 3464 44949 3473
rect 44907 3424 44908 3464
rect 44948 3424 44949 3464
rect 44907 3415 44949 3424
rect 25083 3296 25125 3305
rect 25083 3256 25084 3296
rect 25124 3256 25125 3296
rect 25083 3247 25125 3256
rect 44763 3296 44805 3305
rect 44763 3256 44764 3296
rect 44804 3256 44805 3296
rect 44763 3247 44805 3256
rect 19227 3212 19269 3221
rect 19227 3172 19228 3212
rect 19268 3172 19269 3212
rect 19227 3163 19269 3172
rect 19995 3212 20037 3221
rect 19995 3172 19996 3212
rect 20036 3172 20037 3212
rect 19995 3163 20037 3172
rect 21243 3212 21285 3221
rect 21243 3172 21244 3212
rect 21284 3172 21285 3212
rect 21243 3163 21285 3172
rect 21627 3212 21669 3221
rect 21627 3172 21628 3212
rect 21668 3172 21669 3212
rect 21627 3163 21669 3172
rect 22011 3212 22053 3221
rect 22011 3172 22012 3212
rect 22052 3172 22053 3212
rect 22011 3163 22053 3172
rect 22875 3212 22917 3221
rect 22875 3172 22876 3212
rect 22916 3172 22917 3212
rect 22875 3163 22917 3172
rect 23259 3212 23301 3221
rect 23259 3172 23260 3212
rect 23300 3172 23301 3212
rect 23259 3163 23301 3172
rect 23643 3212 23685 3221
rect 23643 3172 23644 3212
rect 23684 3172 23685 3212
rect 23643 3163 23685 3172
rect 24315 3212 24357 3221
rect 24315 3172 24316 3212
rect 24356 3172 24357 3212
rect 24315 3163 24357 3172
rect 24699 3212 24741 3221
rect 24699 3172 24700 3212
rect 24740 3172 24741 3212
rect 24699 3163 24741 3172
rect 34443 3212 34485 3221
rect 34443 3172 34444 3212
rect 34484 3172 34485 3212
rect 34443 3163 34485 3172
rect 34714 3212 34772 3213
rect 34714 3172 34723 3212
rect 34763 3172 34772 3212
rect 34714 3171 34772 3172
rect 1152 3044 45216 3068
rect 1152 3004 4928 3044
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 5296 3004 20048 3044
rect 20088 3004 20130 3044
rect 20170 3004 20212 3044
rect 20252 3004 20294 3044
rect 20334 3004 20376 3044
rect 20416 3004 35168 3044
rect 35208 3004 35250 3044
rect 35290 3004 35332 3044
rect 35372 3004 35414 3044
rect 35454 3004 35496 3044
rect 35536 3004 45216 3044
rect 1152 2980 45216 3004
rect 18267 2876 18309 2885
rect 18267 2836 18268 2876
rect 18308 2836 18309 2876
rect 18267 2827 18309 2836
rect 45147 2876 45189 2885
rect 45147 2836 45148 2876
rect 45188 2836 45189 2876
rect 45147 2827 45189 2836
rect 11307 2624 11349 2633
rect 11307 2584 11308 2624
rect 11348 2584 11349 2624
rect 11307 2575 11349 2584
rect 18027 2624 18069 2633
rect 18027 2584 18028 2624
rect 18068 2584 18069 2624
rect 18027 2575 18069 2584
rect 27147 2624 27189 2633
rect 27147 2584 27148 2624
rect 27188 2584 27189 2624
rect 27147 2575 27189 2584
rect 28011 2624 28053 2633
rect 28011 2584 28012 2624
rect 28052 2584 28053 2624
rect 28011 2575 28053 2584
rect 44139 2624 44181 2633
rect 44139 2584 44140 2624
rect 44180 2584 44181 2624
rect 44139 2575 44181 2584
rect 44523 2624 44565 2633
rect 44523 2584 44524 2624
rect 44564 2584 44565 2624
rect 44523 2575 44565 2584
rect 44907 2624 44949 2633
rect 44907 2584 44908 2624
rect 44948 2584 44949 2624
rect 44907 2575 44949 2584
rect 27387 2540 27429 2549
rect 27387 2500 27388 2540
rect 27428 2500 27429 2540
rect 27387 2491 27429 2500
rect 44763 2540 44805 2549
rect 44763 2500 44764 2540
rect 44804 2500 44805 2540
rect 44763 2491 44805 2500
rect 11547 2456 11589 2465
rect 11547 2416 11548 2456
rect 11588 2416 11589 2456
rect 11547 2407 11589 2416
rect 28251 2456 28293 2465
rect 28251 2416 28252 2456
rect 28292 2416 28293 2456
rect 28251 2407 28293 2416
rect 44379 2456 44421 2465
rect 44379 2416 44380 2456
rect 44420 2416 44421 2456
rect 44379 2407 44421 2416
rect 1152 2288 45216 2312
rect 1152 2248 3688 2288
rect 3728 2248 3770 2288
rect 3810 2248 3852 2288
rect 3892 2248 3934 2288
rect 3974 2248 4016 2288
rect 4056 2248 18808 2288
rect 18848 2248 18890 2288
rect 18930 2248 18972 2288
rect 19012 2248 19054 2288
rect 19094 2248 19136 2288
rect 19176 2248 33928 2288
rect 33968 2248 34010 2288
rect 34050 2248 34092 2288
rect 34132 2248 34174 2288
rect 34214 2248 34256 2288
rect 34296 2248 45216 2288
rect 1152 2224 45216 2248
rect 45147 2120 45189 2129
rect 45147 2080 45148 2120
rect 45188 2080 45189 2120
rect 45147 2071 45189 2080
rect 43371 1952 43413 1961
rect 43371 1912 43372 1952
rect 43412 1912 43413 1952
rect 43371 1903 43413 1912
rect 43755 1952 43797 1961
rect 43755 1912 43756 1952
rect 43796 1912 43797 1952
rect 43755 1903 43797 1912
rect 44139 1952 44181 1961
rect 44139 1912 44140 1952
rect 44180 1912 44181 1952
rect 44139 1903 44181 1912
rect 44523 1952 44565 1961
rect 44523 1912 44524 1952
rect 44564 1912 44565 1952
rect 44523 1903 44565 1912
rect 44907 1952 44949 1961
rect 44907 1912 44908 1952
rect 44948 1912 44949 1952
rect 44907 1903 44949 1912
rect 43995 1784 44037 1793
rect 43995 1744 43996 1784
rect 44036 1744 44037 1784
rect 43995 1735 44037 1744
rect 43611 1700 43653 1709
rect 43611 1660 43612 1700
rect 43652 1660 43653 1700
rect 43611 1651 43653 1660
rect 44379 1700 44421 1709
rect 44379 1660 44380 1700
rect 44420 1660 44421 1700
rect 44379 1651 44421 1660
rect 44763 1700 44805 1709
rect 44763 1660 44764 1700
rect 44804 1660 44805 1700
rect 44763 1651 44805 1660
rect 1152 1532 45216 1556
rect 1152 1492 4928 1532
rect 4968 1492 5010 1532
rect 5050 1492 5092 1532
rect 5132 1492 5174 1532
rect 5214 1492 5256 1532
rect 5296 1492 20048 1532
rect 20088 1492 20130 1532
rect 20170 1492 20212 1532
rect 20252 1492 20294 1532
rect 20334 1492 20376 1532
rect 20416 1492 35168 1532
rect 35208 1492 35250 1532
rect 35290 1492 35332 1532
rect 35372 1492 35414 1532
rect 35454 1492 35496 1532
rect 35536 1492 45216 1532
rect 1152 1468 45216 1492
<< via1 >>
rect 3688 9808 3728 9848
rect 3770 9808 3810 9848
rect 3852 9808 3892 9848
rect 3934 9808 3974 9848
rect 4016 9808 4056 9848
rect 18808 9808 18848 9848
rect 18890 9808 18930 9848
rect 18972 9808 19012 9848
rect 19054 9808 19094 9848
rect 19136 9808 19176 9848
rect 33928 9808 33968 9848
rect 34010 9808 34050 9848
rect 34092 9808 34132 9848
rect 34174 9808 34214 9848
rect 34256 9808 34296 9848
rect 10972 9640 11012 9680
rect 11356 9640 11396 9680
rect 11740 9640 11780 9680
rect 12124 9640 12164 9680
rect 12508 9640 12548 9680
rect 12892 9640 12932 9680
rect 13276 9640 13316 9680
rect 13660 9640 13700 9680
rect 14044 9640 14084 9680
rect 14428 9640 14468 9680
rect 14812 9640 14852 9680
rect 15196 9640 15236 9680
rect 15580 9640 15620 9680
rect 15964 9640 16004 9680
rect 16348 9640 16388 9680
rect 16732 9640 16772 9680
rect 17116 9640 17156 9680
rect 17500 9640 17540 9680
rect 17884 9640 17924 9680
rect 18268 9640 18308 9680
rect 18652 9640 18692 9680
rect 19036 9640 19076 9680
rect 20188 9640 20228 9680
rect 20668 9640 20708 9680
rect 21436 9640 21476 9680
rect 31228 9640 31268 9680
rect 31996 9640 32036 9680
rect 32764 9640 32804 9680
rect 33148 9640 33188 9680
rect 34684 9640 34724 9680
rect 36220 9640 36260 9680
rect 43228 9640 43268 9680
rect 43612 9640 43652 9680
rect 43996 9640 44036 9680
rect 19420 9556 19460 9596
rect 20284 9556 20324 9596
rect 31612 9556 31652 9596
rect 32380 9556 32420 9596
rect 36604 9556 36644 9596
rect 10732 9472 10772 9512
rect 11116 9472 11156 9512
rect 11500 9472 11540 9512
rect 11884 9472 11924 9512
rect 12268 9472 12308 9512
rect 12652 9472 12692 9512
rect 13036 9472 13076 9512
rect 13420 9472 13460 9512
rect 13804 9472 13844 9512
rect 14188 9472 14228 9512
rect 14572 9472 14612 9512
rect 14956 9472 14996 9512
rect 15340 9472 15380 9512
rect 15724 9472 15764 9512
rect 16108 9472 16148 9512
rect 16492 9472 16532 9512
rect 16876 9472 16916 9512
rect 17260 9472 17300 9512
rect 17644 9472 17684 9512
rect 18028 9472 18068 9512
rect 18412 9472 18452 9512
rect 18796 9472 18836 9512
rect 19180 9472 19220 9512
rect 19564 9472 19604 9512
rect 19948 9472 19988 9512
rect 20524 9472 20564 9512
rect 20908 9472 20948 9512
rect 21676 9472 21716 9512
rect 31468 9472 31508 9512
rect 31852 9472 31892 9512
rect 32236 9472 32276 9512
rect 32620 9472 32660 9512
rect 33004 9472 33044 9512
rect 33388 9472 33428 9512
rect 33532 9472 33572 9512
rect 33772 9472 33812 9512
rect 34156 9472 34196 9512
rect 34540 9472 34580 9512
rect 34924 9472 34964 9512
rect 35308 9472 35348 9512
rect 35692 9472 35732 9512
rect 36076 9472 36116 9512
rect 36460 9472 36500 9512
rect 36844 9472 36884 9512
rect 37132 9472 37172 9512
rect 37708 9472 37748 9512
rect 37900 9472 37940 9512
rect 38476 9472 38516 9512
rect 39052 9472 39092 9512
rect 39628 9472 39668 9512
rect 39916 9472 39956 9512
rect 40492 9472 40532 9512
rect 40780 9472 40820 9512
rect 42988 9472 43028 9512
rect 43372 9472 43412 9512
rect 43756 9472 43796 9512
rect 44140 9472 44180 9512
rect 44524 9472 44564 9512
rect 44908 9472 44948 9512
rect 19804 9304 19844 9344
rect 34300 9304 34340 9344
rect 35836 9304 35876 9344
rect 44380 9304 44420 9344
rect 21100 9220 21140 9260
rect 33916 9220 33956 9260
rect 35068 9220 35108 9260
rect 35452 9220 35492 9260
rect 37036 9220 37076 9260
rect 37315 9220 37355 9260
rect 37891 9220 37931 9260
rect 38188 9220 38228 9260
rect 38764 9220 38804 9260
rect 39331 9220 39371 9260
rect 40204 9220 40244 9260
rect 44764 9220 44804 9260
rect 45148 9220 45188 9260
rect 4928 9052 4968 9092
rect 5010 9052 5050 9092
rect 5092 9052 5132 9092
rect 5174 9052 5214 9092
rect 5256 9052 5296 9092
rect 20048 9052 20088 9092
rect 20130 9052 20170 9092
rect 20212 9052 20252 9092
rect 20294 9052 20334 9092
rect 20376 9052 20416 9092
rect 35168 9052 35208 9092
rect 35250 9052 35290 9092
rect 35332 9052 35372 9092
rect 35414 9052 35454 9092
rect 35496 9052 35536 9092
rect 11068 8884 11108 8924
rect 11452 8884 11492 8924
rect 11836 8884 11876 8924
rect 12220 8884 12260 8924
rect 12604 8884 12644 8924
rect 13372 8884 13412 8924
rect 13756 8884 13796 8924
rect 14140 8884 14180 8924
rect 14524 8884 14564 8924
rect 14908 8884 14948 8924
rect 15292 8884 15332 8924
rect 15676 8884 15716 8924
rect 16060 8884 16100 8924
rect 16444 8884 16484 8924
rect 16828 8884 16868 8924
rect 17212 8884 17252 8924
rect 17596 8884 17636 8924
rect 17980 8884 18020 8924
rect 18364 8884 18404 8924
rect 18748 8884 18788 8924
rect 19132 8884 19172 8924
rect 19516 8884 19556 8924
rect 19900 8884 19940 8924
rect 27196 8884 27236 8924
rect 27580 8884 27620 8924
rect 32188 8884 32228 8924
rect 32572 8884 32612 8924
rect 32956 8884 32996 8924
rect 33340 8884 33380 8924
rect 34243 8884 34283 8924
rect 34876 8884 34916 8924
rect 37219 8884 37259 8924
rect 37756 8884 37796 8924
rect 40003 8884 40043 8924
rect 43996 8884 44036 8924
rect 44380 8884 44420 8924
rect 25852 8800 25892 8840
rect 26428 8800 26468 8840
rect 27964 8800 28004 8840
rect 32092 8800 32132 8840
rect 35260 8800 35300 8840
rect 36316 8800 36356 8840
rect 36700 8800 36740 8840
rect 38140 8800 38180 8840
rect 11251 8632 11291 8672
rect 11692 8632 11732 8672
rect 12076 8632 12116 8672
rect 12460 8632 12500 8672
rect 12844 8632 12884 8672
rect 13228 8632 13268 8672
rect 13612 8632 13652 8672
rect 13996 8632 14036 8672
rect 14380 8632 14420 8672
rect 14764 8632 14804 8672
rect 15148 8632 15188 8672
rect 15532 8632 15572 8672
rect 15916 8632 15956 8672
rect 16300 8632 16340 8672
rect 16684 8632 16724 8672
rect 17068 8632 17108 8672
rect 17452 8632 17492 8672
rect 17836 8632 17876 8672
rect 18220 8632 18260 8672
rect 18604 8632 18644 8672
rect 18988 8632 19028 8672
rect 19372 8632 19412 8672
rect 19756 8632 19796 8672
rect 20140 8632 20180 8672
rect 26092 8632 26132 8672
rect 26668 8632 26708 8672
rect 27436 8632 27476 8672
rect 27820 8632 27860 8672
rect 28204 8632 28244 8672
rect 28348 8632 28388 8672
rect 28588 8632 28628 8672
rect 28732 8632 28772 8672
rect 28972 8632 29012 8672
rect 31852 8632 31892 8672
rect 32428 8632 32468 8672
rect 32812 8632 32852 8672
rect 33196 8632 33236 8672
rect 33580 8632 33620 8672
rect 33868 8632 33908 8672
rect 34252 8632 34292 8672
rect 34540 8632 34580 8672
rect 35116 8632 35156 8672
rect 35500 8632 35540 8672
rect 35788 8632 35828 8672
rect 36076 8632 36116 8672
rect 36460 8632 36500 8672
rect 36844 8632 36884 8672
rect 37228 8632 37268 8672
rect 37516 8632 37556 8672
rect 37900 8632 37940 8672
rect 38284 8632 38324 8672
rect 38572 8632 38612 8672
rect 38860 8632 38900 8672
rect 39148 8632 39188 8672
rect 39436 8632 39476 8672
rect 39724 8632 39764 8672
rect 40300 8632 40340 8672
rect 43756 8632 43796 8672
rect 44140 8632 44180 8672
rect 44524 8632 44564 8672
rect 44908 8632 44948 8672
rect 12988 8548 13028 8588
rect 34780 8548 34820 8588
rect 34108 8464 34148 8504
rect 44764 8464 44804 8504
rect 45148 8464 45188 8504
rect 3688 8296 3728 8336
rect 3770 8296 3810 8336
rect 3852 8296 3892 8336
rect 3934 8296 3974 8336
rect 4016 8296 4056 8336
rect 18808 8296 18848 8336
rect 18890 8296 18930 8336
rect 18972 8296 19012 8336
rect 19054 8296 19094 8336
rect 19136 8296 19176 8336
rect 33928 8296 33968 8336
rect 34010 8296 34050 8336
rect 34092 8296 34132 8336
rect 34174 8296 34214 8336
rect 34256 8296 34296 8336
rect 25564 8128 25604 8168
rect 25948 8128 25988 8168
rect 26716 8128 26756 8168
rect 27100 8128 27140 8168
rect 32956 8128 32996 8168
rect 39772 8128 39812 8168
rect 43132 8128 43172 8168
rect 26332 8044 26372 8084
rect 25180 7960 25220 8000
rect 25420 7960 25460 8000
rect 25804 7960 25844 8000
rect 26188 7960 26228 8000
rect 26572 7960 26612 8000
rect 26956 7960 26996 8000
rect 27340 7960 27380 8000
rect 27484 7960 27524 8000
rect 27724 7960 27764 8000
rect 28204 7960 28244 8000
rect 32716 7960 32756 8000
rect 34348 7960 34388 8000
rect 34636 7960 34676 8000
rect 34924 7960 34964 8000
rect 35212 7960 35252 8000
rect 35500 7960 35540 8000
rect 35788 7960 35828 8000
rect 36076 7960 36116 8000
rect 36460 7960 36500 8000
rect 36700 7960 36740 8000
rect 38380 7960 38420 8000
rect 38668 7960 38708 8000
rect 39532 7960 39572 8000
rect 43372 7960 43412 8000
rect 44524 7960 44564 8000
rect 44908 7960 44948 8000
rect 36940 7876 36980 7916
rect 37132 7876 37172 7916
rect 27964 7708 28004 7748
rect 37411 7708 37451 7748
rect 37699 7708 37739 7748
rect 37987 7708 38027 7748
rect 44764 7708 44804 7748
rect 45148 7708 45188 7748
rect 4928 7540 4968 7580
rect 5010 7540 5050 7580
rect 5092 7540 5132 7580
rect 5174 7540 5214 7580
rect 5256 7540 5296 7580
rect 20048 7540 20088 7580
rect 20130 7540 20170 7580
rect 20212 7540 20252 7580
rect 20294 7540 20334 7580
rect 20376 7540 20416 7580
rect 35168 7540 35208 7580
rect 35250 7540 35290 7580
rect 35332 7540 35372 7580
rect 35414 7540 35454 7580
rect 35496 7540 35536 7580
rect 36076 7372 36116 7412
rect 8332 7120 8372 7160
rect 25900 7120 25940 7160
rect 33292 7120 33332 7160
rect 35692 7120 35732 7160
rect 35932 7120 35972 7160
rect 44524 7120 44564 7160
rect 44908 7120 44948 7160
rect 8572 7036 8612 7076
rect 33532 7036 33572 7076
rect 25660 6952 25700 6992
rect 44764 6952 44804 6992
rect 45148 6952 45188 6992
rect 3688 6784 3728 6824
rect 3770 6784 3810 6824
rect 3852 6784 3892 6824
rect 3934 6784 3974 6824
rect 4016 6784 4056 6824
rect 18808 6784 18848 6824
rect 18890 6784 18930 6824
rect 18972 6784 19012 6824
rect 19054 6784 19094 6824
rect 19136 6784 19176 6824
rect 33928 6784 33968 6824
rect 34010 6784 34050 6824
rect 34092 6784 34132 6824
rect 34174 6784 34214 6824
rect 34256 6784 34296 6824
rect 7612 6616 7652 6656
rect 8668 6532 8708 6572
rect 9052 6532 9092 6572
rect 9436 6532 9476 6572
rect 13948 6532 13988 6572
rect 19132 6532 19172 6572
rect 7372 6448 7412 6488
rect 7756 6448 7796 6488
rect 8428 6448 8468 6488
rect 8812 6448 8852 6488
rect 9196 6448 9236 6488
rect 13708 6448 13748 6488
rect 19372 6448 19412 6488
rect 19804 6448 19844 6488
rect 20044 6448 20084 6488
rect 20428 6448 20468 6488
rect 33772 6448 33812 6488
rect 35788 6448 35828 6488
rect 35980 6448 36020 6488
rect 44524 6448 44564 6488
rect 44908 6448 44948 6488
rect 7996 6280 8036 6320
rect 45148 6280 45188 6320
rect 20188 6196 20228 6236
rect 34012 6196 34052 6236
rect 44764 6196 44804 6236
rect 4928 6028 4968 6068
rect 5010 6028 5050 6068
rect 5092 6028 5132 6068
rect 5174 6028 5214 6068
rect 5256 6028 5296 6068
rect 20048 6028 20088 6068
rect 20130 6028 20170 6068
rect 20212 6028 20252 6068
rect 20294 6028 20334 6068
rect 20376 6028 20416 6068
rect 35168 6028 35208 6068
rect 35250 6028 35290 6068
rect 35332 6028 35372 6068
rect 35414 6028 35454 6068
rect 35496 6028 35536 6068
rect 18268 5776 18308 5816
rect 18652 5776 18692 5816
rect 19036 5776 19076 5816
rect 9100 5608 9140 5648
rect 9484 5608 9524 5648
rect 9868 5608 9908 5648
rect 10252 5608 10292 5648
rect 10636 5608 10676 5648
rect 11020 5608 11060 5648
rect 11356 5608 11396 5648
rect 11596 5608 11636 5648
rect 11827 5608 11867 5648
rect 13228 5608 13268 5648
rect 13564 5608 13604 5648
rect 13804 5608 13844 5648
rect 13996 5608 14036 5648
rect 14236 5608 14276 5648
rect 14572 5608 14612 5648
rect 14956 5608 14996 5648
rect 15100 5608 15140 5648
rect 15340 5608 15380 5648
rect 17884 5608 17924 5648
rect 18124 5608 18164 5648
rect 18508 5608 18548 5648
rect 18892 5608 18932 5648
rect 19276 5608 19316 5648
rect 19660 5608 19700 5648
rect 20044 5608 20084 5648
rect 20428 5608 20468 5648
rect 20812 5608 20852 5648
rect 21196 5608 21236 5648
rect 21580 5608 21620 5648
rect 27340 5608 27380 5648
rect 29452 5608 29492 5648
rect 29836 5608 29876 5648
rect 30076 5608 30116 5648
rect 30259 5608 30299 5648
rect 30604 5608 30644 5648
rect 32044 5608 32084 5648
rect 32428 5608 32468 5648
rect 33004 5608 33044 5648
rect 33244 5608 33284 5648
rect 33964 5608 34004 5648
rect 34204 5608 34244 5648
rect 34636 5608 34676 5648
rect 34876 5608 34916 5648
rect 44524 5608 44564 5648
rect 44908 5608 44948 5648
rect 45148 5608 45188 5648
rect 9724 5524 9764 5564
rect 10108 5524 10148 5564
rect 10492 5524 10532 5564
rect 11260 5524 11300 5564
rect 12028 5524 12068 5564
rect 13468 5524 13508 5564
rect 14332 5524 14372 5564
rect 20188 5524 20228 5564
rect 32284 5524 32324 5564
rect 9340 5440 9380 5480
rect 10876 5440 10916 5480
rect 14716 5440 14756 5480
rect 19420 5440 19460 5480
rect 19804 5440 19844 5480
rect 20572 5440 20612 5480
rect 20956 5440 20996 5480
rect 21340 5440 21380 5480
rect 27580 5440 27620 5480
rect 29692 5440 29732 5480
rect 30460 5440 30500 5480
rect 30844 5440 30884 5480
rect 32668 5440 32708 5480
rect 44764 5440 44804 5480
rect 3688 5272 3728 5312
rect 3770 5272 3810 5312
rect 3852 5272 3892 5312
rect 3934 5272 3974 5312
rect 4016 5272 4056 5312
rect 18808 5272 18848 5312
rect 18890 5272 18930 5312
rect 18972 5272 19012 5312
rect 19054 5272 19094 5312
rect 19136 5272 19176 5312
rect 33928 5272 33968 5312
rect 34010 5272 34050 5312
rect 34092 5272 34132 5312
rect 34174 5272 34214 5312
rect 34256 5272 34296 5312
rect 10108 5104 10148 5144
rect 13948 5104 13988 5144
rect 20188 5104 20228 5144
rect 32284 5104 32324 5144
rect 19804 5020 19844 5060
rect 8524 4936 8564 4976
rect 9868 4936 9908 4976
rect 14188 4936 14228 4976
rect 19564 4936 19604 4976
rect 20044 4936 20084 4976
rect 20428 4936 20468 4976
rect 26092 4936 26132 4976
rect 31660 4936 31700 4976
rect 32044 4936 32084 4976
rect 44524 4936 44564 4976
rect 44908 4936 44948 4976
rect 45148 4936 45188 4976
rect 19324 4768 19364 4808
rect 26332 4768 26372 4808
rect 8764 4684 8804 4724
rect 31900 4684 31940 4724
rect 44764 4684 44804 4724
rect 4928 4516 4968 4556
rect 5010 4516 5050 4556
rect 5092 4516 5132 4556
rect 5174 4516 5214 4556
rect 5256 4516 5296 4556
rect 20048 4516 20088 4556
rect 20130 4516 20170 4556
rect 20212 4516 20252 4556
rect 20294 4516 20334 4556
rect 20376 4516 20416 4556
rect 35168 4516 35208 4556
rect 35250 4516 35290 4556
rect 35332 4516 35372 4556
rect 35414 4516 35454 4556
rect 35496 4516 35536 4556
rect 24028 4264 24068 4304
rect 26044 4264 26084 4304
rect 34684 4264 34724 4304
rect 45148 4264 45188 4304
rect 23788 4096 23828 4136
rect 25804 4096 25844 4136
rect 34444 4096 34484 4136
rect 44524 4096 44564 4136
rect 44908 4096 44948 4136
rect 44764 4012 44804 4052
rect 3688 3760 3728 3800
rect 3770 3760 3810 3800
rect 3852 3760 3892 3800
rect 3934 3760 3974 3800
rect 4016 3760 4056 3800
rect 18808 3760 18848 3800
rect 18890 3760 18930 3800
rect 18972 3760 19012 3800
rect 19054 3760 19094 3800
rect 19136 3760 19176 3800
rect 33928 3760 33968 3800
rect 34010 3760 34050 3800
rect 34092 3760 34132 3800
rect 34174 3760 34214 3800
rect 34256 3760 34296 3800
rect 27004 3592 27044 3632
rect 32092 3592 32132 3632
rect 45148 3592 45188 3632
rect 26140 3508 26180 3548
rect 18988 3424 19028 3464
rect 19756 3424 19796 3464
rect 21004 3424 21044 3464
rect 21388 3424 21428 3464
rect 21772 3424 21812 3464
rect 22636 3424 22676 3464
rect 23020 3424 23060 3464
rect 23404 3424 23444 3464
rect 24076 3424 24116 3464
rect 24460 3424 24500 3464
rect 24844 3424 24884 3464
rect 25900 3424 25940 3464
rect 26764 3424 26804 3464
rect 27628 3424 27668 3464
rect 27868 3424 27908 3464
rect 31852 3424 31892 3464
rect 44524 3424 44564 3464
rect 44908 3424 44948 3464
rect 25084 3256 25124 3296
rect 44764 3256 44804 3296
rect 19228 3172 19268 3212
rect 19996 3172 20036 3212
rect 21244 3172 21284 3212
rect 21628 3172 21668 3212
rect 22012 3172 22052 3212
rect 22876 3172 22916 3212
rect 23260 3172 23300 3212
rect 23644 3172 23684 3212
rect 24316 3172 24356 3212
rect 24700 3172 24740 3212
rect 34444 3172 34484 3212
rect 34723 3172 34763 3212
rect 4928 3004 4968 3044
rect 5010 3004 5050 3044
rect 5092 3004 5132 3044
rect 5174 3004 5214 3044
rect 5256 3004 5296 3044
rect 20048 3004 20088 3044
rect 20130 3004 20170 3044
rect 20212 3004 20252 3044
rect 20294 3004 20334 3044
rect 20376 3004 20416 3044
rect 35168 3004 35208 3044
rect 35250 3004 35290 3044
rect 35332 3004 35372 3044
rect 35414 3004 35454 3044
rect 35496 3004 35536 3044
rect 18268 2836 18308 2876
rect 45148 2836 45188 2876
rect 11308 2584 11348 2624
rect 18028 2584 18068 2624
rect 27148 2584 27188 2624
rect 28012 2584 28052 2624
rect 44140 2584 44180 2624
rect 44524 2584 44564 2624
rect 44908 2584 44948 2624
rect 27388 2500 27428 2540
rect 44764 2500 44804 2540
rect 11548 2416 11588 2456
rect 28252 2416 28292 2456
rect 44380 2416 44420 2456
rect 3688 2248 3728 2288
rect 3770 2248 3810 2288
rect 3852 2248 3892 2288
rect 3934 2248 3974 2288
rect 4016 2248 4056 2288
rect 18808 2248 18848 2288
rect 18890 2248 18930 2288
rect 18972 2248 19012 2288
rect 19054 2248 19094 2288
rect 19136 2248 19176 2288
rect 33928 2248 33968 2288
rect 34010 2248 34050 2288
rect 34092 2248 34132 2288
rect 34174 2248 34214 2288
rect 34256 2248 34296 2288
rect 45148 2080 45188 2120
rect 43372 1912 43412 1952
rect 43756 1912 43796 1952
rect 44140 1912 44180 1952
rect 44524 1912 44564 1952
rect 44908 1912 44948 1952
rect 43996 1744 44036 1784
rect 43612 1660 43652 1700
rect 44380 1660 44420 1700
rect 44764 1660 44804 1700
rect 4928 1492 4968 1532
rect 5010 1492 5050 1532
rect 5092 1492 5132 1532
rect 5174 1492 5214 1532
rect 5256 1492 5296 1532
rect 20048 1492 20088 1532
rect 20130 1492 20170 1532
rect 20212 1492 20252 1532
rect 20294 1492 20334 1532
rect 20376 1492 20416 1532
rect 35168 1492 35208 1532
rect 35250 1492 35290 1532
rect 35332 1492 35372 1532
rect 35414 1492 35454 1532
rect 35496 1492 35536 1532
<< metal2 >>
rect 9571 11740 9580 11780
rect 9620 11740 22156 11780
rect 22196 11740 22205 11780
rect 9859 11656 9868 11696
rect 9908 11656 22348 11696
rect 22388 11656 22397 11696
rect 16483 11572 16492 11612
rect 16532 11572 24460 11612
rect 24500 11572 24509 11612
rect 10051 11488 10060 11528
rect 10100 11488 21964 11528
rect 22004 11488 22013 11528
rect 16291 11320 16300 11360
rect 16340 11320 23308 11360
rect 23348 11320 23357 11360
rect 0 11024 90 11044
rect 46278 11024 46368 11044
rect 0 10984 1324 11024
rect 1364 10984 1373 11024
rect 15331 10984 15340 11024
rect 15380 10984 21772 11024
rect 21812 10984 21821 11024
rect 44131 10984 44140 11024
rect 44180 10984 46368 11024
rect 0 10964 90 10984
rect 46278 10964 46368 10984
rect 0 10688 90 10708
rect 46278 10688 46368 10708
rect 0 10648 268 10688
rect 308 10648 317 10688
rect 19939 10648 19948 10688
rect 19988 10648 23884 10688
rect 23924 10648 23933 10688
rect 43363 10648 43372 10688
rect 43412 10648 46368 10688
rect 0 10628 90 10648
rect 46278 10628 46368 10648
rect 0 10352 90 10372
rect 46278 10352 46368 10372
rect 0 10312 556 10352
rect 596 10312 605 10352
rect 43651 10312 43660 10352
rect 43700 10312 46368 10352
rect 0 10292 90 10312
rect 46278 10292 46368 10312
rect 19555 10228 19564 10268
rect 19604 10228 23692 10268
rect 23732 10228 23741 10268
rect 20332 10144 20756 10184
rect 20332 10100 20372 10144
rect 20716 10100 20756 10144
rect 33484 10144 34772 10184
rect 33484 10100 33524 10144
rect 34732 10100 34772 10144
rect 18019 10060 18028 10100
rect 18068 10060 20372 10100
rect 20640 10060 20716 10100
rect 20756 10060 20765 10100
rect 32611 10060 32620 10100
rect 32660 10060 33524 10100
rect 33580 10060 34484 10100
rect 34732 10060 36076 10100
rect 36116 10060 36125 10100
rect 0 10016 90 10036
rect 33580 10016 33620 10060
rect 0 9976 1420 10016
rect 1460 9976 1469 10016
rect 19372 9976 20524 10016
rect 20564 9976 20573 10016
rect 32419 9976 32428 10016
rect 32468 9976 33620 10016
rect 0 9956 90 9976
rect 19372 9932 19412 9976
rect 34444 9932 34484 10060
rect 46278 10016 46368 10036
rect 34819 9976 34828 10016
rect 34868 9976 35828 10016
rect 44419 9976 44428 10016
rect 44468 9976 46368 10016
rect 17635 9892 17644 9932
rect 17684 9892 19412 9932
rect 19468 9892 27052 9932
rect 27092 9892 27101 9932
rect 30499 9892 30508 9932
rect 30548 9892 34388 9932
rect 34444 9892 35692 9932
rect 35732 9892 35741 9932
rect 3679 9808 3688 9848
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 4056 9808 4065 9848
rect 18799 9808 18808 9848
rect 18848 9808 18890 9848
rect 18930 9808 18972 9848
rect 19012 9808 19054 9848
rect 19094 9808 19136 9848
rect 19176 9808 19185 9848
rect 19468 9764 19508 9892
rect 34348 9848 34388 9892
rect 18595 9724 18604 9764
rect 18644 9724 18653 9764
rect 18892 9724 19508 9764
rect 19852 9808 27532 9848
rect 27572 9808 27581 9848
rect 32323 9808 32332 9848
rect 32372 9808 32468 9848
rect 32995 9808 33004 9848
rect 33044 9808 33620 9848
rect 33919 9808 33928 9848
rect 33968 9808 34010 9848
rect 34050 9808 34092 9848
rect 34132 9808 34174 9848
rect 34214 9808 34256 9848
rect 34296 9808 34305 9848
rect 34348 9808 34964 9848
rect 0 9680 90 9700
rect 18604 9680 18644 9724
rect 0 9640 1420 9680
rect 1460 9640 1469 9680
rect 10963 9640 10972 9680
rect 11012 9640 11212 9680
rect 11252 9640 11261 9680
rect 11347 9640 11356 9680
rect 11396 9640 11596 9680
rect 11636 9640 11645 9680
rect 11731 9640 11740 9680
rect 11780 9640 11980 9680
rect 12020 9640 12029 9680
rect 12115 9640 12124 9680
rect 12164 9640 12364 9680
rect 12404 9640 12413 9680
rect 12499 9640 12508 9680
rect 12548 9640 12748 9680
rect 12788 9640 12797 9680
rect 12883 9640 12892 9680
rect 12932 9640 13132 9680
rect 13172 9640 13181 9680
rect 13267 9640 13276 9680
rect 13316 9640 13516 9680
rect 13556 9640 13565 9680
rect 13651 9640 13660 9680
rect 13700 9640 13900 9680
rect 13940 9640 13949 9680
rect 14035 9640 14044 9680
rect 14084 9640 14284 9680
rect 14324 9640 14333 9680
rect 14419 9640 14428 9680
rect 14468 9640 14668 9680
rect 14708 9640 14717 9680
rect 14803 9640 14812 9680
rect 14852 9640 15052 9680
rect 15092 9640 15101 9680
rect 15187 9640 15196 9680
rect 15236 9640 15436 9680
rect 15476 9640 15485 9680
rect 15571 9640 15580 9680
rect 15620 9640 15820 9680
rect 15860 9640 15869 9680
rect 15955 9640 15964 9680
rect 16004 9640 16204 9680
rect 16244 9640 16253 9680
rect 16339 9640 16348 9680
rect 16388 9640 16588 9680
rect 16628 9640 16637 9680
rect 16723 9640 16732 9680
rect 16772 9640 16972 9680
rect 17012 9640 17021 9680
rect 17107 9640 17116 9680
rect 17156 9640 17356 9680
rect 17396 9640 17405 9680
rect 17491 9640 17500 9680
rect 17540 9640 17740 9680
rect 17780 9640 17789 9680
rect 17875 9640 17884 9680
rect 17924 9640 18124 9680
rect 18164 9640 18173 9680
rect 18259 9640 18268 9680
rect 18308 9640 18508 9680
rect 18548 9640 18557 9680
rect 18604 9640 18652 9680
rect 18692 9640 18701 9680
rect 18787 9640 18796 9680
rect 18836 9640 18845 9680
rect 0 9620 90 9640
rect 18796 9596 18836 9640
rect 10339 9556 10348 9596
rect 10388 9556 12692 9596
rect 12652 9512 12692 9556
rect 16492 9556 18836 9596
rect 18892 9596 18932 9724
rect 19027 9640 19036 9680
rect 19076 9640 19372 9680
rect 19412 9640 19421 9680
rect 18892 9556 19220 9596
rect 19411 9556 19420 9596
rect 19460 9556 19660 9596
rect 19700 9556 19709 9596
rect 16492 9512 16532 9556
rect 19180 9512 19220 9556
rect 19852 9512 19892 9808
rect 32428 9764 32468 9808
rect 20803 9724 20812 9764
rect 20852 9724 21140 9764
rect 31939 9724 31948 9764
rect 31988 9724 32372 9764
rect 32428 9724 33140 9764
rect 21100 9680 21140 9724
rect 32332 9680 32372 9724
rect 33100 9680 33140 9724
rect 20105 9640 20188 9680
rect 20228 9640 20236 9680
rect 20276 9640 20285 9680
rect 20611 9640 20620 9680
rect 20660 9640 20668 9680
rect 20708 9640 20791 9680
rect 21100 9640 21436 9680
rect 21476 9640 21485 9680
rect 31171 9640 31180 9680
rect 31220 9640 31228 9680
rect 31268 9640 31351 9680
rect 31555 9640 31564 9680
rect 31604 9640 31996 9680
rect 32036 9640 32045 9680
rect 32332 9640 32764 9680
rect 32804 9640 32813 9680
rect 33100 9640 33148 9680
rect 33188 9640 33197 9680
rect 33580 9596 33620 9808
rect 33667 9640 33676 9680
rect 33716 9640 34684 9680
rect 34724 9640 34733 9680
rect 20275 9556 20284 9596
rect 20324 9556 20428 9596
rect 20468 9556 20477 9596
rect 20908 9556 28780 9596
rect 28820 9556 28829 9596
rect 31363 9556 31372 9596
rect 31412 9556 31612 9596
rect 31652 9556 31661 9596
rect 31747 9556 31756 9596
rect 31796 9556 32380 9596
rect 32420 9556 32429 9596
rect 32707 9556 32716 9596
rect 32756 9556 33524 9596
rect 33580 9556 33716 9596
rect 20908 9512 20948 9556
rect 33484 9512 33524 9556
rect 33676 9512 33716 9556
rect 34924 9512 34964 9808
rect 35788 9680 35828 9976
rect 46278 9956 46368 9976
rect 46278 9680 46368 9700
rect 35788 9640 36220 9680
rect 36260 9640 36269 9680
rect 43219 9640 43228 9680
rect 43268 9640 43372 9680
rect 43412 9640 43421 9680
rect 43529 9640 43612 9680
rect 43652 9640 43660 9680
rect 43700 9640 43709 9680
rect 43987 9640 43996 9680
rect 44036 9640 46368 9680
rect 46278 9620 46368 9640
rect 35011 9556 35020 9596
rect 35060 9556 36604 9596
rect 36644 9556 36653 9596
rect 36739 9556 36748 9596
rect 36788 9556 44948 9596
rect 44908 9512 44948 9556
rect 9475 9472 9484 9512
rect 9524 9472 10732 9512
rect 10772 9472 10781 9512
rect 11107 9472 11116 9512
rect 11156 9472 11165 9512
rect 11299 9472 11308 9512
rect 11348 9472 11500 9512
rect 11540 9472 11549 9512
rect 11875 9472 11884 9512
rect 11924 9472 11933 9512
rect 12259 9472 12268 9512
rect 12308 9472 12317 9512
rect 12643 9472 12652 9512
rect 12692 9472 12701 9512
rect 13027 9472 13036 9512
rect 13076 9472 13228 9512
rect 13268 9472 13277 9512
rect 13411 9472 13420 9512
rect 13460 9472 13469 9512
rect 13673 9472 13804 9512
rect 13844 9472 13853 9512
rect 14057 9472 14188 9512
rect 14228 9472 14237 9512
rect 14563 9472 14572 9512
rect 14612 9472 14621 9512
rect 14947 9472 14956 9512
rect 14996 9472 15052 9512
rect 15092 9472 15127 9512
rect 15331 9472 15340 9512
rect 15380 9472 15436 9512
rect 15476 9472 15511 9512
rect 15715 9472 15724 9512
rect 15764 9472 15895 9512
rect 16099 9472 16108 9512
rect 16148 9472 16157 9512
rect 16483 9472 16492 9512
rect 16532 9472 16541 9512
rect 16867 9472 16876 9512
rect 16916 9472 16972 9512
rect 17012 9472 17047 9512
rect 17251 9472 17260 9512
rect 17300 9472 17452 9512
rect 17492 9472 17501 9512
rect 17635 9472 17644 9512
rect 17684 9472 17815 9512
rect 18019 9472 18028 9512
rect 18068 9472 18199 9512
rect 18403 9472 18412 9512
rect 18452 9472 18461 9512
rect 18665 9472 18796 9512
rect 18836 9472 18845 9512
rect 19171 9472 19180 9512
rect 19220 9472 19229 9512
rect 19555 9472 19564 9512
rect 19604 9472 19892 9512
rect 19939 9472 19948 9512
rect 19988 9472 20468 9512
rect 20515 9472 20524 9512
rect 20564 9472 20573 9512
rect 20899 9472 20908 9512
rect 20948 9472 20957 9512
rect 21667 9472 21676 9512
rect 21716 9472 27340 9512
rect 27380 9472 27389 9512
rect 31337 9472 31468 9512
rect 31508 9472 31517 9512
rect 31651 9472 31660 9512
rect 31700 9472 31852 9512
rect 31892 9472 31901 9512
rect 32035 9472 32044 9512
rect 32084 9472 32236 9512
rect 32276 9472 32285 9512
rect 32611 9472 32620 9512
rect 32660 9472 32812 9512
rect 32852 9472 32861 9512
rect 32995 9472 33004 9512
rect 33044 9472 33053 9512
rect 33379 9472 33388 9512
rect 33428 9472 33437 9512
rect 33484 9472 33532 9512
rect 33572 9472 33581 9512
rect 33676 9472 33772 9512
rect 33812 9472 33821 9512
rect 33955 9472 33964 9512
rect 34004 9472 34156 9512
rect 34196 9472 34205 9512
rect 34531 9472 34540 9512
rect 34580 9472 34732 9512
rect 34772 9472 34781 9512
rect 34915 9472 34924 9512
rect 34964 9472 34973 9512
rect 35299 9472 35308 9512
rect 35348 9472 35357 9512
rect 35561 9472 35692 9512
rect 35732 9472 35741 9512
rect 35945 9472 36076 9512
rect 36116 9472 36125 9512
rect 36329 9472 36460 9512
rect 36500 9472 36509 9512
rect 36835 9472 36844 9512
rect 36884 9472 36893 9512
rect 37123 9472 37132 9512
rect 37172 9472 37708 9512
rect 37748 9472 37757 9512
rect 37891 9472 37900 9512
rect 37940 9472 38476 9512
rect 38516 9472 39052 9512
rect 39092 9472 39628 9512
rect 39668 9472 39916 9512
rect 39956 9472 40492 9512
rect 40532 9472 40780 9512
rect 40820 9472 40829 9512
rect 42857 9472 42988 9512
rect 43028 9472 43037 9512
rect 43241 9472 43372 9512
rect 43412 9472 43421 9512
rect 43625 9472 43756 9512
rect 43796 9472 43805 9512
rect 44131 9472 44140 9512
rect 44180 9472 44189 9512
rect 44236 9472 44524 9512
rect 44564 9472 44573 9512
rect 44899 9472 44908 9512
rect 44948 9472 44957 9512
rect 11116 9428 11156 9472
rect 11884 9428 11924 9472
rect 8611 9388 8620 9428
rect 8660 9388 11156 9428
rect 11203 9388 11212 9428
rect 11252 9388 11924 9428
rect 0 9344 90 9364
rect 12268 9344 12308 9472
rect 13420 9428 13460 9472
rect 13420 9388 14284 9428
rect 14324 9388 14333 9428
rect 0 9304 1420 9344
rect 1460 9304 1469 9344
rect 10147 9304 10156 9344
rect 10196 9304 12308 9344
rect 14572 9344 14612 9472
rect 16108 9428 16148 9472
rect 18412 9428 18452 9472
rect 16108 9388 17260 9428
rect 17300 9388 17309 9428
rect 18412 9388 19756 9428
rect 19796 9388 19805 9428
rect 19852 9388 20044 9428
rect 20084 9388 20093 9428
rect 19852 9344 19892 9388
rect 14572 9304 18028 9344
rect 18068 9304 18077 9344
rect 19795 9304 19804 9344
rect 19844 9304 19892 9344
rect 20428 9344 20468 9472
rect 20524 9428 20564 9472
rect 33004 9428 33044 9472
rect 20524 9388 28012 9428
rect 28052 9388 28061 9428
rect 32227 9388 32236 9428
rect 32276 9388 33044 9428
rect 33091 9388 33100 9428
rect 33140 9388 33149 9428
rect 33100 9344 33140 9388
rect 20428 9304 27916 9344
rect 27956 9304 27965 9344
rect 30883 9304 30892 9344
rect 30932 9304 33140 9344
rect 0 9284 90 9304
rect 18220 9220 20756 9260
rect 20969 9220 21004 9260
rect 21044 9220 21100 9260
rect 21140 9220 21149 9260
rect 32323 9220 32332 9260
rect 32372 9220 33004 9260
rect 33044 9220 33053 9260
rect 4919 9052 4928 9092
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 5296 9052 5305 9092
rect 0 9008 90 9028
rect 0 8968 1420 9008
rect 1460 8968 1469 9008
rect 9763 8968 9772 9008
rect 9812 8968 12980 9008
rect 0 8948 90 8968
rect 11011 8884 11020 8924
rect 11060 8884 11068 8924
rect 11108 8884 11191 8924
rect 11395 8884 11404 8924
rect 11444 8884 11452 8924
rect 11492 8884 11575 8924
rect 11779 8884 11788 8924
rect 11828 8884 11836 8924
rect 11876 8884 11959 8924
rect 12163 8884 12172 8924
rect 12212 8884 12220 8924
rect 12260 8884 12343 8924
rect 12547 8884 12556 8924
rect 12596 8884 12604 8924
rect 12644 8884 12727 8924
rect 10531 8800 10540 8840
rect 10580 8800 12884 8840
rect 8707 8716 8716 8756
rect 8756 8716 11444 8756
rect 11491 8716 11500 8756
rect 11540 8716 12116 8756
rect 0 8672 90 8692
rect 11404 8672 11444 8716
rect 12076 8672 12116 8716
rect 12844 8672 12884 8800
rect 12940 8672 12980 8968
rect 13315 8884 13324 8924
rect 13364 8884 13372 8924
rect 13412 8884 13495 8924
rect 13699 8884 13708 8924
rect 13748 8884 13756 8924
rect 13796 8884 13879 8924
rect 14083 8884 14092 8924
rect 14132 8884 14140 8924
rect 14180 8884 14263 8924
rect 14467 8884 14476 8924
rect 14516 8884 14524 8924
rect 14564 8884 14647 8924
rect 14851 8884 14860 8924
rect 14900 8884 14908 8924
rect 14948 8884 15031 8924
rect 15235 8884 15244 8924
rect 15284 8884 15292 8924
rect 15332 8884 15415 8924
rect 15619 8884 15628 8924
rect 15668 8884 15676 8924
rect 15716 8884 15799 8924
rect 16003 8884 16012 8924
rect 16052 8884 16060 8924
rect 16100 8884 16183 8924
rect 16387 8884 16396 8924
rect 16436 8884 16444 8924
rect 16484 8884 16567 8924
rect 16771 8884 16780 8924
rect 16820 8884 16828 8924
rect 16868 8884 16951 8924
rect 17155 8884 17164 8924
rect 17204 8884 17212 8924
rect 17252 8884 17335 8924
rect 17539 8884 17548 8924
rect 17588 8884 17596 8924
rect 17636 8884 17719 8924
rect 17923 8884 17932 8924
rect 17972 8884 17980 8924
rect 18020 8884 18103 8924
rect 13507 8716 13516 8756
rect 13556 8716 14804 8756
rect 14764 8672 14804 8716
rect 16300 8716 17164 8756
rect 17204 8716 17213 8756
rect 17452 8716 18124 8756
rect 18164 8716 18173 8756
rect 16300 8672 16340 8716
rect 17452 8672 17492 8716
rect 18220 8672 18260 9220
rect 19747 9136 19756 9176
rect 19796 9136 20620 9176
rect 20660 9136 20669 9176
rect 20716 9092 20756 9220
rect 33388 9176 33428 9472
rect 35308 9428 35348 9472
rect 36844 9428 36884 9472
rect 33475 9388 33484 9428
rect 33524 9388 35348 9428
rect 35587 9388 35596 9428
rect 35636 9388 36884 9428
rect 36931 9388 36940 9428
rect 36980 9388 43948 9428
rect 43988 9388 43997 9428
rect 44140 9344 44180 9472
rect 33571 9304 33580 9344
rect 33620 9304 34300 9344
rect 34340 9304 34349 9344
rect 34435 9304 34444 9344
rect 34484 9304 35836 9344
rect 35876 9304 35885 9344
rect 35971 9304 35980 9344
rect 36020 9304 44180 9344
rect 20803 9136 20812 9176
rect 20852 9136 26668 9176
rect 26708 9136 26717 9176
rect 27235 9136 27244 9176
rect 27284 9136 30604 9176
rect 30644 9136 30653 9176
rect 31747 9136 31756 9176
rect 31796 9136 33428 9176
rect 33484 9220 33916 9260
rect 33956 9220 33965 9260
rect 34444 9220 35068 9260
rect 35108 9220 35117 9260
rect 35212 9220 35452 9260
rect 35492 9220 35501 9260
rect 35779 9220 35788 9260
rect 35828 9220 37036 9260
rect 37076 9220 37085 9260
rect 37306 9220 37315 9260
rect 37355 9220 37364 9260
rect 33484 9092 33524 9220
rect 34444 9176 34484 9220
rect 35212 9176 35252 9220
rect 37324 9176 37364 9220
rect 37708 9220 37891 9260
rect 37931 9220 37940 9260
rect 37987 9220 37996 9260
rect 38036 9220 38188 9260
rect 38228 9220 38764 9260
rect 38804 9220 39331 9260
rect 39371 9220 39380 9260
rect 40073 9220 40204 9260
rect 40244 9220 40253 9260
rect 37708 9176 37748 9220
rect 44236 9176 44276 9472
rect 46278 9344 46368 9364
rect 44371 9304 44380 9344
rect 44420 9304 46368 9344
rect 46278 9284 46368 9304
rect 44755 9220 44764 9260
rect 44804 9220 44813 9260
rect 45139 9220 45148 9260
rect 45188 9220 45772 9260
rect 45812 9220 45821 9260
rect 33763 9136 33772 9176
rect 33812 9136 34484 9176
rect 34531 9136 34540 9176
rect 34580 9136 35252 9176
rect 36355 9136 36364 9176
rect 36404 9136 37748 9176
rect 37795 9136 37804 9176
rect 37844 9136 44276 9176
rect 44764 9092 44804 9220
rect 18883 9052 18892 9092
rect 18932 9052 19948 9092
rect 19988 9052 19997 9092
rect 20039 9052 20048 9092
rect 20088 9052 20130 9092
rect 20170 9052 20212 9092
rect 20252 9052 20294 9092
rect 20334 9052 20376 9092
rect 20416 9052 20425 9092
rect 20716 9052 21524 9092
rect 21667 9052 21676 9092
rect 21716 9052 25132 9092
rect 25172 9052 25181 9092
rect 27340 9052 30796 9092
rect 30836 9052 30845 9092
rect 31939 9052 31948 9092
rect 31988 9052 32812 9092
rect 32852 9052 32861 9092
rect 33187 9052 33196 9092
rect 33236 9052 33524 9092
rect 34435 9052 34444 9092
rect 34484 9052 35020 9092
rect 35060 9052 35069 9092
rect 35159 9052 35168 9092
rect 35208 9052 35250 9092
rect 35290 9052 35332 9092
rect 35372 9052 35414 9092
rect 35454 9052 35496 9092
rect 35536 9052 35545 9092
rect 37891 9052 37900 9092
rect 37940 9052 40052 9092
rect 40099 9052 40108 9092
rect 40148 9052 43220 9092
rect 44764 9052 45620 9092
rect 21484 9008 21524 9052
rect 18604 8968 21428 9008
rect 21484 8968 25172 9008
rect 18307 8884 18316 8924
rect 18356 8884 18364 8924
rect 18404 8884 18487 8924
rect 18604 8672 18644 8968
rect 18691 8884 18700 8924
rect 18740 8884 18748 8924
rect 18788 8884 18871 8924
rect 19123 8884 19132 8924
rect 19172 8884 19276 8924
rect 19316 8884 19325 8924
rect 19459 8884 19468 8924
rect 19508 8884 19516 8924
rect 19556 8884 19639 8924
rect 19843 8884 19852 8924
rect 19892 8884 19900 8924
rect 19940 8884 20023 8924
rect 21388 8840 21428 8968
rect 25132 8924 25172 8968
rect 21667 8884 21676 8924
rect 21716 8884 25036 8924
rect 25076 8884 25085 8924
rect 25132 8884 27196 8924
rect 27236 8884 27245 8924
rect 18988 8800 21332 8840
rect 21388 8800 25852 8840
rect 25892 8800 25901 8840
rect 26371 8800 26380 8840
rect 26420 8800 26428 8840
rect 26468 8800 26551 8840
rect 18988 8672 19028 8800
rect 21292 8756 21332 8800
rect 19372 8716 21236 8756
rect 21292 8716 24268 8756
rect 24308 8716 24317 8756
rect 26092 8716 27244 8756
rect 27284 8716 27293 8756
rect 19372 8672 19412 8716
rect 21196 8672 21236 8716
rect 26092 8672 26132 8716
rect 27340 8672 27380 9052
rect 27436 8968 30988 9008
rect 31028 8968 31037 9008
rect 32428 8968 39916 9008
rect 39956 8968 39965 9008
rect 27436 8672 27476 8968
rect 27523 8884 27532 8924
rect 27572 8884 27580 8924
rect 27620 8884 27703 8924
rect 27820 8884 28876 8924
rect 28916 8884 28925 8924
rect 32131 8884 32140 8924
rect 32180 8884 32188 8924
rect 32228 8884 32311 8924
rect 27820 8672 27860 8884
rect 32428 8840 32468 8968
rect 40012 8924 40052 9052
rect 43180 9008 43220 9052
rect 45580 9008 45620 9052
rect 46278 9008 46368 9028
rect 43180 8968 44948 9008
rect 45580 8968 46368 9008
rect 32515 8884 32524 8924
rect 32564 8884 32572 8924
rect 32612 8884 32695 8924
rect 32899 8884 32908 8924
rect 32948 8884 32956 8924
rect 32996 8884 33079 8924
rect 33283 8884 33292 8924
rect 33332 8884 33340 8924
rect 33380 8884 33463 8924
rect 34121 8884 34243 8924
rect 34292 8884 34301 8924
rect 34348 8884 34876 8924
rect 34916 8884 34925 8924
rect 35011 8884 35020 8924
rect 35060 8884 36460 8924
rect 36500 8884 36509 8924
rect 36556 8884 36748 8924
rect 36788 8884 36797 8924
rect 37097 8884 37219 8924
rect 37268 8884 37277 8924
rect 37673 8884 37756 8924
rect 37796 8884 37804 8924
rect 37844 8884 37853 8924
rect 37996 8884 39820 8924
rect 39860 8884 39869 8924
rect 39994 8884 40003 8924
rect 40043 8884 40052 8924
rect 40291 8884 40300 8924
rect 40340 8884 43756 8924
rect 43796 8884 43805 8924
rect 43987 8884 43996 8924
rect 44036 8884 44140 8924
rect 44180 8884 44189 8924
rect 44297 8884 44380 8924
rect 44420 8884 44428 8924
rect 44468 8884 44477 8924
rect 34348 8840 34388 8884
rect 36556 8840 36596 8884
rect 37996 8840 38036 8884
rect 27907 8800 27916 8840
rect 27956 8800 27964 8840
rect 28004 8800 28087 8840
rect 28291 8800 28300 8840
rect 28340 8800 29012 8840
rect 32083 8800 32092 8840
rect 32132 8800 32468 8840
rect 33187 8800 33196 8840
rect 33236 8800 33964 8840
rect 34004 8800 34013 8840
rect 34339 8800 34348 8840
rect 34388 8800 34397 8840
rect 34627 8800 34636 8840
rect 34676 8800 35260 8840
rect 35300 8800 35309 8840
rect 36307 8800 36316 8840
rect 36356 8800 36596 8840
rect 36691 8800 36700 8840
rect 36740 8800 38036 8840
rect 38131 8800 38140 8840
rect 38180 8800 43372 8840
rect 43412 8800 43421 8840
rect 28204 8716 28684 8756
rect 28724 8716 28733 8756
rect 28204 8672 28244 8716
rect 28972 8672 29012 8800
rect 29155 8716 29164 8756
rect 29204 8716 32468 8756
rect 33379 8716 33388 8756
rect 33428 8716 35540 8756
rect 32428 8672 32468 8716
rect 35500 8672 35540 8716
rect 35596 8716 35980 8756
rect 36020 8716 36029 8756
rect 36172 8716 36940 8756
rect 36980 8716 36989 8756
rect 37411 8716 37420 8756
rect 37460 8716 44564 8756
rect 0 8632 1420 8672
rect 1460 8632 1469 8672
rect 9091 8632 9100 8672
rect 9140 8632 11251 8672
rect 11291 8632 11300 8672
rect 11404 8632 11692 8672
rect 11732 8632 11741 8672
rect 12067 8632 12076 8672
rect 12116 8632 12125 8672
rect 12329 8632 12460 8672
rect 12500 8632 12509 8672
rect 12835 8632 12844 8672
rect 12884 8632 12893 8672
rect 12940 8632 13228 8672
rect 13268 8632 13277 8672
rect 13481 8632 13612 8672
rect 13652 8632 13661 8672
rect 13865 8632 13996 8672
rect 14036 8632 14045 8672
rect 14249 8632 14380 8672
rect 14420 8632 14429 8672
rect 14755 8632 14764 8672
rect 14804 8632 14813 8672
rect 15017 8632 15148 8672
rect 15188 8632 15197 8672
rect 15401 8632 15532 8672
rect 15572 8632 15581 8672
rect 15785 8632 15916 8672
rect 15956 8632 15965 8672
rect 16291 8632 16300 8672
rect 16340 8632 16349 8672
rect 16553 8632 16684 8672
rect 16724 8632 16733 8672
rect 16937 8632 17068 8672
rect 17108 8632 17117 8672
rect 17443 8632 17452 8672
rect 17492 8632 17501 8672
rect 17827 8632 17836 8672
rect 17876 8632 18164 8672
rect 18211 8632 18220 8672
rect 18260 8632 18269 8672
rect 18595 8632 18604 8672
rect 18644 8632 18653 8672
rect 18979 8632 18988 8672
rect 19028 8632 19037 8672
rect 19363 8632 19372 8672
rect 19412 8632 19421 8672
rect 19625 8632 19756 8672
rect 19796 8632 19805 8672
rect 20131 8632 20140 8672
rect 20180 8632 21140 8672
rect 21196 8632 25900 8672
rect 25940 8632 25949 8672
rect 26083 8632 26092 8672
rect 26132 8632 26141 8672
rect 26659 8632 26668 8672
rect 26708 8632 27380 8672
rect 27427 8632 27436 8672
rect 27476 8632 27485 8672
rect 27811 8632 27820 8672
rect 27860 8632 27869 8672
rect 28003 8632 28012 8672
rect 28052 8632 28148 8672
rect 28195 8632 28204 8672
rect 28244 8632 28253 8672
rect 28300 8632 28348 8672
rect 28388 8632 28397 8672
rect 28457 8632 28492 8672
rect 28532 8632 28588 8672
rect 28628 8632 28637 8672
rect 28723 8632 28732 8672
rect 28772 8632 28780 8672
rect 28820 8632 28903 8672
rect 28963 8632 28972 8672
rect 29012 8632 29021 8672
rect 30019 8632 30028 8672
rect 30068 8632 31604 8672
rect 31721 8632 31852 8672
rect 31892 8632 31901 8672
rect 32419 8632 32428 8672
rect 32468 8632 32477 8672
rect 32681 8632 32812 8672
rect 32852 8632 32861 8672
rect 32995 8632 33004 8672
rect 33044 8632 33196 8672
rect 33236 8632 33245 8672
rect 33292 8632 33580 8672
rect 33620 8632 33629 8672
rect 33737 8632 33868 8672
rect 33908 8632 33917 8672
rect 34217 8632 34252 8672
rect 34292 8632 34348 8672
rect 34388 8632 34540 8672
rect 34580 8632 34589 8672
rect 34723 8632 34732 8672
rect 34772 8632 35116 8672
rect 35156 8632 35165 8672
rect 35491 8632 35500 8672
rect 35540 8632 35549 8672
rect 0 8612 90 8632
rect 18124 8588 18164 8632
rect 21100 8588 21140 8632
rect 28108 8588 28148 8632
rect 28300 8588 28340 8632
rect 12979 8548 12988 8588
rect 13028 8548 13036 8588
rect 13076 8548 13159 8588
rect 18124 8548 20524 8588
rect 20564 8548 20573 8588
rect 21100 8548 21676 8588
rect 21716 8548 21725 8588
rect 28108 8548 28340 8588
rect 31564 8588 31604 8632
rect 31564 8548 33140 8588
rect 33100 8504 33140 8548
rect 33292 8504 33332 8632
rect 35596 8588 35636 8716
rect 35779 8632 35788 8672
rect 35828 8632 36076 8672
rect 36116 8632 36125 8672
rect 34771 8548 34780 8588
rect 34820 8548 35636 8588
rect 36172 8504 36212 8716
rect 44524 8672 44564 8716
rect 44908 8672 44948 8968
rect 46278 8948 46368 8968
rect 46278 8672 46368 8692
rect 36355 8632 36364 8672
rect 36404 8632 36460 8672
rect 36500 8632 36844 8672
rect 36884 8632 36893 8672
rect 37219 8632 37228 8672
rect 37268 8632 37516 8672
rect 37556 8632 37565 8672
rect 37769 8632 37900 8672
rect 37940 8632 37949 8672
rect 38275 8632 38284 8672
rect 38324 8632 38572 8672
rect 38612 8632 38668 8672
rect 38708 8632 38860 8672
rect 38900 8632 39148 8672
rect 39188 8632 39436 8672
rect 39476 8632 39724 8672
rect 39764 8632 40204 8672
rect 40244 8632 40300 8672
rect 40340 8632 40375 8672
rect 40483 8632 40492 8672
rect 40532 8632 43756 8672
rect 43796 8632 43805 8672
rect 43939 8632 43948 8672
rect 43988 8632 44140 8672
rect 44180 8632 44189 8672
rect 44515 8632 44524 8672
rect 44564 8632 44573 8672
rect 44899 8632 44908 8672
rect 44948 8632 44957 8672
rect 45763 8632 45772 8672
rect 45812 8632 46368 8672
rect 16771 8464 16780 8504
rect 16820 8464 22540 8504
rect 22580 8464 22589 8504
rect 26188 8464 29836 8504
rect 29876 8464 29885 8504
rect 33100 8464 33332 8504
rect 34099 8464 34108 8504
rect 34148 8464 36212 8504
rect 37516 8504 37556 8632
rect 38284 8504 38324 8632
rect 46278 8612 46368 8632
rect 37516 8464 38324 8504
rect 44755 8464 44764 8504
rect 44804 8464 44813 8504
rect 45139 8464 45148 8504
rect 45188 8464 45772 8504
rect 45812 8464 45821 8504
rect 26188 8420 26228 8464
rect 2947 8380 2956 8420
rect 2996 8380 12980 8420
rect 26179 8380 26188 8420
rect 26228 8380 26237 8420
rect 26563 8380 26572 8420
rect 26612 8380 30412 8420
rect 30452 8380 30461 8420
rect 0 8336 90 8356
rect 0 8296 172 8336
rect 212 8296 221 8336
rect 3679 8296 3688 8336
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 4056 8296 4065 8336
rect 0 8276 90 8296
rect 1315 8212 1324 8252
rect 1364 8212 10100 8252
rect 652 8128 2860 8168
rect 2900 8128 2909 8168
rect 652 8084 692 8128
rect 268 8044 692 8084
rect 10060 8084 10100 8212
rect 12940 8168 12980 8380
rect 44764 8336 44804 8464
rect 46278 8336 46368 8356
rect 18799 8296 18808 8336
rect 18848 8296 18890 8336
rect 18930 8296 18972 8336
rect 19012 8296 19054 8336
rect 19094 8296 19136 8336
rect 19176 8296 19185 8336
rect 26947 8296 26956 8336
rect 26996 8296 29452 8336
rect 29492 8296 29501 8336
rect 33919 8296 33928 8336
rect 33968 8296 34010 8336
rect 34050 8296 34092 8336
rect 34132 8296 34174 8336
rect 34214 8296 34256 8336
rect 34296 8296 34305 8336
rect 44764 8296 46368 8336
rect 46278 8276 46368 8296
rect 16579 8212 16588 8252
rect 16628 8212 22732 8252
rect 22772 8212 22781 8252
rect 23020 8212 31852 8252
rect 31892 8212 31901 8252
rect 23020 8168 23060 8212
rect 12940 8128 23060 8168
rect 24259 8128 24268 8168
rect 24308 8128 25564 8168
rect 25604 8128 25613 8168
rect 25891 8128 25900 8168
rect 25940 8128 25948 8168
rect 25988 8128 26071 8168
rect 26659 8128 26668 8168
rect 26708 8128 26716 8168
rect 26756 8128 26839 8168
rect 27043 8128 27052 8168
rect 27092 8128 27100 8168
rect 27140 8128 27223 8168
rect 32947 8128 32956 8168
rect 32996 8128 39668 8168
rect 39763 8128 39772 8168
rect 39812 8128 40492 8168
rect 40532 8128 40541 8168
rect 42979 8128 42988 8168
rect 43028 8128 43132 8168
rect 43172 8128 43181 8168
rect 39628 8084 39668 8128
rect 10060 8044 20140 8084
rect 20180 8044 20189 8084
rect 20899 8044 20908 8084
rect 20948 8044 26332 8084
rect 26372 8044 26381 8084
rect 27523 8044 27532 8084
rect 27572 8044 39572 8084
rect 39628 8044 44948 8084
rect 0 8000 90 8020
rect 268 8000 308 8044
rect 39532 8000 39572 8044
rect 44908 8000 44948 8044
rect 46278 8000 46368 8020
rect 0 7960 308 8000
rect 13699 7960 13708 8000
rect 13748 7960 24844 8000
rect 24884 7960 24893 8000
rect 25123 7960 25132 8000
rect 25172 7960 25180 8000
rect 25220 7960 25303 8000
rect 25411 7960 25420 8000
rect 25460 7960 25591 8000
rect 25795 7960 25804 8000
rect 25844 7960 25900 8000
rect 25940 7960 25975 8000
rect 26179 7960 26188 8000
rect 26228 7960 26359 8000
rect 26441 7960 26572 8000
rect 26612 7960 26621 8000
rect 26825 7960 26956 8000
rect 26996 7960 27005 8000
rect 27209 7960 27244 8000
rect 27284 7960 27340 8000
rect 27380 7960 27389 8000
rect 27475 7960 27484 8000
rect 27524 7960 27572 8000
rect 27715 7960 27724 8000
rect 27764 7960 27773 8000
rect 28073 7960 28108 8000
rect 28148 7960 28204 8000
rect 28244 7960 28253 8000
rect 32585 7960 32716 8000
rect 32756 7960 32765 8000
rect 34217 7960 34348 8000
rect 34388 7960 34636 8000
rect 34676 7960 34924 8000
rect 34964 7960 35212 8000
rect 35252 7960 35500 8000
rect 35540 7960 35788 8000
rect 35828 7960 36076 8000
rect 36116 7960 36172 8000
rect 36212 7960 36276 8000
rect 36329 7960 36460 8000
rect 36500 7960 36509 8000
rect 36691 7960 36700 8000
rect 36740 7960 37420 8000
rect 37460 7960 37469 8000
rect 37891 7960 37900 8000
rect 37940 7960 38380 8000
rect 38420 7960 38429 8000
rect 38537 7960 38668 8000
rect 38708 7960 38717 8000
rect 39523 7960 39532 8000
rect 39572 7960 39581 8000
rect 43363 7960 43372 8000
rect 43412 7960 43421 8000
rect 43555 7960 43564 8000
rect 43604 7960 44524 8000
rect 44564 7960 44573 8000
rect 44899 7960 44908 8000
rect 44948 7960 44957 8000
rect 45763 7960 45772 8000
rect 45812 7960 46368 8000
rect 0 7940 90 7960
rect 27532 7916 27572 7960
rect 259 7876 268 7916
rect 308 7876 10100 7916
rect 25027 7876 25036 7916
rect 25076 7876 27572 7916
rect 27724 7916 27764 7960
rect 27724 7876 29068 7916
rect 29108 7876 29117 7916
rect 36809 7876 36940 7916
rect 36980 7876 37132 7916
rect 37172 7876 37181 7916
rect 10060 7748 10100 7876
rect 43372 7832 43412 7960
rect 46278 7940 46368 7960
rect 23020 7792 35212 7832
rect 35252 7792 35261 7832
rect 40291 7792 40300 7832
rect 40340 7792 43412 7832
rect 23020 7748 23060 7792
rect 10060 7708 23060 7748
rect 27331 7708 27340 7748
rect 27380 7708 27964 7748
rect 28004 7708 28013 7748
rect 37228 7708 37411 7748
rect 37451 7708 37699 7748
rect 37739 7708 37987 7748
rect 38027 7708 38036 7748
rect 44755 7708 44764 7748
rect 44804 7708 44813 7748
rect 45139 7708 45148 7748
rect 45188 7708 45772 7748
rect 45812 7708 45821 7748
rect 0 7664 90 7684
rect 0 7624 4780 7664
rect 4820 7624 4829 7664
rect 5539 7624 5548 7664
rect 5588 7624 35692 7664
rect 35732 7624 35741 7664
rect 0 7604 90 7624
rect 4919 7540 4928 7580
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 5296 7540 5305 7580
rect 20039 7540 20048 7580
rect 20088 7540 20130 7580
rect 20170 7540 20212 7580
rect 20252 7540 20294 7580
rect 20334 7540 20376 7580
rect 20416 7540 20425 7580
rect 25891 7540 25900 7580
rect 25940 7540 30220 7580
rect 30260 7540 30269 7580
rect 35159 7540 35168 7580
rect 35208 7540 35250 7580
rect 35290 7540 35332 7580
rect 35372 7540 35414 7580
rect 35454 7540 35496 7580
rect 35536 7540 35545 7580
rect 163 7456 172 7496
rect 212 7456 36460 7496
rect 36500 7456 36509 7496
rect 37228 7412 37268 7708
rect 44764 7664 44804 7708
rect 46278 7664 46368 7684
rect 44764 7624 46368 7664
rect 46278 7604 46368 7624
rect 25411 7372 25420 7412
rect 25460 7372 29932 7412
rect 29972 7372 29981 7412
rect 35945 7372 36076 7412
rect 36116 7372 37268 7412
rect 0 7328 90 7348
rect 46278 7328 46368 7348
rect 0 7288 32716 7328
rect 32756 7288 32765 7328
rect 45763 7288 45772 7328
rect 45812 7288 46368 7328
rect 0 7268 90 7288
rect 46278 7268 46368 7288
rect 36076 7204 36308 7244
rect 36076 7160 36116 7204
rect 8323 7120 8332 7160
rect 8372 7120 21196 7160
rect 21236 7120 21245 7160
rect 25891 7120 25900 7160
rect 25940 7120 29644 7160
rect 29684 7120 29693 7160
rect 33161 7120 33292 7160
rect 33332 7120 33341 7160
rect 35561 7120 35692 7160
rect 35732 7120 35741 7160
rect 35923 7120 35932 7160
rect 35972 7120 36116 7160
rect 36268 7160 36308 7204
rect 36268 7120 43564 7160
rect 43604 7120 43613 7160
rect 44393 7120 44524 7160
rect 44564 7120 44573 7160
rect 44899 7120 44908 7160
rect 44948 7120 44957 7160
rect 44908 7076 44948 7120
rect 8489 7036 8572 7076
rect 8612 7036 8620 7076
rect 8660 7036 8669 7076
rect 12940 7036 32044 7076
rect 32084 7036 32093 7076
rect 33523 7036 33532 7076
rect 33572 7036 44948 7076
rect 0 6992 90 7012
rect 12940 6992 12980 7036
rect 46278 6992 46368 7012
rect 0 6952 7852 6992
rect 7892 6952 7901 6992
rect 8035 6952 8044 6992
rect 8084 6952 12980 6992
rect 18691 6952 18700 6992
rect 18740 6952 25660 6992
rect 25700 6952 25709 6992
rect 44755 6952 44764 6992
rect 44804 6952 45044 6992
rect 45139 6952 45148 6992
rect 45188 6952 46368 6992
rect 0 6932 90 6952
rect 15811 6868 15820 6908
rect 15860 6868 24076 6908
rect 24116 6868 24125 6908
rect 3679 6784 3688 6824
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 4056 6784 4065 6824
rect 8803 6784 8812 6824
rect 8852 6784 15340 6824
rect 15380 6784 15389 6824
rect 18799 6784 18808 6824
rect 18848 6784 18890 6824
rect 18930 6784 18972 6824
rect 19012 6784 19054 6824
rect 19094 6784 19136 6824
rect 19176 6784 19185 6824
rect 19843 6784 19852 6824
rect 19892 6784 21388 6824
rect 21428 6784 21437 6824
rect 33919 6784 33928 6824
rect 33968 6784 34010 6824
rect 34050 6784 34092 6824
rect 34132 6784 34174 6824
rect 34214 6784 34256 6824
rect 34296 6784 34305 6824
rect 2860 6700 12980 6740
rect 16867 6700 16876 6740
rect 16916 6700 21580 6740
rect 21620 6700 21629 6740
rect 0 6656 90 6676
rect 2860 6656 2900 6700
rect 12940 6656 12980 6700
rect 45004 6656 45044 6952
rect 46278 6932 46368 6952
rect 46278 6656 46368 6676
rect 0 6616 2900 6656
rect 7603 6616 7612 6656
rect 7652 6616 8044 6656
rect 8084 6616 8093 6656
rect 12940 6616 33140 6656
rect 45004 6616 46368 6656
rect 0 6596 90 6616
rect 8585 6532 8668 6572
rect 8708 6532 8716 6572
rect 8756 6532 8765 6572
rect 8969 6532 9052 6572
rect 9092 6532 9100 6572
rect 9140 6532 9149 6572
rect 9353 6532 9436 6572
rect 9476 6532 9484 6572
rect 9524 6532 9533 6572
rect 13939 6532 13948 6572
rect 13988 6532 14188 6572
rect 14228 6532 14237 6572
rect 15523 6532 15532 6572
rect 15572 6532 19132 6572
rect 19172 6532 19181 6572
rect 19276 6532 23500 6572
rect 23540 6532 23549 6572
rect 19276 6488 19316 6532
rect 33100 6488 33140 6616
rect 46278 6596 46368 6616
rect 6211 6448 6220 6488
rect 6260 6448 7372 6488
rect 7412 6448 7421 6488
rect 7747 6448 7756 6488
rect 7796 6448 7805 6488
rect 8297 6448 8428 6488
rect 8468 6448 8477 6488
rect 8681 6448 8812 6488
rect 8852 6448 8861 6488
rect 9187 6448 9196 6488
rect 9236 6448 12980 6488
rect 13699 6448 13708 6488
rect 13748 6448 19316 6488
rect 19363 6448 19372 6488
rect 19412 6448 19543 6488
rect 19660 6448 19804 6488
rect 19844 6448 19853 6488
rect 20035 6448 20044 6488
rect 20084 6448 20093 6488
rect 20419 6448 20428 6488
rect 20468 6448 26476 6488
rect 26516 6448 26525 6488
rect 33100 6448 33772 6488
rect 33812 6448 33821 6488
rect 35683 6448 35692 6488
rect 35732 6448 35788 6488
rect 35828 6448 35980 6488
rect 36020 6448 36029 6488
rect 41731 6448 41740 6488
rect 41780 6448 44524 6488
rect 44564 6448 44573 6488
rect 44777 6448 44908 6488
rect 44948 6448 44957 6488
rect 7756 6404 7796 6448
rect 4099 6364 4108 6404
rect 4148 6364 7796 6404
rect 12940 6404 12980 6448
rect 19660 6404 19700 6448
rect 12940 6364 16876 6404
rect 16916 6364 16925 6404
rect 17059 6364 17068 6404
rect 17108 6364 19700 6404
rect 20044 6404 20084 6448
rect 20044 6364 25996 6404
rect 26036 6364 26045 6404
rect 0 6320 90 6340
rect 46278 6320 46368 6340
rect 0 6280 748 6320
rect 788 6280 797 6320
rect 7987 6280 7996 6320
rect 8036 6280 31660 6320
rect 31700 6280 31709 6320
rect 45139 6280 45148 6320
rect 45188 6280 46368 6320
rect 0 6260 90 6280
rect 46278 6260 46368 6280
rect 15715 6196 15724 6236
rect 15764 6196 20188 6236
rect 20228 6196 20237 6236
rect 34003 6196 34012 6236
rect 34052 6196 35636 6236
rect 44755 6196 44764 6236
rect 44804 6196 46100 6236
rect 35596 6152 35636 6196
rect 46060 6152 46100 6196
rect 19363 6112 19372 6152
rect 19412 6112 21964 6152
rect 22004 6112 22013 6152
rect 35596 6112 44524 6152
rect 44564 6112 44573 6152
rect 46060 6112 46252 6152
rect 46292 6112 46301 6152
rect 4919 6028 4928 6068
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 5296 6028 5305 6068
rect 8419 6028 8428 6068
rect 8468 6028 19852 6068
rect 19892 6028 19901 6068
rect 20039 6028 20048 6068
rect 20088 6028 20130 6068
rect 20170 6028 20212 6068
rect 20252 6028 20294 6068
rect 20334 6028 20376 6068
rect 20416 6028 20425 6068
rect 24835 6028 24844 6068
rect 24884 6028 27436 6068
rect 27476 6028 27485 6068
rect 35159 6028 35168 6068
rect 35208 6028 35250 6068
rect 35290 6028 35332 6068
rect 35372 6028 35414 6068
rect 35454 6028 35496 6068
rect 35536 6028 35545 6068
rect 0 5984 90 6004
rect 46278 5984 46368 6004
rect 0 5944 34444 5984
rect 34484 5944 34493 5984
rect 46243 5944 46252 5984
rect 46292 5944 46368 5984
rect 0 5924 90 5944
rect 46278 5924 46368 5944
rect 7843 5860 7852 5900
rect 7892 5860 33292 5900
rect 33332 5860 33341 5900
rect 14092 5776 15820 5816
rect 15860 5776 15869 5816
rect 18019 5776 18028 5816
rect 18068 5776 18268 5816
rect 18308 5776 18317 5816
rect 18521 5776 18604 5816
rect 18644 5776 18652 5816
rect 18692 5776 18701 5816
rect 18796 5776 19036 5816
rect 19076 5776 19085 5816
rect 21388 5776 21908 5816
rect 21955 5776 21964 5816
rect 22004 5776 24844 5816
rect 24884 5776 24893 5816
rect 25027 5776 25036 5816
rect 25076 5776 25364 5816
rect 0 5648 90 5668
rect 14092 5648 14132 5776
rect 18796 5732 18836 5776
rect 21388 5732 21428 5776
rect 21868 5732 21908 5776
rect 25324 5732 25364 5776
rect 14275 5692 14284 5732
rect 14324 5692 15092 5732
rect 15139 5692 15148 5732
rect 15188 5692 16532 5732
rect 17251 5692 17260 5732
rect 17300 5692 18836 5732
rect 18892 5692 20044 5732
rect 20084 5692 20093 5732
rect 20236 5692 20524 5732
rect 20564 5692 20573 5732
rect 21100 5692 21428 5732
rect 21484 5692 21812 5732
rect 21868 5692 23020 5732
rect 23060 5692 23069 5732
rect 23116 5692 25228 5732
rect 25268 5692 25277 5732
rect 25324 5692 26860 5732
rect 26900 5692 26909 5732
rect 27331 5692 27340 5732
rect 27380 5692 29492 5732
rect 29539 5692 29548 5732
rect 29588 5692 30356 5732
rect 15052 5648 15092 5692
rect 16492 5648 16532 5692
rect 18892 5648 18932 5692
rect 0 5608 1420 5648
rect 1460 5608 1469 5648
rect 1987 5608 1996 5648
rect 2036 5608 9100 5648
rect 9140 5608 9149 5648
rect 9475 5608 9484 5648
rect 9524 5608 9580 5648
rect 9620 5608 9655 5648
rect 9737 5608 9868 5648
rect 9908 5608 9917 5648
rect 10121 5608 10252 5648
rect 10292 5608 10301 5648
rect 10505 5608 10636 5648
rect 10676 5608 10685 5648
rect 10889 5608 11020 5648
rect 11060 5608 11069 5648
rect 11299 5608 11308 5648
rect 11348 5608 11356 5648
rect 11396 5608 11479 5648
rect 11587 5608 11596 5648
rect 11636 5608 11767 5648
rect 11818 5608 11827 5648
rect 11867 5608 11884 5648
rect 11924 5608 12007 5648
rect 13219 5608 13228 5648
rect 13268 5608 13324 5648
rect 13364 5608 13399 5648
rect 13481 5608 13564 5648
rect 13604 5608 13612 5648
rect 13652 5608 13661 5648
rect 13795 5608 13804 5648
rect 13844 5608 13853 5648
rect 13987 5608 13996 5648
rect 14036 5608 14132 5648
rect 14227 5608 14236 5648
rect 14276 5608 14380 5648
rect 14420 5608 14429 5648
rect 14563 5608 14572 5648
rect 14612 5608 14668 5648
rect 14708 5608 14743 5648
rect 14825 5608 14956 5648
rect 14996 5608 15005 5648
rect 15052 5608 15100 5648
rect 15140 5608 15149 5648
rect 15331 5608 15340 5648
rect 15380 5608 15511 5648
rect 16492 5608 17884 5648
rect 17924 5608 17933 5648
rect 18115 5608 18124 5648
rect 18164 5608 18295 5648
rect 18499 5608 18508 5648
rect 18548 5608 18679 5648
rect 18883 5608 18892 5648
rect 18932 5608 18941 5648
rect 19145 5608 19276 5648
rect 19316 5608 19325 5648
rect 19529 5608 19660 5648
rect 19700 5608 19709 5648
rect 20035 5608 20044 5648
rect 20084 5608 20093 5648
rect 0 5588 90 5608
rect 13804 5564 13844 5608
rect 9641 5524 9724 5564
rect 9764 5524 9772 5564
rect 9812 5524 9821 5564
rect 10025 5524 10108 5564
rect 10148 5524 10156 5564
rect 10196 5524 10205 5564
rect 10409 5524 10492 5564
rect 10532 5524 10540 5564
rect 10580 5524 10589 5564
rect 11251 5524 11260 5564
rect 11300 5524 11500 5564
rect 11540 5524 11549 5564
rect 12019 5524 12028 5564
rect 12068 5524 12460 5564
rect 12500 5524 12509 5564
rect 13385 5524 13468 5564
rect 13508 5524 13516 5564
rect 13556 5524 13565 5564
rect 13699 5524 13708 5564
rect 13748 5524 13844 5564
rect 13987 5524 13996 5564
rect 14036 5524 14332 5564
rect 14372 5524 14381 5564
rect 17932 5524 19852 5564
rect 19892 5524 19901 5564
rect 9331 5440 9340 5480
rect 9380 5440 9620 5480
rect 10867 5440 10876 5480
rect 10916 5440 11212 5480
rect 11252 5440 11261 5480
rect 13219 5440 13228 5480
rect 13268 5440 14716 5480
rect 14756 5440 14765 5480
rect 14851 5440 14860 5480
rect 14900 5440 16492 5480
rect 16532 5440 16541 5480
rect 9580 5396 9620 5440
rect 17932 5396 17972 5524
rect 20044 5480 20084 5608
rect 20236 5564 20276 5692
rect 21100 5648 21140 5692
rect 20419 5608 20428 5648
rect 20468 5608 20477 5648
rect 20803 5608 20812 5648
rect 20852 5608 21140 5648
rect 21187 5608 21196 5648
rect 21236 5608 21367 5648
rect 20179 5524 20188 5564
rect 20228 5524 20276 5564
rect 20428 5564 20468 5608
rect 21484 5564 21524 5692
rect 21772 5648 21812 5692
rect 23116 5648 23156 5692
rect 29452 5648 29492 5692
rect 30316 5648 30356 5692
rect 33100 5692 34484 5732
rect 33100 5648 33140 5692
rect 21571 5608 21580 5648
rect 21620 5608 21629 5648
rect 21772 5608 23156 5648
rect 23203 5608 23212 5648
rect 23252 5608 27340 5648
rect 27380 5608 27389 5648
rect 29443 5608 29452 5648
rect 29492 5608 29501 5648
rect 29705 5608 29836 5648
rect 29876 5608 29885 5648
rect 30019 5608 30028 5648
rect 30068 5608 30076 5648
rect 30116 5608 30199 5648
rect 30250 5608 30259 5648
rect 30299 5608 30356 5648
rect 30595 5608 30604 5648
rect 30644 5608 31564 5648
rect 31604 5608 31613 5648
rect 31913 5608 32044 5648
rect 32084 5608 32093 5648
rect 32419 5608 32428 5648
rect 32468 5608 32948 5648
rect 32995 5608 33004 5648
rect 33044 5608 33140 5648
rect 33235 5608 33244 5648
rect 33284 5608 33388 5648
rect 33428 5608 33437 5648
rect 33763 5608 33772 5648
rect 33812 5608 33964 5648
rect 34004 5608 34013 5648
rect 34195 5608 34204 5648
rect 34244 5608 34348 5648
rect 34388 5608 34397 5648
rect 20428 5524 21524 5564
rect 21580 5480 21620 5608
rect 32908 5564 32948 5608
rect 21763 5524 21772 5564
rect 21812 5524 31468 5564
rect 31508 5524 31517 5564
rect 32275 5524 32284 5564
rect 32324 5524 32852 5564
rect 32908 5524 33908 5564
rect 32812 5480 32852 5524
rect 18796 5440 19420 5480
rect 19460 5440 19469 5480
rect 19564 5440 19804 5480
rect 19844 5440 19853 5480
rect 19948 5440 20084 5480
rect 20419 5440 20428 5480
rect 20468 5440 20572 5480
rect 20612 5440 20621 5480
rect 20707 5440 20716 5480
rect 20756 5440 20956 5480
rect 20996 5440 21005 5480
rect 21283 5440 21292 5480
rect 21332 5440 21340 5480
rect 21380 5440 21463 5480
rect 21580 5440 23020 5480
rect 23060 5440 23069 5480
rect 23299 5440 23308 5480
rect 23348 5440 25324 5480
rect 25364 5440 25373 5480
rect 27571 5440 27580 5480
rect 27620 5440 29588 5480
rect 29683 5440 29692 5480
rect 29732 5440 29932 5480
rect 29972 5440 29981 5480
rect 30377 5440 30460 5480
rect 30500 5440 30508 5480
rect 30548 5440 30557 5480
rect 30761 5440 30844 5480
rect 30884 5440 30892 5480
rect 30932 5440 30941 5480
rect 32537 5440 32620 5480
rect 32660 5440 32668 5480
rect 32708 5440 32717 5480
rect 32812 5440 33716 5480
rect 18796 5396 18836 5440
rect 19564 5396 19604 5440
rect 9580 5356 17972 5396
rect 18499 5356 18508 5396
rect 18548 5356 18836 5396
rect 19372 5356 19604 5396
rect 0 5312 90 5332
rect 0 5272 652 5312
rect 692 5272 701 5312
rect 3679 5272 3688 5312
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 4056 5272 4065 5312
rect 10243 5272 10252 5312
rect 10292 5272 15284 5312
rect 18799 5272 18808 5312
rect 18848 5272 18890 5312
rect 18930 5272 18972 5312
rect 19012 5272 19054 5312
rect 19094 5272 19136 5312
rect 19176 5272 19185 5312
rect 0 5252 90 5272
rect 15244 5144 15284 5272
rect 19372 5144 19412 5356
rect 19948 5312 19988 5440
rect 29548 5396 29588 5440
rect 20035 5356 20044 5396
rect 20084 5356 25036 5396
rect 25076 5356 25085 5396
rect 25132 5356 26764 5396
rect 26804 5356 26813 5396
rect 29548 5356 33100 5396
rect 33140 5356 33149 5396
rect 19948 5272 24940 5312
rect 24980 5272 24989 5312
rect 25132 5228 25172 5356
rect 25219 5272 25228 5312
rect 25268 5272 29836 5312
rect 29876 5272 29885 5312
rect 33676 5228 33716 5440
rect 33868 5396 33908 5524
rect 34444 5480 34484 5692
rect 34636 5692 44236 5732
rect 44276 5692 44285 5732
rect 34636 5648 34676 5692
rect 46278 5648 46368 5668
rect 34627 5608 34636 5648
rect 34676 5608 34685 5648
rect 34867 5608 34876 5648
rect 34916 5608 35596 5648
rect 35636 5608 35645 5648
rect 40771 5608 40780 5648
rect 40820 5608 44524 5648
rect 44564 5608 44573 5648
rect 44899 5608 44908 5648
rect 44948 5608 44957 5648
rect 45139 5608 45148 5648
rect 45188 5608 46368 5648
rect 44908 5564 44948 5608
rect 46278 5588 46368 5608
rect 43267 5524 43276 5564
rect 43316 5524 44948 5564
rect 34444 5440 40012 5480
rect 40052 5440 40061 5480
rect 44755 5440 44764 5480
rect 44804 5440 46252 5480
rect 46292 5440 46301 5480
rect 33868 5356 37900 5396
rect 37940 5356 37949 5396
rect 46278 5312 46368 5332
rect 33919 5272 33928 5312
rect 33968 5272 34010 5312
rect 34050 5272 34092 5312
rect 34132 5272 34174 5312
rect 34214 5272 34256 5312
rect 34296 5272 34305 5312
rect 46243 5272 46252 5312
rect 46292 5272 46368 5312
rect 46278 5252 46368 5272
rect 21187 5188 21196 5228
rect 21236 5188 25172 5228
rect 25900 5188 26284 5228
rect 26324 5188 26333 5228
rect 33676 5188 44908 5228
rect 44948 5188 44957 5228
rect 10099 5104 10108 5144
rect 10148 5104 10348 5144
rect 10388 5104 10397 5144
rect 13795 5104 13804 5144
rect 13844 5104 13948 5144
rect 13988 5104 13997 5144
rect 15244 5104 16780 5144
rect 16820 5104 16829 5144
rect 17443 5104 17452 5144
rect 17492 5104 19412 5144
rect 19660 5104 20188 5144
rect 20228 5104 20237 5144
rect 20332 5104 21620 5144
rect 22339 5104 22348 5144
rect 22388 5104 25612 5144
rect 25652 5104 25661 5144
rect 19660 5060 19700 5104
rect 11587 5020 11596 5060
rect 11636 5020 16108 5060
rect 16148 5020 16157 5060
rect 16675 5020 16684 5060
rect 16724 5020 19700 5060
rect 19795 5020 19804 5060
rect 19844 5020 19948 5060
rect 19988 5020 19997 5060
rect 0 4976 90 4996
rect 20332 4976 20372 5104
rect 21580 4976 21620 5104
rect 25900 5060 25940 5188
rect 21667 5020 21676 5060
rect 21716 5020 25940 5060
rect 25996 5104 32044 5144
rect 32084 5104 32093 5144
rect 32275 5104 32284 5144
rect 32324 5104 34732 5144
rect 34772 5104 34781 5144
rect 0 4936 1132 4976
rect 1172 4936 1181 4976
rect 8323 4936 8332 4976
rect 8372 4936 8524 4976
rect 8564 4936 8573 4976
rect 9859 4936 9868 4976
rect 9908 4936 10060 4976
rect 10100 4936 10109 4976
rect 11011 4936 11020 4976
rect 11060 4936 13900 4976
rect 13940 4936 13949 4976
rect 14057 4936 14188 4976
rect 14228 4936 14237 4976
rect 15907 4936 15916 4976
rect 15956 4936 19180 4976
rect 19220 4936 19229 4976
rect 19433 4936 19564 4976
rect 19604 4936 19613 4976
rect 20035 4936 20044 4976
rect 20084 4936 20372 4976
rect 20419 4936 20428 4976
rect 20468 4936 21484 4976
rect 21524 4936 21533 4976
rect 21580 4936 25708 4976
rect 25748 4936 25757 4976
rect 0 4916 90 4936
rect 25996 4892 26036 5104
rect 29923 5020 29932 5060
rect 29972 5020 34828 5060
rect 34868 5020 34877 5060
rect 46278 4976 46368 4996
rect 26083 4936 26092 4976
rect 26132 4936 26141 4976
rect 31651 4936 31660 4976
rect 31700 4936 31709 4976
rect 32035 4936 32044 4976
rect 32084 4936 35788 4976
rect 35828 4936 35837 4976
rect 40867 4936 40876 4976
rect 40916 4936 44524 4976
rect 44564 4936 44573 4976
rect 44899 4936 44908 4976
rect 44948 4936 44957 4976
rect 45139 4936 45148 4976
rect 45188 4936 46368 4976
rect 739 4852 748 4892
rect 788 4852 26036 4892
rect 10627 4768 10636 4808
rect 10676 4768 13172 4808
rect 15043 4768 15052 4808
rect 15092 4768 19324 4808
rect 19364 4768 19373 4808
rect 19651 4768 19660 4808
rect 19700 4768 22348 4808
rect 22388 4768 22397 4808
rect 22531 4768 22540 4808
rect 22580 4768 25996 4808
rect 26036 4768 26045 4808
rect 8755 4684 8764 4724
rect 8804 4684 10004 4724
rect 0 4640 90 4660
rect 0 4600 1228 4640
rect 1268 4600 1277 4640
rect 0 4580 90 4600
rect 4919 4516 4928 4556
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 5296 4516 5305 4556
rect 9964 4472 10004 4684
rect 13132 4556 13172 4768
rect 26092 4724 26132 4936
rect 31660 4892 31700 4936
rect 44908 4892 44948 4936
rect 46278 4916 46368 4936
rect 31660 4852 33676 4892
rect 33716 4852 33725 4892
rect 43171 4852 43180 4892
rect 43220 4852 44948 4892
rect 26323 4768 26332 4808
rect 26372 4768 32812 4808
rect 32852 4768 32861 4808
rect 33763 4768 33772 4808
rect 33812 4768 42124 4808
rect 42164 4768 42173 4808
rect 13315 4684 13324 4724
rect 13364 4684 19468 4724
rect 19508 4684 19517 4724
rect 20131 4684 20140 4724
rect 20180 4684 26132 4724
rect 31891 4684 31900 4724
rect 31940 4684 32428 4724
rect 32468 4684 32477 4724
rect 44755 4684 44764 4724
rect 44804 4684 45620 4724
rect 45580 4640 45620 4684
rect 46278 4640 46368 4660
rect 13891 4600 13900 4640
rect 13940 4600 16300 4640
rect 16340 4600 16349 4640
rect 19747 4600 19756 4640
rect 19796 4600 20564 4640
rect 23107 4600 23116 4640
rect 23156 4600 27148 4640
rect 27188 4600 27197 4640
rect 45580 4600 46368 4640
rect 20524 4556 20564 4600
rect 46278 4580 46368 4600
rect 13132 4516 16588 4556
rect 16628 4516 16637 4556
rect 20039 4516 20048 4556
rect 20088 4516 20130 4556
rect 20170 4516 20212 4556
rect 20252 4516 20294 4556
rect 20334 4516 20376 4556
rect 20416 4516 20425 4556
rect 20524 4516 24172 4556
rect 24212 4516 24221 4556
rect 25708 4516 31948 4556
rect 31988 4516 31997 4556
rect 35159 4516 35168 4556
rect 35208 4516 35250 4556
rect 35290 4516 35332 4556
rect 35372 4516 35414 4556
rect 35454 4516 35496 4556
rect 35536 4516 35545 4556
rect 25708 4472 25748 4516
rect 9964 4432 25748 4472
rect 25804 4432 27628 4472
rect 27668 4432 27677 4472
rect 25804 4388 25844 4432
rect 14179 4348 14188 4388
rect 14228 4348 19372 4388
rect 19412 4348 19421 4388
rect 19555 4348 19564 4388
rect 19604 4348 25844 4388
rect 0 4304 90 4324
rect 46278 4304 46368 4324
rect 0 4264 22924 4304
rect 22964 4264 22973 4304
rect 24019 4264 24028 4304
rect 24068 4264 25940 4304
rect 26035 4264 26044 4304
rect 26084 4264 31756 4304
rect 31796 4264 31805 4304
rect 34675 4264 34684 4304
rect 34724 4264 41740 4304
rect 41780 4264 41789 4304
rect 45139 4264 45148 4304
rect 45188 4264 46368 4304
rect 0 4244 90 4264
rect 25900 4220 25940 4264
rect 46278 4244 46368 4264
rect 17251 4180 17260 4220
rect 17300 4180 20812 4220
rect 20852 4180 20861 4220
rect 20995 4180 21004 4220
rect 21044 4180 22964 4220
rect 23011 4180 23020 4220
rect 23060 4180 24844 4220
rect 24884 4180 24893 4220
rect 25900 4180 33004 4220
rect 33044 4180 33053 4220
rect 33100 4180 38764 4220
rect 38804 4180 38813 4220
rect 22924 4136 22964 4180
rect 19267 4096 19276 4136
rect 19316 4096 22828 4136
rect 22868 4096 22877 4136
rect 22924 4096 23788 4136
rect 23828 4096 23837 4136
rect 25673 4096 25804 4136
rect 25844 4096 25853 4136
rect 26275 4096 26284 4136
rect 26324 4096 32332 4136
rect 32372 4096 32381 4136
rect 33100 4052 33140 4180
rect 34313 4096 34444 4136
rect 34484 4096 34493 4136
rect 40291 4096 40300 4136
rect 40340 4096 44524 4136
rect 44564 4096 44573 4136
rect 44620 4096 44908 4136
rect 44948 4096 44957 4136
rect 44620 4052 44660 4096
rect 14659 4012 14668 4052
rect 14708 4012 21676 4052
rect 21716 4012 21725 4052
rect 21859 4012 21868 4052
rect 21908 4012 33140 4052
rect 33187 4012 33196 4052
rect 33236 4012 44660 4052
rect 44755 4012 44764 4052
rect 44804 4012 45812 4052
rect 0 3968 90 3988
rect 45772 3968 45812 4012
rect 46278 3968 46368 3988
rect 0 3928 20140 3968
rect 20180 3928 20189 3968
rect 24067 3928 24076 3968
rect 24116 3928 38572 3968
rect 38612 3928 38621 3968
rect 45772 3928 46368 3968
rect 0 3908 90 3928
rect 46278 3908 46368 3928
rect 18499 3844 18508 3884
rect 18548 3844 21388 3884
rect 21428 3844 21437 3884
rect 25891 3844 25900 3884
rect 25940 3844 44564 3884
rect 3679 3760 3688 3800
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 4056 3760 4065 3800
rect 18799 3760 18808 3800
rect 18848 3760 18890 3800
rect 18930 3760 18972 3800
rect 19012 3760 19054 3800
rect 19094 3760 19136 3800
rect 19176 3760 19185 3800
rect 19843 3760 19852 3800
rect 19892 3760 22636 3800
rect 22676 3760 22685 3800
rect 28003 3760 28012 3800
rect 28052 3760 33140 3800
rect 33919 3760 33928 3800
rect 33968 3760 34010 3800
rect 34050 3760 34092 3800
rect 34132 3760 34174 3800
rect 34214 3760 34256 3800
rect 34296 3760 34305 3800
rect 33100 3716 33140 3760
rect 1411 3676 1420 3716
rect 1460 3676 31852 3716
rect 31892 3676 31901 3716
rect 32332 3676 32660 3716
rect 33100 3676 38860 3716
rect 38900 3676 38909 3716
rect 0 3632 90 3652
rect 32332 3632 32372 3676
rect 0 3592 25940 3632
rect 26995 3592 27004 3632
rect 27044 3592 31756 3632
rect 31796 3592 31805 3632
rect 32083 3592 32092 3632
rect 32132 3592 32372 3632
rect 32620 3632 32660 3676
rect 32620 3592 43276 3632
rect 43316 3592 43325 3632
rect 0 3572 90 3592
rect 1123 3508 1132 3548
rect 1172 3508 24116 3548
rect 24163 3508 24172 3548
rect 24212 3508 25804 3548
rect 25844 3508 25853 3548
rect 24076 3464 24116 3508
rect 25900 3464 25940 3592
rect 26131 3508 26140 3548
rect 26180 3508 27764 3548
rect 1315 3424 1324 3464
rect 1364 3424 17932 3464
rect 17972 3424 17981 3464
rect 18691 3424 18700 3464
rect 18740 3424 18988 3464
rect 19028 3424 19037 3464
rect 19180 3424 19756 3464
rect 19796 3424 19805 3464
rect 19939 3424 19948 3464
rect 19988 3424 21004 3464
rect 21044 3424 21053 3464
rect 21257 3424 21388 3464
rect 21428 3424 21437 3464
rect 21641 3424 21772 3464
rect 21812 3424 21821 3464
rect 22505 3424 22636 3464
rect 22676 3424 22685 3464
rect 22819 3424 22828 3464
rect 22868 3424 23020 3464
rect 23060 3424 23069 3464
rect 23395 3424 23404 3464
rect 23444 3424 23453 3464
rect 24067 3424 24076 3464
rect 24116 3424 24125 3464
rect 24451 3424 24460 3464
rect 24500 3424 24509 3464
rect 24713 3424 24844 3464
rect 24884 3424 24893 3464
rect 25891 3424 25900 3464
rect 25940 3424 25949 3464
rect 26633 3424 26764 3464
rect 26804 3424 26813 3464
rect 27619 3424 27628 3464
rect 27668 3424 27677 3464
rect 19180 3380 19220 3424
rect 23404 3380 23444 3424
rect 24460 3380 24500 3424
rect 27628 3380 27668 3424
rect 10051 3340 10060 3380
rect 10100 3340 19220 3380
rect 19276 3340 23444 3380
rect 23491 3340 23500 3380
rect 23540 3340 24500 3380
rect 24556 3340 27668 3380
rect 27724 3380 27764 3508
rect 44524 3464 44564 3844
rect 46278 3632 46368 3652
rect 45139 3592 45148 3632
rect 45188 3592 46368 3632
rect 46278 3572 46368 3592
rect 27859 3424 27868 3464
rect 27908 3424 30548 3464
rect 31721 3424 31852 3464
rect 31892 3424 31901 3464
rect 32419 3424 32428 3464
rect 32468 3424 43084 3464
rect 43124 3424 43133 3464
rect 44515 3424 44524 3464
rect 44564 3424 44573 3464
rect 44899 3424 44908 3464
rect 44948 3424 44957 3464
rect 30508 3380 30548 3424
rect 44908 3380 44948 3424
rect 27724 3340 29684 3380
rect 30508 3340 33100 3380
rect 33140 3340 33149 3380
rect 33292 3340 33388 3380
rect 33428 3340 33437 3380
rect 43180 3340 44948 3380
rect 0 3296 90 3316
rect 19276 3296 19316 3340
rect 24556 3296 24596 3340
rect 29644 3296 29684 3340
rect 33292 3296 33332 3340
rect 43180 3296 43220 3340
rect 46278 3296 46368 3316
rect 0 3256 2188 3296
rect 2228 3256 2237 3296
rect 8131 3256 8140 3296
rect 8180 3256 19316 3296
rect 19852 3256 22924 3296
rect 22964 3256 22973 3296
rect 23107 3256 23116 3296
rect 23156 3256 24596 3296
rect 25075 3256 25084 3296
rect 25124 3256 29108 3296
rect 29644 3256 33332 3296
rect 33475 3256 33484 3296
rect 33524 3256 43220 3296
rect 44755 3256 44764 3296
rect 44804 3256 46368 3296
rect 0 3236 90 3256
rect 19219 3172 19228 3212
rect 19268 3172 19564 3212
rect 19604 3172 19613 3212
rect 19852 3128 19892 3256
rect 29068 3212 29108 3256
rect 46278 3236 46368 3256
rect 19987 3172 19996 3212
rect 20036 3172 21140 3212
rect 21235 3172 21244 3212
rect 21284 3172 21484 3212
rect 21524 3172 21533 3212
rect 21619 3172 21628 3212
rect 21668 3172 21868 3212
rect 21908 3172 21917 3212
rect 22003 3172 22012 3212
rect 22052 3172 22772 3212
rect 22867 3172 22876 3212
rect 22916 3172 23060 3212
rect 23251 3172 23260 3212
rect 23300 3172 23404 3212
rect 23444 3172 23453 3212
rect 23635 3172 23644 3212
rect 23684 3172 24212 3212
rect 24307 3172 24316 3212
rect 24356 3172 24596 3212
rect 24691 3172 24700 3212
rect 24740 3172 28780 3212
rect 28820 3172 28829 3212
rect 29068 3172 33388 3212
rect 33428 3172 33437 3212
rect 34313 3172 34444 3212
rect 34484 3172 34723 3212
rect 34763 3172 34772 3212
rect 1411 3088 1420 3128
rect 1460 3088 17396 3128
rect 17923 3088 17932 3128
rect 17972 3088 19892 3128
rect 21100 3128 21140 3172
rect 21100 3088 21908 3128
rect 4919 3004 4928 3044
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 5296 3004 5305 3044
rect 0 2960 90 2980
rect 17356 2960 17396 3088
rect 18595 3004 18604 3044
rect 18644 3004 19948 3044
rect 19988 3004 19997 3044
rect 20039 3004 20048 3044
rect 20088 3004 20130 3044
rect 20170 3004 20212 3044
rect 20252 3004 20294 3044
rect 20334 3004 20376 3044
rect 20416 3004 20425 3044
rect 20524 3004 21772 3044
rect 21812 3004 21821 3044
rect 20524 2960 20564 3004
rect 0 2920 17260 2960
rect 17300 2920 17309 2960
rect 17356 2920 20564 2960
rect 21868 2960 21908 3088
rect 22732 3044 22772 3172
rect 23020 3128 23060 3172
rect 23020 3088 23348 3128
rect 22732 3004 23116 3044
rect 23156 3004 23165 3044
rect 23308 2960 23348 3088
rect 24172 3044 24212 3172
rect 24556 3128 24596 3172
rect 24556 3088 32428 3128
rect 32468 3088 32477 3128
rect 33196 3088 44620 3128
rect 44660 3088 44669 3128
rect 33196 3044 33236 3088
rect 24172 3004 33236 3044
rect 35159 3004 35168 3044
rect 35208 3004 35250 3044
rect 35290 3004 35332 3044
rect 35372 3004 35414 3044
rect 35454 3004 35496 3044
rect 35536 3004 35545 3044
rect 35884 3004 44140 3044
rect 44180 3004 44189 3044
rect 21868 2920 23020 2960
rect 23060 2920 23069 2960
rect 23308 2920 28012 2960
rect 28052 2920 28061 2960
rect 28771 2920 28780 2960
rect 28820 2920 35732 2960
rect 0 2900 90 2920
rect 35692 2876 35732 2920
rect 35884 2876 35924 3004
rect 46278 2960 46368 2980
rect 40291 2920 40300 2960
rect 40340 2920 44948 2960
rect 18259 2836 18268 2876
rect 18308 2836 28876 2876
rect 28916 2836 28925 2876
rect 35692 2836 35924 2876
rect 1219 2752 1228 2792
rect 1268 2752 27188 2792
rect 7180 2668 19948 2708
rect 19988 2668 19997 2708
rect 0 2624 90 2644
rect 7180 2624 7220 2668
rect 27148 2624 27188 2752
rect 38851 2668 38860 2708
rect 38900 2668 44564 2708
rect 44524 2624 44564 2668
rect 44908 2624 44948 2920
rect 45484 2920 46368 2960
rect 45484 2876 45524 2920
rect 46278 2900 46368 2920
rect 45139 2836 45148 2876
rect 45188 2836 45524 2876
rect 46278 2624 46368 2644
rect 0 2584 7220 2624
rect 10435 2584 10444 2624
rect 10484 2584 11308 2624
rect 11348 2584 11357 2624
rect 12547 2584 12556 2624
rect 12596 2584 18028 2624
rect 18068 2584 18077 2624
rect 27139 2584 27148 2624
rect 27188 2584 27197 2624
rect 27244 2584 28012 2624
rect 28052 2584 28061 2624
rect 44009 2584 44140 2624
rect 44180 2584 44189 2624
rect 44515 2584 44524 2624
rect 44564 2584 44573 2624
rect 44899 2584 44908 2624
rect 44948 2584 44957 2624
rect 45772 2584 46368 2624
rect 0 2564 90 2584
rect 27244 2540 27284 2584
rect 45772 2540 45812 2584
rect 46278 2564 46368 2584
rect 7180 2500 27284 2540
rect 27379 2500 27388 2540
rect 27428 2500 40876 2540
rect 40916 2500 40925 2540
rect 44755 2500 44764 2540
rect 44804 2500 45812 2540
rect 7180 2372 7220 2500
rect 11539 2416 11548 2456
rect 11588 2416 17300 2456
rect 28243 2416 28252 2456
rect 28292 2416 40780 2456
rect 40820 2416 40829 2456
rect 44371 2416 44380 2456
rect 44420 2416 45044 2456
rect 643 2332 652 2372
rect 692 2332 7220 2372
rect 0 2288 90 2308
rect 0 2248 3572 2288
rect 3679 2248 3688 2288
rect 3728 2248 3770 2288
rect 3810 2248 3852 2288
rect 3892 2248 3934 2288
rect 3974 2248 4016 2288
rect 4056 2248 4065 2288
rect 0 2228 90 2248
rect 3532 2204 3572 2248
rect 3532 2164 8140 2204
rect 8180 2164 8189 2204
rect 17260 2120 17300 2416
rect 18799 2248 18808 2288
rect 18848 2248 18890 2288
rect 18930 2248 18972 2288
rect 19012 2248 19054 2288
rect 19094 2248 19136 2288
rect 19176 2248 19185 2288
rect 33919 2248 33928 2288
rect 33968 2248 34010 2288
rect 34050 2248 34092 2288
rect 34132 2248 34174 2288
rect 34214 2248 34256 2288
rect 34296 2248 34305 2288
rect 19555 2164 19564 2204
rect 19604 2164 44564 2204
rect 17260 2080 32236 2120
rect 32276 2080 32285 2120
rect 21475 1996 21484 2036
rect 21524 1996 44180 2036
rect 0 1952 90 1972
rect 44140 1952 44180 1996
rect 44524 1952 44564 2164
rect 44611 1996 44620 2036
rect 44660 1996 44669 2036
rect 44620 1952 44660 1996
rect 45004 1952 45044 2416
rect 46278 2288 46368 2308
rect 45772 2248 46368 2288
rect 45772 2120 45812 2248
rect 46278 2228 46368 2248
rect 45139 2080 45148 2120
rect 45188 2080 45812 2120
rect 46278 1952 46368 1972
rect 0 1912 1324 1952
rect 1364 1912 1373 1952
rect 38563 1912 38572 1952
rect 38612 1912 43372 1952
rect 43412 1912 43421 1952
rect 43747 1912 43756 1952
rect 43796 1912 43805 1952
rect 44131 1912 44140 1952
rect 44180 1912 44189 1952
rect 44515 1912 44524 1952
rect 44564 1912 44573 1952
rect 44620 1912 44908 1952
rect 44948 1912 44957 1952
rect 45004 1912 46368 1952
rect 0 1892 90 1912
rect 43756 1868 43796 1912
rect 46278 1892 46368 1912
rect 38755 1828 38764 1868
rect 38804 1828 43796 1868
rect 43987 1744 43996 1784
rect 44036 1744 45676 1784
rect 45716 1744 45725 1784
rect 43603 1660 43612 1700
rect 43652 1660 44276 1700
rect 44371 1660 44380 1700
rect 44420 1660 44620 1700
rect 44660 1660 44669 1700
rect 44755 1660 44764 1700
rect 44804 1660 45044 1700
rect 0 1616 90 1636
rect 0 1576 18700 1616
rect 18740 1576 18749 1616
rect 0 1556 90 1576
rect 44236 1532 44276 1660
rect 45004 1616 45044 1660
rect 46278 1616 46368 1636
rect 45004 1576 46368 1616
rect 46278 1556 46368 1576
rect 4919 1492 4928 1532
rect 4968 1492 5010 1532
rect 5050 1492 5092 1532
rect 5132 1492 5174 1532
rect 5214 1492 5256 1532
rect 5296 1492 5305 1532
rect 20039 1492 20048 1532
rect 20088 1492 20130 1532
rect 20170 1492 20212 1532
rect 20252 1492 20294 1532
rect 20334 1492 20376 1532
rect 20416 1492 20425 1532
rect 35159 1492 35168 1532
rect 35208 1492 35250 1532
rect 35290 1492 35332 1532
rect 35372 1492 35414 1532
rect 35454 1492 35496 1532
rect 35536 1492 35545 1532
rect 44236 1492 45044 1532
rect 0 1280 90 1300
rect 45004 1280 45044 1492
rect 46278 1280 46368 1300
rect 0 1240 1420 1280
rect 1460 1240 1469 1280
rect 45004 1240 46368 1280
rect 0 1220 90 1240
rect 46278 1220 46368 1240
rect 0 944 90 964
rect 46278 944 46368 964
rect 0 904 18508 944
rect 18548 904 18557 944
rect 45667 904 45676 944
rect 45716 904 46368 944
rect 0 884 90 904
rect 46278 884 46368 904
rect 0 608 90 628
rect 46278 608 46368 628
rect 0 568 18604 608
rect 18644 568 18653 608
rect 44611 568 44620 608
rect 44660 568 46368 608
rect 0 548 90 568
rect 46278 548 46368 568
<< via2 >>
rect 9580 11740 9620 11780
rect 22156 11740 22196 11780
rect 9868 11656 9908 11696
rect 22348 11656 22388 11696
rect 16492 11572 16532 11612
rect 24460 11572 24500 11612
rect 10060 11488 10100 11528
rect 21964 11488 22004 11528
rect 16300 11320 16340 11360
rect 23308 11320 23348 11360
rect 1324 10984 1364 11024
rect 15340 10984 15380 11024
rect 21772 10984 21812 11024
rect 44140 10984 44180 11024
rect 268 10648 308 10688
rect 19948 10648 19988 10688
rect 23884 10648 23924 10688
rect 43372 10648 43412 10688
rect 556 10312 596 10352
rect 43660 10312 43700 10352
rect 19564 10228 19604 10268
rect 23692 10228 23732 10268
rect 18028 10060 18068 10100
rect 20716 10060 20756 10100
rect 32620 10060 32660 10100
rect 36076 10060 36116 10100
rect 1420 9976 1460 10016
rect 20524 9976 20564 10016
rect 32428 9976 32468 10016
rect 34828 9976 34868 10016
rect 44428 9976 44468 10016
rect 17644 9892 17684 9932
rect 27052 9892 27092 9932
rect 30508 9892 30548 9932
rect 35692 9892 35732 9932
rect 3688 9808 3728 9848
rect 3770 9808 3810 9848
rect 3852 9808 3892 9848
rect 3934 9808 3974 9848
rect 4016 9808 4056 9848
rect 18808 9808 18848 9848
rect 18890 9808 18930 9848
rect 18972 9808 19012 9848
rect 19054 9808 19094 9848
rect 19136 9808 19176 9848
rect 18604 9724 18644 9764
rect 27532 9808 27572 9848
rect 32332 9808 32372 9848
rect 33004 9808 33044 9848
rect 33928 9808 33968 9848
rect 34010 9808 34050 9848
rect 34092 9808 34132 9848
rect 34174 9808 34214 9848
rect 34256 9808 34296 9848
rect 1420 9640 1460 9680
rect 11212 9640 11252 9680
rect 11596 9640 11636 9680
rect 11980 9640 12020 9680
rect 12364 9640 12404 9680
rect 12748 9640 12788 9680
rect 13132 9640 13172 9680
rect 13516 9640 13556 9680
rect 13900 9640 13940 9680
rect 14284 9640 14324 9680
rect 14668 9640 14708 9680
rect 15052 9640 15092 9680
rect 15436 9640 15476 9680
rect 15820 9640 15860 9680
rect 16204 9640 16244 9680
rect 16588 9640 16628 9680
rect 16972 9640 17012 9680
rect 17356 9640 17396 9680
rect 17740 9640 17780 9680
rect 18124 9640 18164 9680
rect 18508 9640 18548 9680
rect 18796 9640 18836 9680
rect 10348 9556 10388 9596
rect 19372 9640 19412 9680
rect 19660 9556 19700 9596
rect 20812 9724 20852 9764
rect 31948 9724 31988 9764
rect 20236 9640 20276 9680
rect 20620 9640 20660 9680
rect 31180 9640 31220 9680
rect 31564 9640 31604 9680
rect 33676 9640 33716 9680
rect 20428 9556 20468 9596
rect 28780 9556 28820 9596
rect 31372 9556 31412 9596
rect 31756 9556 31796 9596
rect 32716 9556 32756 9596
rect 43372 9640 43412 9680
rect 43660 9640 43700 9680
rect 35020 9556 35060 9596
rect 36748 9556 36788 9596
rect 9484 9472 9524 9512
rect 11308 9472 11348 9512
rect 13228 9472 13268 9512
rect 13804 9472 13844 9512
rect 14188 9472 14228 9512
rect 15052 9472 15092 9512
rect 15436 9472 15476 9512
rect 15724 9472 15764 9512
rect 16972 9472 17012 9512
rect 17452 9472 17492 9512
rect 17644 9472 17684 9512
rect 18028 9472 18068 9512
rect 18796 9472 18836 9512
rect 27340 9472 27380 9512
rect 31468 9472 31508 9512
rect 31660 9472 31700 9512
rect 32044 9472 32084 9512
rect 32812 9472 32852 9512
rect 33964 9472 34004 9512
rect 34732 9472 34772 9512
rect 35692 9472 35732 9512
rect 36076 9472 36116 9512
rect 36460 9472 36500 9512
rect 37708 9472 37748 9512
rect 42988 9472 43028 9512
rect 43372 9472 43412 9512
rect 43756 9472 43796 9512
rect 8620 9388 8660 9428
rect 11212 9388 11252 9428
rect 14284 9388 14324 9428
rect 1420 9304 1460 9344
rect 10156 9304 10196 9344
rect 17260 9388 17300 9428
rect 19756 9388 19796 9428
rect 20044 9388 20084 9428
rect 18028 9304 18068 9344
rect 28012 9388 28052 9428
rect 32236 9388 32276 9428
rect 33100 9388 33140 9428
rect 27916 9304 27956 9344
rect 30892 9304 30932 9344
rect 21004 9220 21044 9260
rect 32332 9220 32372 9260
rect 33004 9220 33044 9260
rect 4928 9052 4968 9092
rect 5010 9052 5050 9092
rect 5092 9052 5132 9092
rect 5174 9052 5214 9092
rect 5256 9052 5296 9092
rect 1420 8968 1460 9008
rect 9772 8968 9812 9008
rect 11020 8884 11060 8924
rect 11404 8884 11444 8924
rect 11788 8884 11828 8924
rect 12172 8884 12212 8924
rect 12556 8884 12596 8924
rect 10540 8800 10580 8840
rect 8716 8716 8756 8756
rect 11500 8716 11540 8756
rect 13324 8884 13364 8924
rect 13708 8884 13748 8924
rect 14092 8884 14132 8924
rect 14476 8884 14516 8924
rect 14860 8884 14900 8924
rect 15244 8884 15284 8924
rect 15628 8884 15668 8924
rect 16012 8884 16052 8924
rect 16396 8884 16436 8924
rect 16780 8884 16820 8924
rect 17164 8884 17204 8924
rect 17548 8884 17588 8924
rect 17932 8884 17972 8924
rect 13516 8716 13556 8756
rect 17164 8716 17204 8756
rect 18124 8716 18164 8756
rect 19756 9136 19796 9176
rect 20620 9136 20660 9176
rect 33484 9388 33524 9428
rect 35596 9388 35636 9428
rect 36940 9388 36980 9428
rect 43948 9388 43988 9428
rect 33580 9304 33620 9344
rect 34444 9304 34484 9344
rect 35980 9304 36020 9344
rect 20812 9136 20852 9176
rect 26668 9136 26708 9176
rect 27244 9136 27284 9176
rect 30604 9136 30644 9176
rect 31756 9136 31796 9176
rect 35788 9220 35828 9260
rect 37996 9220 38036 9260
rect 40204 9220 40244 9260
rect 45772 9220 45812 9260
rect 33772 9136 33812 9176
rect 34540 9136 34580 9176
rect 36364 9136 36404 9176
rect 37804 9136 37844 9176
rect 18892 9052 18932 9092
rect 19948 9052 19988 9092
rect 20048 9052 20088 9092
rect 20130 9052 20170 9092
rect 20212 9052 20252 9092
rect 20294 9052 20334 9092
rect 20376 9052 20416 9092
rect 21676 9052 21716 9092
rect 25132 9052 25172 9092
rect 30796 9052 30836 9092
rect 31948 9052 31988 9092
rect 32812 9052 32852 9092
rect 33196 9052 33236 9092
rect 34444 9052 34484 9092
rect 35020 9052 35060 9092
rect 35168 9052 35208 9092
rect 35250 9052 35290 9092
rect 35332 9052 35372 9092
rect 35414 9052 35454 9092
rect 35496 9052 35536 9092
rect 37900 9052 37940 9092
rect 40108 9052 40148 9092
rect 18316 8884 18356 8924
rect 18700 8884 18740 8924
rect 19276 8884 19316 8924
rect 19468 8884 19508 8924
rect 19852 8884 19892 8924
rect 21676 8884 21716 8924
rect 25036 8884 25076 8924
rect 26380 8800 26420 8840
rect 24268 8716 24308 8756
rect 27244 8716 27284 8756
rect 30988 8968 31028 9008
rect 39916 8968 39956 9008
rect 27532 8884 27572 8924
rect 28876 8884 28916 8924
rect 32140 8884 32180 8924
rect 32524 8884 32564 8924
rect 32908 8884 32948 8924
rect 33292 8884 33332 8924
rect 34252 8884 34283 8924
rect 34283 8884 34292 8924
rect 35020 8884 35060 8924
rect 36460 8884 36500 8924
rect 36748 8884 36788 8924
rect 37228 8884 37259 8924
rect 37259 8884 37268 8924
rect 37804 8884 37844 8924
rect 39820 8884 39860 8924
rect 40300 8884 40340 8924
rect 43756 8884 43796 8924
rect 44140 8884 44180 8924
rect 44428 8884 44468 8924
rect 27916 8800 27956 8840
rect 28300 8800 28340 8840
rect 33196 8800 33236 8840
rect 33964 8800 34004 8840
rect 34348 8800 34388 8840
rect 34636 8800 34676 8840
rect 43372 8800 43412 8840
rect 28684 8716 28724 8756
rect 29164 8716 29204 8756
rect 33388 8716 33428 8756
rect 35980 8716 36020 8756
rect 36940 8716 36980 8756
rect 37420 8716 37460 8756
rect 1420 8632 1460 8672
rect 9100 8632 9140 8672
rect 12460 8632 12500 8672
rect 13612 8632 13652 8672
rect 13996 8632 14036 8672
rect 14380 8632 14420 8672
rect 15148 8632 15188 8672
rect 15532 8632 15572 8672
rect 15916 8632 15956 8672
rect 16684 8632 16724 8672
rect 17068 8632 17108 8672
rect 19756 8632 19796 8672
rect 25900 8632 25940 8672
rect 28012 8632 28052 8672
rect 28492 8632 28532 8672
rect 28780 8632 28820 8672
rect 30028 8632 30068 8672
rect 31852 8632 31892 8672
rect 32812 8632 32852 8672
rect 33004 8632 33044 8672
rect 33868 8632 33908 8672
rect 34348 8632 34388 8672
rect 34732 8632 34772 8672
rect 13036 8548 13076 8588
rect 20524 8548 20564 8588
rect 21676 8548 21716 8588
rect 35788 8632 35828 8672
rect 36076 8632 36116 8672
rect 36364 8632 36404 8672
rect 37900 8632 37940 8672
rect 38668 8632 38708 8672
rect 40204 8632 40244 8672
rect 40492 8632 40532 8672
rect 43948 8632 43988 8672
rect 45772 8632 45812 8672
rect 16780 8464 16820 8504
rect 22540 8464 22580 8504
rect 29836 8464 29876 8504
rect 45772 8464 45812 8504
rect 2956 8380 2996 8420
rect 26188 8380 26228 8420
rect 26572 8380 26612 8420
rect 30412 8380 30452 8420
rect 172 8296 212 8336
rect 3688 8296 3728 8336
rect 3770 8296 3810 8336
rect 3852 8296 3892 8336
rect 3934 8296 3974 8336
rect 4016 8296 4056 8336
rect 1324 8212 1364 8252
rect 2860 8128 2900 8168
rect 18808 8296 18848 8336
rect 18890 8296 18930 8336
rect 18972 8296 19012 8336
rect 19054 8296 19094 8336
rect 19136 8296 19176 8336
rect 26956 8296 26996 8336
rect 29452 8296 29492 8336
rect 33928 8296 33968 8336
rect 34010 8296 34050 8336
rect 34092 8296 34132 8336
rect 34174 8296 34214 8336
rect 34256 8296 34296 8336
rect 16588 8212 16628 8252
rect 22732 8212 22772 8252
rect 31852 8212 31892 8252
rect 24268 8128 24308 8168
rect 25900 8128 25940 8168
rect 26668 8128 26708 8168
rect 27052 8128 27092 8168
rect 40492 8128 40532 8168
rect 42988 8128 43028 8168
rect 20140 8044 20180 8084
rect 20908 8044 20948 8084
rect 27532 8044 27572 8084
rect 13708 7960 13748 8000
rect 24844 7960 24884 8000
rect 25132 7960 25172 8000
rect 25420 7960 25460 8000
rect 25900 7960 25940 8000
rect 26188 7960 26228 8000
rect 26572 7960 26612 8000
rect 26956 7960 26996 8000
rect 27244 7960 27284 8000
rect 28108 7960 28148 8000
rect 32716 7960 32756 8000
rect 34348 7960 34388 8000
rect 36172 7960 36212 8000
rect 36460 7960 36500 8000
rect 37420 7960 37460 8000
rect 37900 7960 37940 8000
rect 38668 7960 38708 8000
rect 43564 7960 43604 8000
rect 45772 7960 45812 8000
rect 268 7876 308 7916
rect 25036 7876 25076 7916
rect 29068 7876 29108 7916
rect 36940 7876 36980 7916
rect 35212 7792 35252 7832
rect 40300 7792 40340 7832
rect 27340 7708 27380 7748
rect 45772 7708 45812 7748
rect 4780 7624 4820 7664
rect 5548 7624 5588 7664
rect 35692 7624 35732 7664
rect 4928 7540 4968 7580
rect 5010 7540 5050 7580
rect 5092 7540 5132 7580
rect 5174 7540 5214 7580
rect 5256 7540 5296 7580
rect 20048 7540 20088 7580
rect 20130 7540 20170 7580
rect 20212 7540 20252 7580
rect 20294 7540 20334 7580
rect 20376 7540 20416 7580
rect 25900 7540 25940 7580
rect 30220 7540 30260 7580
rect 35168 7540 35208 7580
rect 35250 7540 35290 7580
rect 35332 7540 35372 7580
rect 35414 7540 35454 7580
rect 35496 7540 35536 7580
rect 172 7456 212 7496
rect 36460 7456 36500 7496
rect 25420 7372 25460 7412
rect 29932 7372 29972 7412
rect 36076 7372 36116 7412
rect 32716 7288 32756 7328
rect 45772 7288 45812 7328
rect 21196 7120 21236 7160
rect 29644 7120 29684 7160
rect 33292 7120 33332 7160
rect 35692 7120 35732 7160
rect 43564 7120 43604 7160
rect 44524 7120 44564 7160
rect 8620 7036 8660 7076
rect 32044 7036 32084 7076
rect 7852 6952 7892 6992
rect 8044 6952 8084 6992
rect 18700 6952 18740 6992
rect 15820 6868 15860 6908
rect 24076 6868 24116 6908
rect 3688 6784 3728 6824
rect 3770 6784 3810 6824
rect 3852 6784 3892 6824
rect 3934 6784 3974 6824
rect 4016 6784 4056 6824
rect 8812 6784 8852 6824
rect 15340 6784 15380 6824
rect 18808 6784 18848 6824
rect 18890 6784 18930 6824
rect 18972 6784 19012 6824
rect 19054 6784 19094 6824
rect 19136 6784 19176 6824
rect 19852 6784 19892 6824
rect 21388 6784 21428 6824
rect 33928 6784 33968 6824
rect 34010 6784 34050 6824
rect 34092 6784 34132 6824
rect 34174 6784 34214 6824
rect 34256 6784 34296 6824
rect 16876 6700 16916 6740
rect 21580 6700 21620 6740
rect 8044 6616 8084 6656
rect 8716 6532 8756 6572
rect 9100 6532 9140 6572
rect 9484 6532 9524 6572
rect 14188 6532 14228 6572
rect 15532 6532 15572 6572
rect 23500 6532 23540 6572
rect 6220 6448 6260 6488
rect 8428 6448 8468 6488
rect 8812 6448 8852 6488
rect 19372 6448 19412 6488
rect 26476 6448 26516 6488
rect 35692 6448 35732 6488
rect 41740 6448 41780 6488
rect 44908 6448 44948 6488
rect 4108 6364 4148 6404
rect 16876 6364 16916 6404
rect 17068 6364 17108 6404
rect 25996 6364 26036 6404
rect 748 6280 788 6320
rect 31660 6280 31700 6320
rect 15724 6196 15764 6236
rect 19372 6112 19412 6152
rect 21964 6112 22004 6152
rect 44524 6112 44564 6152
rect 46252 6112 46292 6152
rect 4928 6028 4968 6068
rect 5010 6028 5050 6068
rect 5092 6028 5132 6068
rect 5174 6028 5214 6068
rect 5256 6028 5296 6068
rect 8428 6028 8468 6068
rect 19852 6028 19892 6068
rect 20048 6028 20088 6068
rect 20130 6028 20170 6068
rect 20212 6028 20252 6068
rect 20294 6028 20334 6068
rect 20376 6028 20416 6068
rect 24844 6028 24884 6068
rect 27436 6028 27476 6068
rect 35168 6028 35208 6068
rect 35250 6028 35290 6068
rect 35332 6028 35372 6068
rect 35414 6028 35454 6068
rect 35496 6028 35536 6068
rect 34444 5944 34484 5984
rect 46252 5944 46292 5984
rect 7852 5860 7892 5900
rect 33292 5860 33332 5900
rect 15820 5776 15860 5816
rect 18028 5776 18068 5816
rect 18604 5776 18644 5816
rect 21964 5776 22004 5816
rect 24844 5776 24884 5816
rect 25036 5776 25076 5816
rect 14284 5692 14324 5732
rect 15148 5692 15188 5732
rect 17260 5692 17300 5732
rect 20044 5692 20084 5732
rect 20524 5692 20564 5732
rect 23020 5692 23060 5732
rect 25228 5692 25268 5732
rect 26860 5692 26900 5732
rect 27340 5692 27380 5732
rect 29548 5692 29588 5732
rect 1420 5608 1460 5648
rect 1996 5608 2036 5648
rect 9580 5608 9620 5648
rect 9868 5608 9908 5648
rect 10252 5608 10292 5648
rect 10636 5608 10676 5648
rect 11020 5608 11060 5648
rect 11308 5608 11348 5648
rect 11596 5608 11636 5648
rect 11884 5608 11924 5648
rect 13324 5608 13364 5648
rect 13612 5608 13652 5648
rect 14380 5608 14420 5648
rect 14668 5608 14708 5648
rect 14956 5608 14996 5648
rect 15340 5608 15380 5648
rect 18124 5608 18164 5648
rect 18508 5608 18548 5648
rect 19276 5608 19316 5648
rect 19660 5608 19700 5648
rect 9772 5524 9812 5564
rect 10156 5524 10196 5564
rect 10540 5524 10580 5564
rect 11500 5524 11540 5564
rect 12460 5524 12500 5564
rect 13516 5524 13556 5564
rect 13708 5524 13748 5564
rect 13996 5524 14036 5564
rect 19852 5524 19892 5564
rect 11212 5440 11252 5480
rect 13228 5440 13268 5480
rect 14860 5440 14900 5480
rect 16492 5440 16532 5480
rect 21196 5608 21236 5648
rect 23212 5608 23252 5648
rect 29836 5608 29876 5648
rect 30028 5608 30068 5648
rect 31564 5608 31604 5648
rect 32044 5608 32084 5648
rect 33388 5608 33428 5648
rect 33772 5608 33812 5648
rect 34348 5608 34388 5648
rect 21772 5524 21812 5564
rect 31468 5524 31508 5564
rect 20428 5440 20468 5480
rect 20716 5440 20756 5480
rect 21292 5440 21332 5480
rect 23020 5440 23060 5480
rect 23308 5440 23348 5480
rect 25324 5440 25364 5480
rect 29932 5440 29972 5480
rect 30508 5440 30548 5480
rect 30892 5440 30932 5480
rect 32620 5440 32660 5480
rect 18508 5356 18548 5396
rect 652 5272 692 5312
rect 3688 5272 3728 5312
rect 3770 5272 3810 5312
rect 3852 5272 3892 5312
rect 3934 5272 3974 5312
rect 4016 5272 4056 5312
rect 10252 5272 10292 5312
rect 18808 5272 18848 5312
rect 18890 5272 18930 5312
rect 18972 5272 19012 5312
rect 19054 5272 19094 5312
rect 19136 5272 19176 5312
rect 20044 5356 20084 5396
rect 25036 5356 25076 5396
rect 26764 5356 26804 5396
rect 33100 5356 33140 5396
rect 24940 5272 24980 5312
rect 25228 5272 25268 5312
rect 29836 5272 29876 5312
rect 44236 5692 44276 5732
rect 35596 5608 35636 5648
rect 40780 5608 40820 5648
rect 43276 5524 43316 5564
rect 40012 5440 40052 5480
rect 46252 5440 46292 5480
rect 37900 5356 37940 5396
rect 33928 5272 33968 5312
rect 34010 5272 34050 5312
rect 34092 5272 34132 5312
rect 34174 5272 34214 5312
rect 34256 5272 34296 5312
rect 46252 5272 46292 5312
rect 21196 5188 21236 5228
rect 26284 5188 26324 5228
rect 44908 5188 44948 5228
rect 10348 5104 10388 5144
rect 13804 5104 13844 5144
rect 16780 5104 16820 5144
rect 17452 5104 17492 5144
rect 22348 5104 22388 5144
rect 25612 5104 25652 5144
rect 11596 5020 11636 5060
rect 16108 5020 16148 5060
rect 16684 5020 16724 5060
rect 19948 5020 19988 5060
rect 21676 5020 21716 5060
rect 32044 5104 32084 5144
rect 34732 5104 34772 5144
rect 1132 4936 1172 4976
rect 8332 4936 8372 4976
rect 10060 4936 10100 4976
rect 11020 4936 11060 4976
rect 13900 4936 13940 4976
rect 14188 4936 14228 4976
rect 15916 4936 15956 4976
rect 19180 4936 19220 4976
rect 19564 4936 19604 4976
rect 21484 4936 21524 4976
rect 25708 4936 25748 4976
rect 29932 5020 29972 5060
rect 34828 5020 34868 5060
rect 35788 4936 35828 4976
rect 40876 4936 40916 4976
rect 748 4852 788 4892
rect 10636 4768 10676 4808
rect 15052 4768 15092 4808
rect 19660 4768 19700 4808
rect 22348 4768 22388 4808
rect 22540 4768 22580 4808
rect 25996 4768 26036 4808
rect 1228 4600 1268 4640
rect 4928 4516 4968 4556
rect 5010 4516 5050 4556
rect 5092 4516 5132 4556
rect 5174 4516 5214 4556
rect 5256 4516 5296 4556
rect 33676 4852 33716 4892
rect 43180 4852 43220 4892
rect 32812 4768 32852 4808
rect 33772 4768 33812 4808
rect 42124 4768 42164 4808
rect 13324 4684 13364 4724
rect 19468 4684 19508 4724
rect 20140 4684 20180 4724
rect 32428 4684 32468 4724
rect 13900 4600 13940 4640
rect 16300 4600 16340 4640
rect 19756 4600 19796 4640
rect 23116 4600 23156 4640
rect 27148 4600 27188 4640
rect 16588 4516 16628 4556
rect 20048 4516 20088 4556
rect 20130 4516 20170 4556
rect 20212 4516 20252 4556
rect 20294 4516 20334 4556
rect 20376 4516 20416 4556
rect 24172 4516 24212 4556
rect 31948 4516 31988 4556
rect 35168 4516 35208 4556
rect 35250 4516 35290 4556
rect 35332 4516 35372 4556
rect 35414 4516 35454 4556
rect 35496 4516 35536 4556
rect 27628 4432 27668 4472
rect 14188 4348 14228 4388
rect 19372 4348 19412 4388
rect 19564 4348 19604 4388
rect 22924 4264 22964 4304
rect 31756 4264 31796 4304
rect 41740 4264 41780 4304
rect 17260 4180 17300 4220
rect 20812 4180 20852 4220
rect 21004 4180 21044 4220
rect 23020 4180 23060 4220
rect 24844 4180 24884 4220
rect 33004 4180 33044 4220
rect 38764 4180 38804 4220
rect 19276 4096 19316 4136
rect 22828 4096 22868 4136
rect 25804 4096 25844 4136
rect 26284 4096 26324 4136
rect 32332 4096 32372 4136
rect 34444 4096 34484 4136
rect 40300 4096 40340 4136
rect 14668 4012 14708 4052
rect 21676 4012 21716 4052
rect 21868 4012 21908 4052
rect 33196 4012 33236 4052
rect 20140 3928 20180 3968
rect 24076 3928 24116 3968
rect 38572 3928 38612 3968
rect 18508 3844 18548 3884
rect 21388 3844 21428 3884
rect 25900 3844 25940 3884
rect 3688 3760 3728 3800
rect 3770 3760 3810 3800
rect 3852 3760 3892 3800
rect 3934 3760 3974 3800
rect 4016 3760 4056 3800
rect 18808 3760 18848 3800
rect 18890 3760 18930 3800
rect 18972 3760 19012 3800
rect 19054 3760 19094 3800
rect 19136 3760 19176 3800
rect 19852 3760 19892 3800
rect 22636 3760 22676 3800
rect 28012 3760 28052 3800
rect 33928 3760 33968 3800
rect 34010 3760 34050 3800
rect 34092 3760 34132 3800
rect 34174 3760 34214 3800
rect 34256 3760 34296 3800
rect 1420 3676 1460 3716
rect 31852 3676 31892 3716
rect 38860 3676 38900 3716
rect 31756 3592 31796 3632
rect 43276 3592 43316 3632
rect 1132 3508 1172 3548
rect 24172 3508 24212 3548
rect 25804 3508 25844 3548
rect 1324 3424 1364 3464
rect 17932 3424 17972 3464
rect 18700 3424 18740 3464
rect 19948 3424 19988 3464
rect 21388 3424 21428 3464
rect 21772 3424 21812 3464
rect 22636 3424 22676 3464
rect 22828 3424 22868 3464
rect 24844 3424 24884 3464
rect 26764 3424 26804 3464
rect 10060 3340 10100 3380
rect 23500 3340 23540 3380
rect 31852 3424 31892 3464
rect 32428 3424 32468 3464
rect 43084 3424 43124 3464
rect 33100 3340 33140 3380
rect 33388 3340 33428 3380
rect 2188 3256 2228 3296
rect 8140 3256 8180 3296
rect 22924 3256 22964 3296
rect 23116 3256 23156 3296
rect 33484 3256 33524 3296
rect 19564 3172 19604 3212
rect 21484 3172 21524 3212
rect 21868 3172 21908 3212
rect 23404 3172 23444 3212
rect 28780 3172 28820 3212
rect 33388 3172 33428 3212
rect 34444 3172 34484 3212
rect 1420 3088 1460 3128
rect 17932 3088 17972 3128
rect 4928 3004 4968 3044
rect 5010 3004 5050 3044
rect 5092 3004 5132 3044
rect 5174 3004 5214 3044
rect 5256 3004 5296 3044
rect 18604 3004 18644 3044
rect 19948 3004 19988 3044
rect 20048 3004 20088 3044
rect 20130 3004 20170 3044
rect 20212 3004 20252 3044
rect 20294 3004 20334 3044
rect 20376 3004 20416 3044
rect 21772 3004 21812 3044
rect 17260 2920 17300 2960
rect 23116 3004 23156 3044
rect 32428 3088 32468 3128
rect 44620 3088 44660 3128
rect 35168 3004 35208 3044
rect 35250 3004 35290 3044
rect 35332 3004 35372 3044
rect 35414 3004 35454 3044
rect 35496 3004 35536 3044
rect 44140 3004 44180 3044
rect 23020 2920 23060 2960
rect 28012 2920 28052 2960
rect 28780 2920 28820 2960
rect 40300 2920 40340 2960
rect 28876 2836 28916 2876
rect 1228 2752 1268 2792
rect 19948 2668 19988 2708
rect 38860 2668 38900 2708
rect 10444 2584 10484 2624
rect 12556 2584 12596 2624
rect 44140 2584 44180 2624
rect 40876 2500 40916 2540
rect 40780 2416 40820 2456
rect 652 2332 692 2372
rect 3688 2248 3728 2288
rect 3770 2248 3810 2288
rect 3852 2248 3892 2288
rect 3934 2248 3974 2288
rect 4016 2248 4056 2288
rect 8140 2164 8180 2204
rect 18808 2248 18848 2288
rect 18890 2248 18930 2288
rect 18972 2248 19012 2288
rect 19054 2248 19094 2288
rect 19136 2248 19176 2288
rect 33928 2248 33968 2288
rect 34010 2248 34050 2288
rect 34092 2248 34132 2288
rect 34174 2248 34214 2288
rect 34256 2248 34296 2288
rect 19564 2164 19604 2204
rect 32236 2080 32276 2120
rect 21484 1996 21524 2036
rect 44620 1996 44660 2036
rect 1324 1912 1364 1952
rect 38572 1912 38612 1952
rect 38764 1828 38804 1868
rect 45676 1744 45716 1784
rect 44620 1660 44660 1700
rect 18700 1576 18740 1616
rect 4928 1492 4968 1532
rect 5010 1492 5050 1532
rect 5092 1492 5132 1532
rect 5174 1492 5214 1532
rect 5256 1492 5296 1532
rect 20048 1492 20088 1532
rect 20130 1492 20170 1532
rect 20212 1492 20252 1532
rect 20294 1492 20334 1532
rect 20376 1492 20416 1532
rect 35168 1492 35208 1532
rect 35250 1492 35290 1532
rect 35332 1492 35372 1532
rect 35414 1492 35454 1532
rect 35496 1492 35536 1532
rect 1420 1240 1460 1280
rect 18508 904 18548 944
rect 45676 904 45716 944
rect 18604 568 18644 608
rect 44620 568 44660 608
<< metal3 >>
rect 9580 11780 9620 11789
rect 11000 11764 11080 11844
rect 11192 11764 11272 11844
rect 11384 11764 11464 11844
rect 11576 11764 11656 11844
rect 11768 11764 11848 11844
rect 11960 11764 12040 11844
rect 12152 11764 12232 11844
rect 12344 11764 12424 11844
rect 12536 11764 12616 11844
rect 12728 11764 12808 11844
rect 12920 11764 13000 11844
rect 13112 11764 13192 11844
rect 13304 11764 13384 11844
rect 13496 11764 13576 11844
rect 13688 11764 13768 11844
rect 13880 11764 13960 11844
rect 14072 11764 14152 11844
rect 14264 11764 14344 11844
rect 14456 11764 14536 11844
rect 14648 11764 14728 11844
rect 14840 11764 14920 11844
rect 15032 11764 15112 11844
rect 15224 11764 15304 11844
rect 15416 11764 15496 11844
rect 15608 11764 15688 11844
rect 15800 11764 15880 11844
rect 15992 11764 16072 11844
rect 16184 11764 16264 11844
rect 16376 11764 16456 11844
rect 16568 11764 16648 11844
rect 16760 11764 16840 11844
rect 16952 11764 17032 11844
rect 17144 11764 17224 11844
rect 17336 11764 17416 11844
rect 17528 11764 17608 11844
rect 17720 11764 17800 11844
rect 17912 11764 17992 11844
rect 18104 11764 18184 11844
rect 18296 11764 18376 11844
rect 18488 11764 18568 11844
rect 18680 11764 18760 11844
rect 18872 11764 18952 11844
rect 19064 11764 19144 11844
rect 19256 11764 19336 11844
rect 19448 11764 19528 11844
rect 19640 11764 19720 11844
rect 19832 11764 19912 11844
rect 20024 11764 20104 11844
rect 20216 11764 20296 11844
rect 20408 11764 20488 11844
rect 20600 11764 20680 11844
rect 20792 11764 20872 11844
rect 20984 11764 21064 11844
rect 21176 11764 21256 11844
rect 21368 11764 21448 11844
rect 21560 11764 21640 11844
rect 21752 11764 21832 11844
rect 21944 11764 22024 11844
rect 22136 11780 22216 11844
rect 22136 11764 22156 11780
rect 1324 11024 1364 11033
rect 268 10688 308 10697
rect 172 8336 212 8345
rect 172 7496 212 8296
rect 268 7916 308 10648
rect 556 10352 596 10361
rect 556 8672 596 10312
rect 556 8623 596 8632
rect 1324 8252 1364 10984
rect 1420 10016 1460 10025
rect 1420 9881 1460 9976
rect 3688 9848 4056 9857
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 3688 9799 4056 9808
rect 1420 9680 1460 9689
rect 1420 9545 1460 9640
rect 9484 9512 9524 9521
rect 8620 9428 8660 9437
rect 1420 9344 1460 9353
rect 1420 9209 1460 9304
rect 4928 9092 5296 9101
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 4928 9043 5296 9052
rect 1420 9008 1460 9017
rect 1420 8873 1460 8968
rect 1420 8756 1460 8765
rect 1420 8672 1460 8716
rect 1420 8621 1460 8632
rect 1324 8203 1364 8212
rect 2956 8420 2996 8429
rect 2860 8168 2900 8177
rect 2956 8168 2996 8380
rect 3688 8336 4056 8345
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 3688 8287 4056 8296
rect 2900 8128 2996 8168
rect 2860 8119 2900 8128
rect 268 7867 308 7876
rect 4780 7664 4820 7673
rect 4780 7529 4820 7624
rect 5548 7664 5588 7673
rect 4928 7580 5296 7589
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 4928 7531 5296 7540
rect 5548 7529 5588 7624
rect 172 7447 212 7456
rect 8620 7076 8660 9388
rect 8620 7027 8660 7036
rect 8716 8756 8756 8765
rect 7852 6992 7892 7001
rect 3688 6824 4056 6833
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 3688 6775 4056 6784
rect 6220 6488 6260 6497
rect 4108 6404 4148 6413
rect 748 6320 788 6329
rect 652 5312 692 5321
rect 652 2372 692 5272
rect 748 4892 788 6280
rect 1420 5648 1460 5657
rect 748 4843 788 4852
rect 1132 4976 1172 4985
rect 1132 3548 1172 4936
rect 1132 3499 1172 3508
rect 1228 4640 1268 4649
rect 1228 2792 1268 4600
rect 1420 3716 1460 5608
rect 1420 3667 1460 3676
rect 1996 5648 2036 5657
rect 1228 2743 1268 2752
rect 1324 3464 1364 3473
rect 652 2323 692 2332
rect 1324 1952 1364 3424
rect 1324 1903 1364 1912
rect 1420 3128 1460 3137
rect 1420 1280 1460 3088
rect 1420 1231 1460 1240
rect 1996 80 2036 5608
rect 3688 5312 4056 5321
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 3688 5263 4056 5272
rect 3688 3800 4056 3809
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 3688 3751 4056 3760
rect 2188 3380 2228 3389
rect 2188 3296 2228 3340
rect 2188 3245 2228 3256
rect 3688 2288 4056 2297
rect 3728 2248 3770 2288
rect 3810 2248 3852 2288
rect 3892 2248 3934 2288
rect 3974 2248 4016 2288
rect 3688 2239 4056 2248
rect 4108 80 4148 6364
rect 4928 6068 5296 6077
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 4928 6019 5296 6028
rect 4928 4556 5296 4565
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 4928 4507 5296 4516
rect 4928 3044 5296 3053
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 4928 2995 5296 3004
rect 4928 1532 5296 1541
rect 4968 1492 5010 1532
rect 5050 1492 5092 1532
rect 5132 1492 5174 1532
rect 5214 1492 5256 1532
rect 4928 1483 5296 1492
rect 6220 80 6260 6448
rect 7852 5900 7892 6952
rect 8044 6992 8084 7001
rect 8044 6656 8084 6952
rect 8044 6607 8084 6616
rect 8716 6572 8756 8716
rect 9100 8672 9140 8681
rect 8716 6523 8756 6532
rect 8812 6824 8852 6833
rect 8428 6488 8468 6497
rect 8428 6068 8468 6448
rect 8812 6488 8852 6784
rect 9100 6572 9140 8632
rect 9100 6523 9140 6532
rect 9484 6572 9524 9472
rect 9484 6523 9524 6532
rect 8812 6439 8852 6448
rect 8428 6019 8468 6028
rect 7852 5851 7892 5860
rect 9580 5648 9620 11740
rect 9868 11696 9908 11705
rect 9580 5599 9620 5608
rect 9772 9008 9812 9017
rect 9772 5564 9812 8968
rect 9868 5648 9908 11656
rect 9868 5599 9908 5608
rect 10060 11528 10100 11537
rect 9772 5515 9812 5524
rect 8332 4976 8372 4985
rect 8140 3296 8180 3305
rect 8140 2204 8180 3256
rect 8140 2155 8180 2164
rect 8332 80 8372 4936
rect 10060 4976 10100 11488
rect 10348 9596 10388 9605
rect 10156 9344 10196 9353
rect 10156 5564 10196 9304
rect 10156 5515 10196 5524
rect 10252 5648 10292 5657
rect 10252 5312 10292 5608
rect 10252 5263 10292 5272
rect 10348 5144 10388 9556
rect 11020 8924 11060 11764
rect 11212 9680 11252 11764
rect 11212 9631 11252 9640
rect 11308 9512 11348 9521
rect 11020 8875 11060 8884
rect 11212 9428 11252 9437
rect 10540 8840 10580 8849
rect 10540 5564 10580 8800
rect 10540 5515 10580 5524
rect 10636 5648 10676 5657
rect 10348 5095 10388 5104
rect 10060 4927 10100 4936
rect 10636 4808 10676 5608
rect 11020 5648 11060 5657
rect 11020 4976 11060 5608
rect 11212 5480 11252 9388
rect 11308 5648 11348 9472
rect 11404 8924 11444 11764
rect 11596 9680 11636 11764
rect 11596 9631 11636 9640
rect 11404 8875 11444 8884
rect 11788 8924 11828 11764
rect 11788 8875 11828 8884
rect 11884 11696 11924 11705
rect 11308 5599 11348 5608
rect 11500 8756 11540 8765
rect 11500 5564 11540 8716
rect 11500 5515 11540 5524
rect 11596 5648 11636 5657
rect 11212 5431 11252 5440
rect 11596 5060 11636 5608
rect 11884 5648 11924 11656
rect 11980 9680 12020 11764
rect 11980 9631 12020 9640
rect 12172 8924 12212 11764
rect 12364 9680 12404 11764
rect 12364 9631 12404 9640
rect 12172 8875 12212 8884
rect 12556 8924 12596 11764
rect 12748 9680 12788 11764
rect 12940 11444 12980 11764
rect 12940 11404 13076 11444
rect 12748 9631 12788 9640
rect 12556 8875 12596 8884
rect 11884 5599 11924 5608
rect 12460 8672 12500 8681
rect 12460 5564 12500 8632
rect 13036 8588 13076 11404
rect 13132 9680 13172 11764
rect 13132 9631 13172 9640
rect 13036 8539 13076 8548
rect 13228 9512 13268 9521
rect 12460 5515 12500 5524
rect 13228 5480 13268 9472
rect 13324 8924 13364 11764
rect 13516 9680 13556 11764
rect 13516 9631 13556 9640
rect 13324 8875 13364 8884
rect 13708 8924 13748 11764
rect 13900 9680 13940 11764
rect 13900 9631 13940 9640
rect 13708 8875 13748 8884
rect 13804 9512 13844 9521
rect 13516 8756 13556 8765
rect 13228 5431 13268 5440
rect 13324 5648 13364 5657
rect 11596 5011 11636 5020
rect 11020 4927 11060 4936
rect 10636 4759 10676 4768
rect 13324 4724 13364 5608
rect 13516 5564 13556 8716
rect 13612 8672 13652 8681
rect 13612 5648 13652 8632
rect 13612 5599 13652 5608
rect 13708 8000 13748 8009
rect 13516 5515 13556 5524
rect 13708 5564 13748 7960
rect 13708 5515 13748 5524
rect 13804 5144 13844 9472
rect 14092 8924 14132 11764
rect 14284 9680 14324 11764
rect 14284 9631 14324 9640
rect 14092 8875 14132 8884
rect 14188 9512 14228 9521
rect 13996 8672 14036 8681
rect 13996 5564 14036 8632
rect 14188 6572 14228 9472
rect 14188 6523 14228 6532
rect 14284 9428 14324 9437
rect 14284 5732 14324 9388
rect 14476 8924 14516 11764
rect 14668 9680 14708 11764
rect 14668 9631 14708 9640
rect 14476 8875 14516 8884
rect 14860 8924 14900 11764
rect 15052 9680 15092 11764
rect 15052 9631 15092 9640
rect 14860 8875 14900 8884
rect 15052 9512 15092 9521
rect 14284 5683 14324 5692
rect 14380 8672 14420 8681
rect 14380 5648 14420 8632
rect 14956 7916 14996 7925
rect 14380 5599 14420 5608
rect 14668 5648 14708 5657
rect 13996 5515 14036 5524
rect 14668 5480 14708 5608
rect 14956 5648 14996 7876
rect 14956 5599 14996 5608
rect 14860 5480 14900 5489
rect 14668 5440 14860 5480
rect 14860 5431 14900 5440
rect 13804 5095 13844 5104
rect 13324 4675 13364 4684
rect 13900 4976 13940 4985
rect 13900 4640 13940 4936
rect 13900 4591 13940 4600
rect 14188 4976 14228 4985
rect 14188 4388 14228 4936
rect 15052 4808 15092 9472
rect 15244 8924 15284 11764
rect 15244 8875 15284 8884
rect 15340 11024 15380 11033
rect 15148 8672 15188 8681
rect 15148 5732 15188 8632
rect 15340 6824 15380 10984
rect 15436 9680 15476 11764
rect 15436 9631 15476 9640
rect 15340 6775 15380 6784
rect 15436 9512 15476 9521
rect 15436 5816 15476 9472
rect 15628 8924 15668 11764
rect 15820 9680 15860 11764
rect 15820 9631 15860 9640
rect 15628 8875 15668 8884
rect 15724 9512 15764 9521
rect 15532 8672 15572 8681
rect 15532 6572 15572 8632
rect 15532 6523 15572 6532
rect 15724 6236 15764 9472
rect 16012 8924 16052 11764
rect 16204 9680 16244 11764
rect 16204 9631 16244 9640
rect 16300 11360 16340 11369
rect 16012 8875 16052 8884
rect 15916 8672 15956 8681
rect 15724 6187 15764 6196
rect 15820 6908 15860 6917
rect 15436 5767 15476 5776
rect 15820 5816 15860 6868
rect 15820 5767 15860 5776
rect 15148 5683 15188 5692
rect 15052 4759 15092 4768
rect 15340 5648 15380 5657
rect 15340 4640 15380 5608
rect 15916 4976 15956 8632
rect 16108 6656 16148 6665
rect 16108 5060 16148 6616
rect 16108 5011 16148 5020
rect 15916 4927 15956 4936
rect 15340 4591 15380 4600
rect 16300 4640 16340 11320
rect 16396 8924 16436 11764
rect 16396 8875 16436 8884
rect 16492 11612 16532 11621
rect 16492 5480 16532 11572
rect 16588 9680 16628 11764
rect 16588 9631 16628 9640
rect 16780 8924 16820 11764
rect 16972 9680 17012 11764
rect 16972 9631 17012 9640
rect 16780 8875 16820 8884
rect 16972 9512 17012 9521
rect 16684 8672 16724 8681
rect 16492 5431 16532 5440
rect 16588 8252 16628 8261
rect 16300 4591 16340 4600
rect 16588 4556 16628 8212
rect 16684 5060 16724 8632
rect 16780 8504 16820 8513
rect 16780 5144 16820 8464
rect 16876 6740 16916 6749
rect 16876 6404 16916 6700
rect 16876 6355 16916 6364
rect 16972 5564 17012 9472
rect 17164 8924 17204 11764
rect 17356 9680 17396 11764
rect 17356 9631 17396 9640
rect 17452 9512 17492 9521
rect 17164 8875 17204 8884
rect 17260 9428 17300 9437
rect 17164 8756 17204 8765
rect 17068 8672 17108 8681
rect 17068 6404 17108 8632
rect 17068 6355 17108 6364
rect 16972 5515 17012 5524
rect 17164 5480 17204 8716
rect 17260 5732 17300 9388
rect 17260 5683 17300 5692
rect 17164 5431 17204 5440
rect 16780 5095 16820 5104
rect 17452 5144 17492 9472
rect 17548 8924 17588 11764
rect 17644 9932 17684 9941
rect 17644 9512 17684 9892
rect 17740 9680 17780 11764
rect 17740 9631 17780 9640
rect 17644 9463 17684 9472
rect 17548 8875 17588 8884
rect 17932 8924 17972 11764
rect 18028 10100 18068 10109
rect 18028 9512 18068 10060
rect 18124 9680 18164 11764
rect 18124 9631 18164 9640
rect 18028 9463 18068 9472
rect 17932 8875 17972 8884
rect 18028 9344 18068 9353
rect 18028 5816 18068 9304
rect 18316 8924 18356 11764
rect 18508 9680 18548 11764
rect 18604 10100 18644 10109
rect 18604 9764 18644 10060
rect 18604 9715 18644 9724
rect 18508 9631 18548 9640
rect 18316 8875 18356 8884
rect 18700 8924 18740 11764
rect 18892 10100 18932 11764
rect 19084 10184 19124 11764
rect 19276 10268 19316 11764
rect 19276 10228 19412 10268
rect 19084 10144 19316 10184
rect 18892 10051 18932 10060
rect 18808 9848 19176 9857
rect 18848 9808 18890 9848
rect 18930 9808 18972 9848
rect 19012 9808 19054 9848
rect 19094 9808 19136 9848
rect 18808 9799 19176 9808
rect 18796 9680 18836 9689
rect 18836 9640 18932 9680
rect 18796 9631 18836 9640
rect 18700 8875 18740 8884
rect 18796 9512 18836 9521
rect 18124 8756 18164 8765
rect 18164 8716 18356 8756
rect 18124 8707 18164 8716
rect 18028 5767 18068 5776
rect 18124 6488 18164 6497
rect 18124 5648 18164 6448
rect 18124 5599 18164 5608
rect 18316 5396 18356 8716
rect 18796 8504 18836 9472
rect 18892 9092 18932 9640
rect 18892 9043 18932 9052
rect 19276 8924 19316 10144
rect 19372 9680 19412 10228
rect 19372 9631 19412 9640
rect 19276 8875 19316 8884
rect 19372 9512 19412 9521
rect 19372 8756 19412 9472
rect 19468 8924 19508 11764
rect 19468 8875 19508 8884
rect 19564 10268 19604 10277
rect 19564 8756 19604 10228
rect 19660 9596 19700 11764
rect 19660 9547 19700 9556
rect 19756 9428 19796 9437
rect 19756 9293 19796 9388
rect 18700 8464 18836 8504
rect 19276 8716 19412 8756
rect 19468 8716 19604 8756
rect 19756 9176 19796 9185
rect 18700 6992 18740 8464
rect 18808 8336 19176 8345
rect 18848 8296 18890 8336
rect 18930 8296 18972 8336
rect 19012 8296 19054 8336
rect 19094 8296 19136 8336
rect 18808 8287 19176 8296
rect 18700 6943 18740 6952
rect 18808 6824 19176 6833
rect 18848 6784 18890 6824
rect 18930 6784 18972 6824
rect 19012 6784 19054 6824
rect 19094 6784 19136 6824
rect 18808 6775 19176 6784
rect 18508 6572 18548 6581
rect 18508 5648 18548 6532
rect 19276 5984 19316 8716
rect 19372 6488 19412 6497
rect 19372 6152 19412 6448
rect 19372 6103 19412 6112
rect 19276 5944 19412 5984
rect 18604 5816 18644 5825
rect 18604 5681 18644 5776
rect 18508 5599 18548 5608
rect 19276 5648 19316 5657
rect 18508 5396 18548 5405
rect 18316 5356 18508 5396
rect 18508 5347 18548 5356
rect 18808 5312 19176 5321
rect 18848 5272 18890 5312
rect 18930 5272 18972 5312
rect 19012 5272 19054 5312
rect 19094 5272 19136 5312
rect 18808 5263 19176 5272
rect 17452 5095 17492 5104
rect 16684 5011 16724 5020
rect 19180 4976 19220 4985
rect 19180 4841 19220 4936
rect 19276 4808 19316 5608
rect 19276 4759 19316 4768
rect 16588 4507 16628 4516
rect 16780 4724 16820 4733
rect 14188 4339 14228 4348
rect 14668 4052 14708 4061
rect 10060 3380 10100 3389
rect 10060 3245 10100 3340
rect 10444 2624 10484 2633
rect 10444 80 10484 2584
rect 12556 2624 12596 2633
rect 12556 80 12596 2584
rect 14668 80 14708 4012
rect 16780 80 16820 4684
rect 19372 4388 19412 5944
rect 19468 4724 19508 8716
rect 19756 8672 19796 9136
rect 19852 8924 19892 11764
rect 19948 10688 19988 10697
rect 19948 9512 19988 10648
rect 19948 9463 19988 9472
rect 20044 9428 20084 11764
rect 20236 9680 20276 11764
rect 20236 9631 20276 9640
rect 20428 9596 20468 11764
rect 20428 9547 20468 9556
rect 20524 10016 20564 10025
rect 20044 9379 20084 9388
rect 19852 8875 19892 8884
rect 19948 9092 19988 9101
rect 19756 8623 19796 8632
rect 19852 6824 19892 6833
rect 19852 6068 19892 6784
rect 19852 6019 19892 6028
rect 19660 5648 19700 5657
rect 19468 4675 19508 4684
rect 19564 4976 19604 4985
rect 19372 4339 19412 4348
rect 19564 4388 19604 4936
rect 19660 4808 19700 5608
rect 19852 5648 19892 5657
rect 19852 5564 19892 5608
rect 19852 5513 19892 5524
rect 19948 5060 19988 9052
rect 20048 9092 20416 9101
rect 20088 9052 20130 9092
rect 20170 9052 20212 9092
rect 20252 9052 20294 9092
rect 20334 9052 20376 9092
rect 20048 9043 20416 9052
rect 20524 8840 20564 9976
rect 20620 9680 20660 11764
rect 20620 9631 20660 9640
rect 20716 10100 20756 10109
rect 20716 9344 20756 10060
rect 20812 9764 20852 11764
rect 20812 9715 20852 9724
rect 20716 9304 20948 9344
rect 20620 9176 20660 9185
rect 20812 9176 20852 9185
rect 20660 9136 20812 9176
rect 20620 9127 20660 9136
rect 20812 9127 20852 9136
rect 20524 8791 20564 8800
rect 20524 8588 20564 8597
rect 20140 8084 20180 8093
rect 20140 7949 20180 8044
rect 20048 7580 20416 7589
rect 20088 7540 20130 7580
rect 20170 7540 20212 7580
rect 20252 7540 20294 7580
rect 20334 7540 20376 7580
rect 20048 7531 20416 7540
rect 20048 6068 20416 6077
rect 20088 6028 20130 6068
rect 20170 6028 20212 6068
rect 20252 6028 20294 6068
rect 20334 6028 20376 6068
rect 20048 6019 20416 6028
rect 20044 5732 20084 5741
rect 20044 5396 20084 5692
rect 20524 5732 20564 8548
rect 20908 8084 20948 9304
rect 21004 9260 21044 11764
rect 21004 9211 21044 9220
rect 20908 8035 20948 8044
rect 21196 7160 21236 11764
rect 21196 7111 21236 7120
rect 21388 6824 21428 11764
rect 21388 6775 21428 6784
rect 21580 6740 21620 11764
rect 21772 11024 21812 11764
rect 21964 11528 22004 11764
rect 22196 11764 22216 11780
rect 22328 11764 22408 11844
rect 22520 11764 22600 11844
rect 22712 11764 22792 11844
rect 22904 11764 22984 11844
rect 23096 11764 23176 11844
rect 23288 11764 23368 11844
rect 23480 11764 23560 11844
rect 23672 11764 23752 11844
rect 23864 11764 23944 11844
rect 24056 11764 24136 11844
rect 24248 11764 24328 11844
rect 24440 11764 24520 11844
rect 24632 11764 24712 11844
rect 24824 11764 24904 11844
rect 25016 11764 25096 11844
rect 25208 11764 25288 11844
rect 25400 11764 25480 11844
rect 25592 11764 25672 11844
rect 25784 11764 25864 11844
rect 25976 11764 26056 11844
rect 26168 11764 26248 11844
rect 26360 11764 26440 11844
rect 26552 11764 26632 11844
rect 26744 11764 26824 11844
rect 26936 11764 27016 11844
rect 27128 11764 27208 11844
rect 27320 11764 27400 11844
rect 27512 11764 27592 11844
rect 27704 11764 27784 11844
rect 27896 11764 27976 11844
rect 28088 11764 28168 11844
rect 28280 11764 28360 11844
rect 28472 11764 28552 11844
rect 28664 11764 28744 11844
rect 28856 11764 28936 11844
rect 29048 11764 29128 11844
rect 29240 11764 29320 11844
rect 29432 11764 29512 11844
rect 29624 11764 29704 11844
rect 29816 11764 29896 11844
rect 30008 11764 30088 11844
rect 30200 11764 30280 11844
rect 30392 11764 30472 11844
rect 30584 11764 30664 11844
rect 30776 11764 30856 11844
rect 30968 11764 31048 11844
rect 31160 11764 31240 11844
rect 31352 11764 31432 11844
rect 31544 11764 31624 11844
rect 31736 11764 31816 11844
rect 31928 11764 32008 11844
rect 32120 11764 32200 11844
rect 32312 11764 32392 11844
rect 32504 11764 32584 11844
rect 32696 11764 32776 11844
rect 32888 11764 32968 11844
rect 33080 11764 33160 11844
rect 33272 11764 33352 11844
rect 33464 11764 33544 11844
rect 33656 11764 33736 11844
rect 33848 11764 33928 11844
rect 34040 11764 34120 11844
rect 34232 11764 34312 11844
rect 34424 11764 34504 11844
rect 34616 11764 34696 11844
rect 34808 11764 34888 11844
rect 35000 11764 35080 11844
rect 22156 11731 22196 11740
rect 22348 11696 22388 11764
rect 22348 11647 22388 11656
rect 21964 11479 22004 11488
rect 21772 10975 21812 10984
rect 21676 9428 21716 9437
rect 21676 9092 21716 9388
rect 21676 9043 21716 9052
rect 21676 8924 21716 8933
rect 21676 8588 21716 8884
rect 21676 8539 21716 8548
rect 22540 8504 22580 11764
rect 22540 8455 22580 8464
rect 22732 8252 22772 11764
rect 22924 11696 22964 11764
rect 22924 11647 22964 11656
rect 22732 8203 22772 8212
rect 21580 6691 21620 6700
rect 23116 6656 23156 11764
rect 23308 11360 23348 11764
rect 23308 11311 23348 11320
rect 23116 6607 23156 6616
rect 23500 6572 23540 11764
rect 23692 10268 23732 11764
rect 23884 10688 23924 11764
rect 23884 10639 23924 10648
rect 23692 10219 23732 10228
rect 24076 6908 24116 11764
rect 24268 8924 24308 11764
rect 24460 11612 24500 11764
rect 24460 11563 24500 11572
rect 24076 6859 24116 6868
rect 24172 8884 24308 8924
rect 23500 6523 23540 6532
rect 21964 6152 22004 6161
rect 21964 5816 22004 6112
rect 21964 5767 22004 5776
rect 23116 5776 23348 5816
rect 20524 5683 20564 5692
rect 23020 5732 23060 5741
rect 23116 5732 23156 5776
rect 23060 5692 23156 5732
rect 23020 5683 23060 5692
rect 21196 5648 21236 5657
rect 20428 5564 20468 5573
rect 20428 5480 20468 5524
rect 20428 5429 20468 5440
rect 20716 5480 20756 5489
rect 20044 5347 20084 5356
rect 20716 5345 20756 5440
rect 21196 5228 21236 5608
rect 21772 5648 21812 5659
rect 21772 5564 21812 5608
rect 21772 5515 21812 5524
rect 23212 5648 23252 5657
rect 21196 5179 21236 5188
rect 21292 5480 21332 5489
rect 19948 5011 19988 5020
rect 21292 4976 21332 5440
rect 23020 5480 23060 5489
rect 23020 5312 23060 5440
rect 23020 5272 23156 5312
rect 22348 5144 22388 5153
rect 21676 5060 21716 5069
rect 21292 4927 21332 4936
rect 21484 5020 21676 5060
rect 21484 4976 21524 5020
rect 21676 5011 21716 5020
rect 21484 4927 21524 4936
rect 19660 4759 19700 4768
rect 20140 4724 20180 4819
rect 22348 4808 22388 5104
rect 22348 4759 22388 4768
rect 22540 4808 22580 4817
rect 20140 4675 20180 4684
rect 22540 4673 22580 4768
rect 19756 4640 19796 4649
rect 19756 4505 19796 4600
rect 23116 4640 23156 5272
rect 23116 4591 23156 4600
rect 20048 4556 20416 4565
rect 20088 4516 20130 4556
rect 20170 4516 20212 4556
rect 20252 4516 20294 4556
rect 20334 4516 20376 4556
rect 20048 4507 20416 4516
rect 19564 4339 19604 4348
rect 22924 4304 22964 4313
rect 17260 4220 17300 4229
rect 17260 2960 17300 4180
rect 20812 4220 20852 4229
rect 19276 4136 19316 4145
rect 18508 3884 18548 3893
rect 17932 3464 17972 3473
rect 17932 3128 17972 3424
rect 17932 3079 17972 3088
rect 17260 2911 17300 2920
rect 18508 944 18548 3844
rect 18808 3800 19176 3809
rect 18848 3760 18890 3800
rect 18930 3760 18972 3800
rect 19012 3760 19054 3800
rect 19094 3760 19136 3800
rect 18808 3751 19176 3760
rect 18700 3464 18740 3473
rect 18508 895 18548 904
rect 18604 3044 18644 3053
rect 18604 608 18644 3004
rect 18700 1616 18740 3424
rect 18808 2288 19176 2297
rect 18848 2248 18890 2288
rect 18930 2248 18972 2288
rect 19012 2248 19054 2288
rect 19094 2248 19136 2288
rect 18808 2239 19176 2248
rect 18700 1567 18740 1576
rect 18604 559 18644 568
rect 18892 148 19124 188
rect 18892 80 18932 148
rect 1976 0 2056 80
rect 4088 0 4168 80
rect 6200 0 6280 80
rect 8312 0 8392 80
rect 10424 0 10504 80
rect 12536 0 12616 80
rect 14648 0 14728 80
rect 16760 0 16840 80
rect 18872 0 18952 80
rect 19084 60 19124 148
rect 19276 60 19316 4096
rect 20812 4085 20852 4180
rect 21004 4220 21044 4229
rect 20140 3968 20180 3977
rect 20140 3833 20180 3928
rect 19852 3800 19892 3809
rect 19564 3212 19604 3221
rect 19564 2204 19604 3172
rect 19852 2900 19892 3760
rect 19948 3464 19988 3473
rect 19948 3044 19988 3424
rect 19948 2995 19988 3004
rect 20048 3044 20416 3053
rect 20088 3004 20130 3044
rect 20170 3004 20212 3044
rect 20252 3004 20294 3044
rect 20334 3004 20376 3044
rect 20048 2995 20416 3004
rect 19852 2860 19988 2900
rect 19948 2708 19988 2860
rect 19948 2659 19988 2668
rect 19564 2155 19604 2164
rect 20048 1532 20416 1541
rect 20088 1492 20130 1532
rect 20170 1492 20212 1532
rect 20252 1492 20294 1532
rect 20334 1492 20376 1532
rect 20048 1483 20416 1492
rect 21004 80 21044 4180
rect 22828 4136 22868 4145
rect 21676 4052 21716 4061
rect 21676 3917 21716 4012
rect 21868 4052 21908 4061
rect 21388 3884 21428 3893
rect 21388 3464 21428 3844
rect 21388 3415 21428 3424
rect 21772 3464 21812 3473
rect 21484 3212 21524 3221
rect 21484 2036 21524 3172
rect 21772 3044 21812 3424
rect 21868 3212 21908 4012
rect 22636 3800 22676 3809
rect 22636 3464 22676 3760
rect 22636 3415 22676 3424
rect 22828 3464 22868 4096
rect 22924 3548 22964 4264
rect 23020 4220 23060 4229
rect 23020 4085 23060 4180
rect 22924 3508 23156 3548
rect 22828 3415 22868 3424
rect 22924 3380 22964 3389
rect 22924 3296 22964 3340
rect 22924 3245 22964 3256
rect 23116 3296 23156 3508
rect 23116 3247 23156 3256
rect 21868 3163 21908 3172
rect 21772 2995 21812 3004
rect 23020 2960 23060 3055
rect 23116 3044 23156 3139
rect 23116 2995 23156 3004
rect 23020 2911 23060 2920
rect 23212 2900 23252 5608
rect 23308 5480 23348 5776
rect 23308 5431 23348 5440
rect 24172 4556 24212 8884
rect 24268 8756 24308 8765
rect 24268 8168 24308 8716
rect 24268 8119 24308 8128
rect 24652 7916 24692 11764
rect 24844 8000 24884 11764
rect 25036 9092 25076 11764
rect 24844 7951 24884 7960
rect 24940 9052 25076 9092
rect 25132 9092 25172 9101
rect 24652 7867 24692 7876
rect 24844 6068 24884 6077
rect 24844 5816 24884 6028
rect 24844 5767 24884 5776
rect 24940 5312 24980 9052
rect 25036 8924 25076 8933
rect 25036 7916 25076 8884
rect 25132 8000 25172 9052
rect 25132 7951 25172 7960
rect 25036 7867 25076 7876
rect 25036 5816 25076 5825
rect 25036 5396 25076 5776
rect 25228 5732 25268 11764
rect 25420 9260 25460 11764
rect 25228 5683 25268 5692
rect 25324 9220 25460 9260
rect 25324 5480 25364 9220
rect 25420 8000 25460 8009
rect 25420 7412 25460 7960
rect 25420 7363 25460 7372
rect 25324 5431 25364 5440
rect 25036 5347 25076 5356
rect 24940 5263 24980 5272
rect 25228 5312 25268 5321
rect 24172 4507 24212 4516
rect 24844 4220 24884 4229
rect 24076 3968 24116 3977
rect 23500 3380 23540 3389
rect 23500 3245 23540 3340
rect 23404 3212 23444 3221
rect 23404 3077 23444 3172
rect 24076 3044 24116 3928
rect 24076 2995 24116 3004
rect 24172 3548 24212 3557
rect 24172 2960 24212 3508
rect 24844 3464 24884 4180
rect 24844 3415 24884 3424
rect 24172 2911 24212 2920
rect 21484 1987 21524 1996
rect 23116 2860 23252 2900
rect 23116 80 23156 2860
rect 25228 80 25268 5272
rect 25612 5144 25652 11764
rect 25804 10184 25844 11764
rect 25612 5095 25652 5104
rect 25708 10144 25844 10184
rect 25708 4976 25748 10144
rect 25900 8672 25940 8681
rect 25900 8168 25940 8632
rect 25900 8119 25940 8128
rect 25900 8000 25940 8009
rect 25900 7580 25940 7960
rect 25900 7531 25940 7540
rect 25996 6404 26036 11764
rect 26188 8588 26228 11764
rect 26380 10268 26420 11764
rect 26572 11024 26612 11764
rect 25996 6355 26036 6364
rect 26092 8548 26228 8588
rect 26284 10228 26420 10268
rect 26476 10984 26612 11024
rect 25708 4927 25748 4936
rect 25996 4808 26036 4817
rect 26092 4808 26132 8548
rect 26188 8420 26228 8429
rect 26188 8000 26228 8380
rect 26188 7951 26228 7960
rect 26284 5228 26324 10228
rect 26380 8840 26420 8849
rect 26380 8705 26420 8800
rect 26476 6488 26516 10984
rect 26668 9176 26708 9185
rect 26572 8420 26612 8429
rect 26572 8000 26612 8380
rect 26668 8168 26708 9136
rect 26668 8119 26708 8128
rect 26572 7951 26612 7960
rect 26476 6439 26516 6448
rect 26764 5396 26804 11764
rect 26956 8588 26996 11764
rect 26860 8548 26996 8588
rect 27052 9932 27092 9941
rect 26860 5732 26900 8548
rect 26956 8336 26996 8345
rect 26956 8000 26996 8296
rect 27052 8168 27092 9892
rect 27052 8119 27092 8128
rect 26956 7951 26996 7960
rect 26860 5683 26900 5692
rect 26764 5347 26804 5356
rect 26284 5179 26324 5188
rect 26036 4768 26132 4808
rect 25996 4759 26036 4768
rect 27148 4640 27188 11764
rect 27340 11696 27380 11764
rect 27340 11647 27380 11656
rect 27532 10016 27572 11764
rect 27436 9976 27572 10016
rect 27628 11696 27668 11705
rect 27340 9512 27380 9521
rect 27244 9176 27284 9185
rect 27244 8756 27284 9136
rect 27244 8707 27284 8716
rect 27244 8000 27284 8009
rect 27244 7865 27284 7960
rect 27340 7748 27380 9472
rect 27340 7699 27380 7708
rect 27436 6068 27476 9976
rect 27532 9848 27572 9857
rect 27532 8924 27572 9808
rect 27532 8875 27572 8884
rect 27532 8084 27572 8093
rect 27532 7949 27572 8044
rect 27436 6019 27476 6028
rect 27148 4591 27188 4600
rect 27340 5732 27380 5741
rect 25804 4136 25844 4145
rect 25804 4052 25844 4096
rect 25804 4001 25844 4012
rect 26284 4136 26324 4145
rect 25900 3884 25940 3893
rect 25804 3844 25900 3884
rect 25804 3548 25844 3844
rect 25900 3835 25940 3844
rect 25804 3499 25844 3508
rect 26284 3212 26324 4096
rect 26764 3968 26804 3977
rect 26764 3464 26804 3928
rect 26764 3415 26804 3424
rect 26284 3163 26324 3172
rect 27340 2900 27380 5692
rect 27628 4472 27668 11656
rect 27724 6572 27764 11764
rect 27916 9512 27956 11764
rect 27724 6523 27764 6532
rect 27820 9472 27956 9512
rect 27820 6488 27860 9472
rect 28012 9428 28052 9437
rect 27916 9344 27956 9353
rect 27916 8840 27956 9304
rect 27916 8791 27956 8800
rect 28012 8672 28052 9388
rect 28012 8623 28052 8632
rect 28108 8000 28148 11764
rect 28300 8840 28340 11764
rect 28300 8791 28340 8800
rect 28492 8672 28532 11764
rect 28684 8756 28724 11764
rect 28684 8707 28724 8716
rect 28780 9596 28820 9605
rect 28492 8623 28532 8632
rect 28780 8672 28820 9556
rect 28876 8924 28916 11764
rect 28876 8875 28916 8884
rect 28780 8623 28820 8632
rect 28108 7951 28148 7960
rect 29068 7916 29108 11764
rect 29068 7867 29108 7876
rect 29164 8756 29204 8765
rect 27820 6439 27860 6448
rect 27628 4423 27668 4432
rect 28012 3800 28052 3809
rect 28012 2960 28052 3760
rect 28012 2911 28052 2920
rect 28780 3212 28820 3221
rect 28780 2960 28820 3172
rect 28780 2911 28820 2920
rect 29164 2900 29204 8716
rect 29260 8000 29300 11764
rect 29452 8336 29492 11764
rect 29452 8287 29492 8296
rect 29260 7951 29300 7960
rect 29644 7160 29684 11764
rect 29836 8504 29876 11764
rect 30028 9932 30068 11764
rect 29836 8455 29876 8464
rect 29932 9892 30068 9932
rect 29932 7412 29972 9892
rect 29932 7363 29972 7372
rect 30028 8672 30068 8681
rect 29644 7111 29684 7120
rect 27244 2860 27380 2900
rect 28876 2876 29204 2900
rect 27244 440 27284 2860
rect 28916 2860 29204 2876
rect 29548 5732 29588 5741
rect 28876 2827 28916 2836
rect 29548 608 29588 5692
rect 29836 5648 29876 5657
rect 29836 5312 29876 5608
rect 30028 5648 30068 8632
rect 30220 7580 30260 11764
rect 30412 8420 30452 11764
rect 30412 8371 30452 8380
rect 30508 9932 30548 9941
rect 30220 7531 30260 7540
rect 30028 5599 30068 5608
rect 29836 5263 29876 5272
rect 29932 5480 29972 5489
rect 29932 5060 29972 5440
rect 30508 5480 30548 9892
rect 30604 9176 30644 11764
rect 30604 9127 30644 9136
rect 30796 9092 30836 11764
rect 30796 9043 30836 9052
rect 30892 9344 30932 9353
rect 30508 5431 30548 5440
rect 30892 5480 30932 9304
rect 30988 9008 31028 11764
rect 31180 9680 31220 11764
rect 31180 9631 31220 9640
rect 31372 9596 31412 11764
rect 31564 9680 31604 11764
rect 31564 9631 31604 9640
rect 31372 9547 31412 9556
rect 31756 9596 31796 11764
rect 31948 9764 31988 11764
rect 31948 9715 31988 9724
rect 31756 9547 31796 9556
rect 30988 8959 31028 8968
rect 31468 9512 31508 9521
rect 31468 5564 31508 9472
rect 31660 9512 31700 9521
rect 31660 6320 31700 9472
rect 32044 9512 32084 9521
rect 31660 6271 31700 6280
rect 31756 9176 31796 9185
rect 31468 5515 31508 5524
rect 31564 5648 31604 5657
rect 30892 5431 30932 5440
rect 29932 5011 29972 5020
rect 29452 568 29588 608
rect 27244 400 27380 440
rect 27340 80 27380 400
rect 29452 80 29492 568
rect 31564 80 31604 5608
rect 31756 4304 31796 9136
rect 31948 9092 31988 9101
rect 31852 8672 31892 8681
rect 31852 8252 31892 8632
rect 31852 8203 31892 8212
rect 31948 4556 31988 9052
rect 32044 7076 32084 9472
rect 32140 8924 32180 11764
rect 32332 9848 32372 11764
rect 32332 9799 32372 9808
rect 32428 10016 32468 10025
rect 32140 8875 32180 8884
rect 32236 9428 32276 9437
rect 32044 7027 32084 7036
rect 32044 5648 32084 5657
rect 32044 5144 32084 5608
rect 32044 5095 32084 5104
rect 31948 4507 31988 4516
rect 31756 4255 31796 4264
rect 31756 4136 31796 4145
rect 31756 3632 31796 4096
rect 31756 3583 31796 3592
rect 31852 3716 31892 3725
rect 31852 3464 31892 3676
rect 31852 3415 31892 3424
rect 32236 2120 32276 9388
rect 32332 9260 32372 9269
rect 32332 4136 32372 9220
rect 32428 4724 32468 9976
rect 32524 8924 32564 11764
rect 32524 8875 32564 8884
rect 32620 10100 32660 10109
rect 32620 5480 32660 10060
rect 32716 9596 32756 11764
rect 32716 9547 32756 9556
rect 32812 9512 32852 9521
rect 32812 9092 32852 9472
rect 32812 9043 32852 9052
rect 32908 8924 32948 11764
rect 33100 11444 33140 11764
rect 33100 11404 33236 11444
rect 33004 9848 33044 9857
rect 33004 9260 33044 9808
rect 33100 9428 33140 9437
rect 33100 9293 33140 9388
rect 33004 9211 33044 9220
rect 33196 9092 33236 11404
rect 33196 9043 33236 9052
rect 32908 8875 32948 8884
rect 33292 8924 33332 11764
rect 33484 9596 33524 11764
rect 33676 9680 33716 11764
rect 33868 10352 33908 11764
rect 33676 9631 33716 9640
rect 33772 10312 33908 10352
rect 33484 9556 33620 9596
rect 33484 9428 33524 9437
rect 33484 9293 33524 9388
rect 33580 9344 33620 9556
rect 33580 9295 33620 9304
rect 33772 9176 33812 10312
rect 34060 10016 34100 11764
rect 34252 10016 34292 11764
rect 34252 9976 34388 10016
rect 34060 9967 34100 9976
rect 33928 9848 34296 9857
rect 33968 9808 34010 9848
rect 34050 9808 34092 9848
rect 34132 9808 34174 9848
rect 34214 9808 34256 9848
rect 33928 9799 34296 9808
rect 33772 9127 33812 9136
rect 33868 9680 33908 9689
rect 33292 8875 33332 8884
rect 33196 8840 33236 8849
rect 32812 8672 32852 8681
rect 32716 8000 32756 8009
rect 32716 7328 32756 7960
rect 32716 7279 32756 7288
rect 32620 5431 32660 5440
rect 32812 4808 32852 8632
rect 32812 4759 32852 4768
rect 33004 8672 33044 8681
rect 32428 4675 32468 4684
rect 33004 4220 33044 8632
rect 33100 5396 33140 5405
rect 33196 5396 33236 8800
rect 33388 8756 33428 8765
rect 33292 7160 33332 7169
rect 33292 5900 33332 7120
rect 33292 5851 33332 5860
rect 33388 5648 33428 8716
rect 33868 8672 33908 9640
rect 33964 9512 34004 9521
rect 33964 8840 34004 9472
rect 34252 9344 34292 9353
rect 34252 8924 34292 9304
rect 34252 8875 34292 8884
rect 33964 8791 34004 8800
rect 34348 8840 34388 9976
rect 34444 9344 34484 11764
rect 34444 9295 34484 9304
rect 34540 10016 34580 10025
rect 34540 9176 34580 9976
rect 34540 9127 34580 9136
rect 34348 8791 34388 8800
rect 34444 9092 34484 9101
rect 33868 8623 33908 8632
rect 34348 8672 34388 8681
rect 33928 8336 34296 8345
rect 33968 8296 34010 8336
rect 34050 8296 34092 8336
rect 34132 8296 34174 8336
rect 34214 8296 34256 8336
rect 33928 8287 34296 8296
rect 34348 8000 34388 8632
rect 34348 7951 34388 7960
rect 33928 6824 34296 6833
rect 33968 6784 34010 6824
rect 34050 6784 34092 6824
rect 34132 6784 34174 6824
rect 34214 6784 34256 6824
rect 33928 6775 34296 6784
rect 34444 6152 34484 9052
rect 34636 8840 34676 11764
rect 34828 10016 34868 11764
rect 34828 9967 34868 9976
rect 35020 9596 35060 11764
rect 44140 11024 44180 11033
rect 43372 10688 43412 10697
rect 36076 10100 36116 10109
rect 35020 9547 35060 9556
rect 35692 9932 35732 9941
rect 34732 9512 34772 9521
rect 35692 9512 35732 9892
rect 34772 9472 34868 9512
rect 34732 9463 34772 9472
rect 34636 8791 34676 8800
rect 34348 6112 34484 6152
rect 34732 8672 34772 8681
rect 33388 5599 33428 5608
rect 33772 5648 33812 5657
rect 33140 5356 33236 5396
rect 33100 5328 33140 5356
rect 33004 4171 33044 4180
rect 33676 4892 33716 4901
rect 32332 4087 32372 4096
rect 33196 4052 33236 4061
rect 32428 3464 32468 3473
rect 32428 3128 32468 3424
rect 33100 3380 33140 3389
rect 33196 3380 33236 4012
rect 33140 3340 33236 3380
rect 33388 3380 33428 3389
rect 33428 3340 33524 3380
rect 33100 3312 33140 3340
rect 33388 3331 33428 3340
rect 33484 3296 33524 3340
rect 33484 3247 33524 3256
rect 32428 3079 32468 3088
rect 33388 3212 33428 3221
rect 33388 2960 33428 3172
rect 33388 2911 33428 2920
rect 32236 2071 32276 2080
rect 33676 80 33716 4852
rect 33772 4808 33812 5608
rect 34348 5648 34388 6112
rect 34348 5599 34388 5608
rect 34444 5984 34484 5993
rect 33928 5312 34296 5321
rect 33968 5272 34010 5312
rect 34050 5272 34092 5312
rect 34132 5272 34174 5312
rect 34214 5272 34256 5312
rect 33928 5263 34296 5272
rect 33772 4759 33812 4768
rect 34444 4136 34484 5944
rect 34732 5144 34772 8632
rect 34732 5095 34772 5104
rect 34828 5060 34868 9472
rect 35692 9463 35732 9472
rect 36076 9512 36116 10060
rect 43372 9680 43412 10648
rect 43372 9631 43412 9640
rect 43660 10352 43700 10361
rect 43660 9680 43700 10312
rect 43660 9631 43700 9640
rect 36076 9463 36116 9472
rect 36364 9596 36404 9605
rect 35596 9428 35636 9437
rect 35020 9092 35060 9101
rect 35020 8924 35060 9052
rect 35168 9092 35536 9101
rect 35208 9052 35250 9092
rect 35290 9052 35332 9092
rect 35372 9052 35414 9092
rect 35454 9052 35496 9092
rect 35168 9043 35536 9052
rect 35020 8875 35060 8884
rect 35212 7832 35252 7927
rect 35212 7783 35252 7792
rect 35168 7580 35536 7589
rect 35208 7540 35250 7580
rect 35290 7540 35332 7580
rect 35372 7540 35414 7580
rect 35454 7540 35496 7580
rect 35168 7531 35536 7540
rect 35168 6068 35536 6077
rect 35208 6028 35250 6068
rect 35290 6028 35332 6068
rect 35372 6028 35414 6068
rect 35454 6028 35496 6068
rect 35168 6019 35536 6028
rect 35596 5648 35636 9388
rect 35980 9344 36020 9353
rect 35788 9260 35828 9269
rect 35788 8756 35828 9220
rect 35788 8672 35828 8716
rect 35980 8756 36020 9304
rect 35980 8707 36020 8716
rect 36364 9176 36404 9556
rect 36748 9596 36788 9605
rect 35788 8621 35828 8632
rect 36076 8672 36116 8681
rect 35692 7664 35732 7673
rect 35692 7160 35732 7624
rect 36076 7412 36116 8632
rect 36364 8672 36404 9136
rect 36460 9512 36500 9521
rect 36460 8924 36500 9472
rect 36460 8875 36500 8884
rect 36748 8924 36788 9556
rect 37708 9512 37748 9521
rect 42988 9512 43028 9521
rect 37748 9472 38036 9512
rect 37708 9463 37748 9472
rect 36748 8875 36788 8884
rect 36940 9428 36980 9437
rect 36940 8756 36980 9388
rect 37996 9260 38036 9472
rect 37996 9211 38036 9220
rect 40204 9260 40244 9269
rect 37804 9176 37844 9185
rect 37228 9008 37268 9017
rect 37228 8924 37268 8968
rect 37228 8873 37268 8884
rect 37804 8924 37844 9136
rect 37804 8875 37844 8884
rect 37900 9092 37940 9101
rect 40108 9092 40148 9101
rect 36940 8707 36980 8716
rect 37420 8756 37460 8765
rect 36364 8623 36404 8632
rect 36172 8000 36212 8009
rect 36172 7916 36212 7960
rect 36172 7865 36212 7876
rect 36460 8000 36500 8009
rect 36460 7496 36500 7960
rect 37420 8000 37460 8716
rect 37420 7951 37460 7960
rect 37900 8672 37940 9052
rect 39916 9052 40108 9092
rect 39916 9008 39956 9052
rect 40108 9043 40148 9052
rect 39916 8959 39956 8968
rect 39820 8924 39860 8933
rect 39820 8789 39860 8884
rect 37900 8000 37940 8632
rect 37900 7951 37940 7960
rect 38668 8672 38708 8681
rect 38668 8000 38708 8632
rect 40204 8672 40244 9220
rect 40300 8924 40340 8933
rect 40300 8789 40340 8884
rect 40204 8623 40244 8632
rect 40492 8672 40532 8681
rect 40492 8168 40532 8632
rect 40492 8119 40532 8128
rect 42988 8168 43028 9472
rect 43372 9512 43412 9521
rect 43372 8840 43412 9472
rect 43756 9512 43796 9521
rect 43756 8924 43796 9472
rect 43756 8875 43796 8884
rect 43948 9428 43988 9437
rect 43372 8791 43412 8800
rect 43948 8672 43988 9388
rect 44140 8924 44180 10984
rect 44140 8875 44180 8884
rect 44428 10016 44468 10025
rect 44428 8924 44468 9976
rect 44428 8875 44468 8884
rect 45772 9260 45812 9269
rect 43948 8623 43988 8632
rect 45772 8672 45812 9220
rect 45772 8623 45812 8632
rect 42988 8119 43028 8128
rect 45772 8504 45812 8513
rect 38668 7951 38708 7960
rect 43564 8000 43604 8009
rect 36940 7916 36980 7925
rect 36940 7781 36980 7876
rect 40300 7832 40340 7841
rect 40300 7697 40340 7792
rect 36460 7447 36500 7456
rect 36076 7363 36116 7372
rect 35692 6488 35732 7120
rect 43564 7160 43604 7960
rect 45772 8000 45812 8464
rect 45772 7951 45812 7960
rect 45772 7748 45812 7757
rect 45772 7328 45812 7708
rect 45772 7279 45812 7288
rect 43564 7111 43604 7120
rect 44524 7160 44564 7169
rect 35692 6439 35732 6448
rect 41740 6488 41780 6497
rect 35596 5599 35636 5608
rect 40780 5648 40820 5657
rect 40012 5480 40052 5489
rect 34828 5011 34868 5020
rect 37900 5396 37940 5405
rect 35788 4976 35828 4985
rect 35168 4556 35536 4565
rect 35208 4516 35250 4556
rect 35290 4516 35332 4556
rect 35372 4516 35414 4556
rect 35454 4516 35496 4556
rect 35168 4507 35536 4516
rect 33928 3800 34296 3809
rect 33968 3760 34010 3800
rect 34050 3760 34092 3800
rect 34132 3760 34174 3800
rect 34214 3760 34256 3800
rect 33928 3751 34296 3760
rect 34444 3212 34484 4096
rect 34444 3163 34484 3172
rect 35168 3044 35536 3053
rect 35208 3004 35250 3044
rect 35290 3004 35332 3044
rect 35372 3004 35414 3044
rect 35454 3004 35496 3044
rect 35168 2995 35536 3004
rect 33928 2288 34296 2297
rect 33968 2248 34010 2288
rect 34050 2248 34092 2288
rect 34132 2248 34174 2288
rect 34214 2248 34256 2288
rect 33928 2239 34296 2248
rect 35168 1532 35536 1541
rect 35208 1492 35250 1532
rect 35290 1492 35332 1532
rect 35372 1492 35414 1532
rect 35454 1492 35496 1532
rect 35168 1483 35536 1492
rect 35788 80 35828 4936
rect 37900 80 37940 5356
rect 38764 4220 38804 4229
rect 38572 3968 38612 3977
rect 38572 1952 38612 3928
rect 38572 1903 38612 1912
rect 38764 1868 38804 4180
rect 38860 3716 38900 3725
rect 38860 2708 38900 3676
rect 38860 2659 38900 2668
rect 38764 1819 38804 1828
rect 40012 80 40052 5440
rect 40300 4136 40340 4145
rect 40300 4001 40340 4096
rect 40300 2960 40340 2969
rect 40300 2825 40340 2920
rect 40780 2456 40820 5608
rect 40876 4976 40916 4985
rect 40876 2540 40916 4936
rect 41740 4304 41780 6448
rect 44524 6152 44564 7120
rect 44524 6103 44564 6112
rect 44908 6488 44948 6497
rect 44236 5732 44276 5741
rect 43276 5564 43316 5573
rect 43180 4892 43220 4901
rect 43084 4852 43180 4892
rect 41740 4255 41780 4264
rect 42124 4808 42164 4817
rect 40876 2491 40916 2500
rect 40780 2407 40820 2416
rect 42124 80 42164 4768
rect 43084 3464 43124 4852
rect 43180 4843 43220 4852
rect 43276 3632 43316 5524
rect 43276 3583 43316 3592
rect 43084 3415 43124 3424
rect 44140 3044 44180 3053
rect 44140 2624 44180 3004
rect 44140 2575 44180 2584
rect 44236 80 44276 5692
rect 44908 5228 44948 6448
rect 46252 6152 46292 6161
rect 46252 5984 46292 6112
rect 46252 5935 46292 5944
rect 46252 5480 46292 5489
rect 46252 5312 46292 5440
rect 46252 5263 46292 5272
rect 44908 5179 44948 5188
rect 44620 3128 44660 3137
rect 44620 2036 44660 3088
rect 44620 1987 44660 1996
rect 45676 1784 45716 1793
rect 44620 1700 44660 1709
rect 44620 608 44660 1660
rect 45676 944 45716 1744
rect 45676 895 45716 904
rect 44620 559 44660 568
rect 19084 20 19316 60
rect 20984 0 21064 80
rect 23096 0 23176 80
rect 25208 0 25288 80
rect 27320 0 27400 80
rect 29432 0 29512 80
rect 31544 0 31624 80
rect 33656 0 33736 80
rect 35768 0 35848 80
rect 37880 0 37960 80
rect 39992 0 40072 80
rect 42104 0 42184 80
rect 44216 0 44296 80
<< via3 >>
rect 556 8632 596 8672
rect 1420 9976 1460 10016
rect 3688 9808 3728 9848
rect 3770 9808 3810 9848
rect 3852 9808 3892 9848
rect 3934 9808 3974 9848
rect 4016 9808 4056 9848
rect 1420 9640 1460 9680
rect 1420 9304 1460 9344
rect 4928 9052 4968 9092
rect 5010 9052 5050 9092
rect 5092 9052 5132 9092
rect 5174 9052 5214 9092
rect 5256 9052 5296 9092
rect 1420 8968 1460 9008
rect 1420 8716 1460 8756
rect 3688 8296 3728 8336
rect 3770 8296 3810 8336
rect 3852 8296 3892 8336
rect 3934 8296 3974 8336
rect 4016 8296 4056 8336
rect 4780 7624 4820 7664
rect 5548 7624 5588 7664
rect 4928 7540 4968 7580
rect 5010 7540 5050 7580
rect 5092 7540 5132 7580
rect 5174 7540 5214 7580
rect 5256 7540 5296 7580
rect 3688 6784 3728 6824
rect 3770 6784 3810 6824
rect 3852 6784 3892 6824
rect 3934 6784 3974 6824
rect 4016 6784 4056 6824
rect 3688 5272 3728 5312
rect 3770 5272 3810 5312
rect 3852 5272 3892 5312
rect 3934 5272 3974 5312
rect 4016 5272 4056 5312
rect 3688 3760 3728 3800
rect 3770 3760 3810 3800
rect 3852 3760 3892 3800
rect 3934 3760 3974 3800
rect 4016 3760 4056 3800
rect 2188 3340 2228 3380
rect 3688 2248 3728 2288
rect 3770 2248 3810 2288
rect 3852 2248 3892 2288
rect 3934 2248 3974 2288
rect 4016 2248 4056 2288
rect 4928 6028 4968 6068
rect 5010 6028 5050 6068
rect 5092 6028 5132 6068
rect 5174 6028 5214 6068
rect 5256 6028 5296 6068
rect 4928 4516 4968 4556
rect 5010 4516 5050 4556
rect 5092 4516 5132 4556
rect 5174 4516 5214 4556
rect 5256 4516 5296 4556
rect 4928 3004 4968 3044
rect 5010 3004 5050 3044
rect 5092 3004 5132 3044
rect 5174 3004 5214 3044
rect 5256 3004 5296 3044
rect 4928 1492 4968 1532
rect 5010 1492 5050 1532
rect 5092 1492 5132 1532
rect 5174 1492 5214 1532
rect 5256 1492 5296 1532
rect 11884 11656 11924 11696
rect 14956 7876 14996 7916
rect 15436 5776 15476 5816
rect 16108 6616 16148 6656
rect 15340 4600 15380 4640
rect 16972 5524 17012 5564
rect 17164 5440 17204 5480
rect 18604 10060 18644 10100
rect 18892 10060 18932 10100
rect 18808 9808 18848 9848
rect 18890 9808 18930 9848
rect 18972 9808 19012 9848
rect 19054 9808 19094 9848
rect 19136 9808 19176 9848
rect 18124 6448 18164 6488
rect 19372 9472 19412 9512
rect 19756 9388 19796 9428
rect 18808 8296 18848 8336
rect 18890 8296 18930 8336
rect 18972 8296 19012 8336
rect 19054 8296 19094 8336
rect 19136 8296 19176 8336
rect 18808 6784 18848 6824
rect 18890 6784 18930 6824
rect 18972 6784 19012 6824
rect 19054 6784 19094 6824
rect 19136 6784 19176 6824
rect 18508 6532 18548 6572
rect 18604 5776 18644 5816
rect 18808 5272 18848 5312
rect 18890 5272 18930 5312
rect 18972 5272 19012 5312
rect 19054 5272 19094 5312
rect 19136 5272 19176 5312
rect 19180 4936 19220 4976
rect 19276 4768 19316 4808
rect 16780 4684 16820 4724
rect 10060 3340 10100 3380
rect 19948 9472 19988 9512
rect 19852 5608 19892 5648
rect 20048 9052 20088 9092
rect 20130 9052 20170 9092
rect 20212 9052 20252 9092
rect 20294 9052 20334 9092
rect 20376 9052 20416 9092
rect 20524 8800 20564 8840
rect 20140 8044 20180 8084
rect 20048 7540 20088 7580
rect 20130 7540 20170 7580
rect 20212 7540 20252 7580
rect 20294 7540 20334 7580
rect 20376 7540 20416 7580
rect 20048 6028 20088 6068
rect 20130 6028 20170 6068
rect 20212 6028 20252 6068
rect 20294 6028 20334 6068
rect 20376 6028 20416 6068
rect 21676 9388 21716 9428
rect 22924 11656 22964 11696
rect 23116 6616 23156 6656
rect 20428 5524 20468 5564
rect 20716 5440 20756 5480
rect 21772 5608 21812 5648
rect 21292 4936 21332 4976
rect 22540 4768 22580 4808
rect 20140 4684 20180 4724
rect 19756 4600 19796 4640
rect 20048 4516 20088 4556
rect 20130 4516 20170 4556
rect 20212 4516 20252 4556
rect 20294 4516 20334 4556
rect 20376 4516 20416 4556
rect 20812 4180 20852 4220
rect 18808 3760 18848 3800
rect 18890 3760 18930 3800
rect 18972 3760 19012 3800
rect 19054 3760 19094 3800
rect 19136 3760 19176 3800
rect 18808 2248 18848 2288
rect 18890 2248 18930 2288
rect 18972 2248 19012 2288
rect 19054 2248 19094 2288
rect 19136 2248 19176 2288
rect 20140 3928 20180 3968
rect 20048 3004 20088 3044
rect 20130 3004 20170 3044
rect 20212 3004 20252 3044
rect 20294 3004 20334 3044
rect 20376 3004 20416 3044
rect 20048 1492 20088 1532
rect 20130 1492 20170 1532
rect 20212 1492 20252 1532
rect 20294 1492 20334 1532
rect 20376 1492 20416 1532
rect 21676 4012 21716 4052
rect 23020 4180 23060 4220
rect 22924 3340 22964 3380
rect 23116 3004 23156 3044
rect 23020 2920 23060 2960
rect 24652 7876 24692 7916
rect 23500 3340 23540 3380
rect 23404 3172 23444 3212
rect 24076 3004 24116 3044
rect 24172 2920 24212 2960
rect 26380 8800 26420 8840
rect 27340 11656 27380 11696
rect 27628 11656 27668 11696
rect 27244 7960 27284 8000
rect 27532 8044 27572 8084
rect 25804 4012 25844 4052
rect 26764 3928 26804 3968
rect 26284 3172 26324 3212
rect 27724 6532 27764 6572
rect 27820 6448 27860 6488
rect 29260 7960 29300 8000
rect 31756 4096 31796 4136
rect 33100 9388 33140 9428
rect 33484 9388 33524 9428
rect 34060 9976 34100 10016
rect 33928 9808 33968 9848
rect 34010 9808 34050 9848
rect 34092 9808 34132 9848
rect 34174 9808 34214 9848
rect 34256 9808 34296 9848
rect 33868 9640 33908 9680
rect 34252 9304 34292 9344
rect 34540 9976 34580 10016
rect 33928 8296 33968 8336
rect 34010 8296 34050 8336
rect 34092 8296 34132 8336
rect 34174 8296 34214 8336
rect 34256 8296 34296 8336
rect 33928 6784 33968 6824
rect 34010 6784 34050 6824
rect 34092 6784 34132 6824
rect 34174 6784 34214 6824
rect 34256 6784 34296 6824
rect 33388 2920 33428 2960
rect 33928 5272 33968 5312
rect 34010 5272 34050 5312
rect 34092 5272 34132 5312
rect 34174 5272 34214 5312
rect 34256 5272 34296 5312
rect 36364 9556 36404 9596
rect 35168 9052 35208 9092
rect 35250 9052 35290 9092
rect 35332 9052 35372 9092
rect 35414 9052 35454 9092
rect 35496 9052 35536 9092
rect 35212 7792 35252 7832
rect 35168 7540 35208 7580
rect 35250 7540 35290 7580
rect 35332 7540 35372 7580
rect 35414 7540 35454 7580
rect 35496 7540 35536 7580
rect 35168 6028 35208 6068
rect 35250 6028 35290 6068
rect 35332 6028 35372 6068
rect 35414 6028 35454 6068
rect 35496 6028 35536 6068
rect 35788 8716 35828 8756
rect 37228 8968 37268 9008
rect 36172 7876 36212 7916
rect 39820 8884 39860 8924
rect 37900 8632 37940 8672
rect 40300 8884 40340 8924
rect 36940 7876 36980 7916
rect 40300 7792 40340 7832
rect 35168 4516 35208 4556
rect 35250 4516 35290 4556
rect 35332 4516 35372 4556
rect 35414 4516 35454 4556
rect 35496 4516 35536 4556
rect 33928 3760 33968 3800
rect 34010 3760 34050 3800
rect 34092 3760 34132 3800
rect 34174 3760 34214 3800
rect 34256 3760 34296 3800
rect 35168 3004 35208 3044
rect 35250 3004 35290 3044
rect 35332 3004 35372 3044
rect 35414 3004 35454 3044
rect 35496 3004 35536 3044
rect 33928 2248 33968 2288
rect 34010 2248 34050 2288
rect 34092 2248 34132 2288
rect 34174 2248 34214 2288
rect 34256 2248 34296 2288
rect 35168 1492 35208 1532
rect 35250 1492 35290 1532
rect 35332 1492 35372 1532
rect 35414 1492 35454 1532
rect 35496 1492 35536 1532
rect 40300 4096 40340 4136
rect 40300 2920 40340 2960
<< metal4 >>
rect 11875 11656 11884 11696
rect 11924 11656 22924 11696
rect 22964 11656 22973 11696
rect 27331 11656 27340 11696
rect 27380 11656 27628 11696
rect 27668 11656 27677 11696
rect 18595 10060 18604 10100
rect 18644 10060 18892 10100
rect 18932 10060 18941 10100
rect 1411 9976 1420 10016
rect 1460 9976 33140 10016
rect 34051 9976 34060 10016
rect 34100 9976 34540 10016
rect 34580 9976 34589 10016
rect 3679 9808 3688 9848
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 4056 9808 4065 9848
rect 18799 9808 18808 9848
rect 18848 9808 18890 9848
rect 18930 9808 18972 9848
rect 19012 9808 19054 9848
rect 19094 9808 19136 9848
rect 19176 9808 19185 9848
rect 33100 9680 33140 9976
rect 33919 9808 33928 9848
rect 33968 9808 34010 9848
rect 34050 9808 34092 9848
rect 34132 9808 34174 9848
rect 34214 9808 34256 9848
rect 34296 9808 34305 9848
rect 1411 9640 1420 9680
rect 1460 9640 23060 9680
rect 33100 9640 33868 9680
rect 33908 9640 33917 9680
rect 23020 9596 23060 9640
rect 23020 9556 36364 9596
rect 36404 9556 36413 9596
rect 19363 9472 19372 9512
rect 19412 9472 19948 9512
rect 19988 9472 19997 9512
rect 19747 9388 19756 9428
rect 19796 9388 21676 9428
rect 21716 9388 21725 9428
rect 33091 9388 33100 9428
rect 33140 9388 33484 9428
rect 33524 9388 33533 9428
rect 1411 9304 1420 9344
rect 1460 9304 34252 9344
rect 34292 9304 34301 9344
rect 4919 9052 4928 9092
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 5296 9052 5305 9092
rect 20039 9052 20048 9092
rect 20088 9052 20130 9092
rect 20170 9052 20212 9092
rect 20252 9052 20294 9092
rect 20334 9052 20376 9092
rect 20416 9052 20425 9092
rect 35159 9052 35168 9092
rect 35208 9052 35250 9092
rect 35290 9052 35332 9092
rect 35372 9052 35414 9092
rect 35454 9052 35496 9092
rect 35536 9052 35545 9092
rect 1411 8968 1420 9008
rect 1460 8968 37228 9008
rect 37268 8968 37277 9008
rect 39811 8884 39820 8924
rect 39860 8884 40300 8924
rect 40340 8884 40349 8924
rect 20515 8800 20524 8840
rect 20564 8800 26380 8840
rect 26420 8800 26429 8840
rect 1411 8716 1420 8756
rect 1460 8716 35788 8756
rect 35828 8716 35837 8756
rect 547 8632 556 8672
rect 596 8632 37900 8672
rect 37940 8632 37949 8672
rect 3679 8296 3688 8336
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 4056 8296 4065 8336
rect 18799 8296 18808 8336
rect 18848 8296 18890 8336
rect 18930 8296 18972 8336
rect 19012 8296 19054 8336
rect 19094 8296 19136 8336
rect 19176 8296 19185 8336
rect 33919 8296 33928 8336
rect 33968 8296 34010 8336
rect 34050 8296 34092 8336
rect 34132 8296 34174 8336
rect 34214 8296 34256 8336
rect 34296 8296 34305 8336
rect 20131 8044 20140 8084
rect 20180 8044 27532 8084
rect 27572 8044 27581 8084
rect 27235 7960 27244 8000
rect 27284 7960 29260 8000
rect 29300 7960 29309 8000
rect 14947 7876 14956 7916
rect 14996 7876 24652 7916
rect 24692 7876 24701 7916
rect 36163 7876 36172 7916
rect 36212 7876 36940 7916
rect 36980 7876 36989 7916
rect 35203 7792 35212 7832
rect 35252 7792 40300 7832
rect 40340 7792 40349 7832
rect 4771 7624 4780 7664
rect 4820 7624 5548 7664
rect 5588 7624 5597 7664
rect 4919 7540 4928 7580
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 5296 7540 5305 7580
rect 20039 7540 20048 7580
rect 20088 7540 20130 7580
rect 20170 7540 20212 7580
rect 20252 7540 20294 7580
rect 20334 7540 20376 7580
rect 20416 7540 20425 7580
rect 35159 7540 35168 7580
rect 35208 7540 35250 7580
rect 35290 7540 35332 7580
rect 35372 7540 35414 7580
rect 35454 7540 35496 7580
rect 35536 7540 35545 7580
rect 3679 6784 3688 6824
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 4056 6784 4065 6824
rect 18799 6784 18808 6824
rect 18848 6784 18890 6824
rect 18930 6784 18972 6824
rect 19012 6784 19054 6824
rect 19094 6784 19136 6824
rect 19176 6784 19185 6824
rect 33919 6784 33928 6824
rect 33968 6784 34010 6824
rect 34050 6784 34092 6824
rect 34132 6784 34174 6824
rect 34214 6784 34256 6824
rect 34296 6784 34305 6824
rect 16099 6616 16108 6656
rect 16148 6616 23116 6656
rect 23156 6616 23165 6656
rect 18499 6532 18508 6572
rect 18548 6532 27724 6572
rect 27764 6532 27773 6572
rect 18115 6448 18124 6488
rect 18164 6448 27820 6488
rect 27860 6448 27869 6488
rect 4919 6028 4928 6068
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 5296 6028 5305 6068
rect 20039 6028 20048 6068
rect 20088 6028 20130 6068
rect 20170 6028 20212 6068
rect 20252 6028 20294 6068
rect 20334 6028 20376 6068
rect 20416 6028 20425 6068
rect 35159 6028 35168 6068
rect 35208 6028 35250 6068
rect 35290 6028 35332 6068
rect 35372 6028 35414 6068
rect 35454 6028 35496 6068
rect 35536 6028 35545 6068
rect 15427 5776 15436 5816
rect 15476 5776 18604 5816
rect 18644 5776 18653 5816
rect 19843 5608 19852 5648
rect 19892 5608 21772 5648
rect 21812 5608 21821 5648
rect 16963 5524 16972 5564
rect 17012 5524 20428 5564
rect 20468 5524 20477 5564
rect 17155 5440 17164 5480
rect 17204 5440 20716 5480
rect 20756 5440 20765 5480
rect 3679 5272 3688 5312
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 4056 5272 4065 5312
rect 18799 5272 18808 5312
rect 18848 5272 18890 5312
rect 18930 5272 18972 5312
rect 19012 5272 19054 5312
rect 19094 5272 19136 5312
rect 19176 5272 19185 5312
rect 33919 5272 33928 5312
rect 33968 5272 34010 5312
rect 34050 5272 34092 5312
rect 34132 5272 34174 5312
rect 34214 5272 34256 5312
rect 34296 5272 34305 5312
rect 19171 4936 19180 4976
rect 19220 4936 21292 4976
rect 21332 4936 21341 4976
rect 19267 4768 19276 4808
rect 19316 4768 22540 4808
rect 22580 4768 22589 4808
rect 16771 4684 16780 4724
rect 16820 4684 20140 4724
rect 20180 4684 20189 4724
rect 15331 4600 15340 4640
rect 15380 4600 19756 4640
rect 19796 4600 19805 4640
rect 4919 4516 4928 4556
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 5296 4516 5305 4556
rect 20039 4516 20048 4556
rect 20088 4516 20130 4556
rect 20170 4516 20212 4556
rect 20252 4516 20294 4556
rect 20334 4516 20376 4556
rect 20416 4516 20425 4556
rect 35159 4516 35168 4556
rect 35208 4516 35250 4556
rect 35290 4516 35332 4556
rect 35372 4516 35414 4556
rect 35454 4516 35496 4556
rect 35536 4516 35545 4556
rect 20803 4180 20812 4220
rect 20852 4180 23020 4220
rect 23060 4180 23069 4220
rect 31747 4096 31756 4136
rect 31796 4096 40300 4136
rect 40340 4096 40349 4136
rect 21667 4012 21676 4052
rect 21716 4012 25804 4052
rect 25844 4012 25853 4052
rect 20131 3928 20140 3968
rect 20180 3928 26764 3968
rect 26804 3928 26813 3968
rect 3679 3760 3688 3800
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 4056 3760 4065 3800
rect 18799 3760 18808 3800
rect 18848 3760 18890 3800
rect 18930 3760 18972 3800
rect 19012 3760 19054 3800
rect 19094 3760 19136 3800
rect 19176 3760 19185 3800
rect 33919 3760 33928 3800
rect 33968 3760 34010 3800
rect 34050 3760 34092 3800
rect 34132 3760 34174 3800
rect 34214 3760 34256 3800
rect 34296 3760 34305 3800
rect 2179 3340 2188 3380
rect 2228 3340 10060 3380
rect 10100 3340 10109 3380
rect 22915 3340 22924 3380
rect 22964 3340 23500 3380
rect 23540 3340 23549 3380
rect 23395 3172 23404 3212
rect 23444 3172 26284 3212
rect 26324 3172 26333 3212
rect 4919 3004 4928 3044
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 5296 3004 5305 3044
rect 20039 3004 20048 3044
rect 20088 3004 20130 3044
rect 20170 3004 20212 3044
rect 20252 3004 20294 3044
rect 20334 3004 20376 3044
rect 20416 3004 20425 3044
rect 23107 3004 23116 3044
rect 23156 3004 24076 3044
rect 24116 3004 24125 3044
rect 35159 3004 35168 3044
rect 35208 3004 35250 3044
rect 35290 3004 35332 3044
rect 35372 3004 35414 3044
rect 35454 3004 35496 3044
rect 35536 3004 35545 3044
rect 23011 2920 23020 2960
rect 23060 2920 24172 2960
rect 24212 2920 24221 2960
rect 33379 2920 33388 2960
rect 33428 2920 40300 2960
rect 40340 2920 40349 2960
rect 3679 2248 3688 2288
rect 3728 2248 3770 2288
rect 3810 2248 3852 2288
rect 3892 2248 3934 2288
rect 3974 2248 4016 2288
rect 4056 2248 4065 2288
rect 18799 2248 18808 2288
rect 18848 2248 18890 2288
rect 18930 2248 18972 2288
rect 19012 2248 19054 2288
rect 19094 2248 19136 2288
rect 19176 2248 19185 2288
rect 33919 2248 33928 2288
rect 33968 2248 34010 2288
rect 34050 2248 34092 2288
rect 34132 2248 34174 2288
rect 34214 2248 34256 2288
rect 34296 2248 34305 2288
rect 4919 1492 4928 1532
rect 4968 1492 5010 1532
rect 5050 1492 5092 1532
rect 5132 1492 5174 1532
rect 5214 1492 5256 1532
rect 5296 1492 5305 1532
rect 20039 1492 20048 1532
rect 20088 1492 20130 1532
rect 20170 1492 20212 1532
rect 20252 1492 20294 1532
rect 20334 1492 20376 1532
rect 20416 1492 20425 1532
rect 35159 1492 35168 1532
rect 35208 1492 35250 1532
rect 35290 1492 35332 1532
rect 35372 1492 35414 1532
rect 35454 1492 35496 1532
rect 35536 1492 35545 1532
<< via4 >>
rect 3688 9808 3728 9848
rect 3770 9808 3810 9848
rect 3852 9808 3892 9848
rect 3934 9808 3974 9848
rect 4016 9808 4056 9848
rect 18808 9808 18848 9848
rect 18890 9808 18930 9848
rect 18972 9808 19012 9848
rect 19054 9808 19094 9848
rect 19136 9808 19176 9848
rect 33928 9808 33968 9848
rect 34010 9808 34050 9848
rect 34092 9808 34132 9848
rect 34174 9808 34214 9848
rect 34256 9808 34296 9848
rect 4928 9052 4968 9092
rect 5010 9052 5050 9092
rect 5092 9052 5132 9092
rect 5174 9052 5214 9092
rect 5256 9052 5296 9092
rect 20048 9052 20088 9092
rect 20130 9052 20170 9092
rect 20212 9052 20252 9092
rect 20294 9052 20334 9092
rect 20376 9052 20416 9092
rect 35168 9052 35208 9092
rect 35250 9052 35290 9092
rect 35332 9052 35372 9092
rect 35414 9052 35454 9092
rect 35496 9052 35536 9092
rect 3688 8296 3728 8336
rect 3770 8296 3810 8336
rect 3852 8296 3892 8336
rect 3934 8296 3974 8336
rect 4016 8296 4056 8336
rect 18808 8296 18848 8336
rect 18890 8296 18930 8336
rect 18972 8296 19012 8336
rect 19054 8296 19094 8336
rect 19136 8296 19176 8336
rect 33928 8296 33968 8336
rect 34010 8296 34050 8336
rect 34092 8296 34132 8336
rect 34174 8296 34214 8336
rect 34256 8296 34296 8336
rect 4928 7540 4968 7580
rect 5010 7540 5050 7580
rect 5092 7540 5132 7580
rect 5174 7540 5214 7580
rect 5256 7540 5296 7580
rect 20048 7540 20088 7580
rect 20130 7540 20170 7580
rect 20212 7540 20252 7580
rect 20294 7540 20334 7580
rect 20376 7540 20416 7580
rect 35168 7540 35208 7580
rect 35250 7540 35290 7580
rect 35332 7540 35372 7580
rect 35414 7540 35454 7580
rect 35496 7540 35536 7580
rect 3688 6784 3728 6824
rect 3770 6784 3810 6824
rect 3852 6784 3892 6824
rect 3934 6784 3974 6824
rect 4016 6784 4056 6824
rect 18808 6784 18848 6824
rect 18890 6784 18930 6824
rect 18972 6784 19012 6824
rect 19054 6784 19094 6824
rect 19136 6784 19176 6824
rect 33928 6784 33968 6824
rect 34010 6784 34050 6824
rect 34092 6784 34132 6824
rect 34174 6784 34214 6824
rect 34256 6784 34296 6824
rect 4928 6028 4968 6068
rect 5010 6028 5050 6068
rect 5092 6028 5132 6068
rect 5174 6028 5214 6068
rect 5256 6028 5296 6068
rect 20048 6028 20088 6068
rect 20130 6028 20170 6068
rect 20212 6028 20252 6068
rect 20294 6028 20334 6068
rect 20376 6028 20416 6068
rect 35168 6028 35208 6068
rect 35250 6028 35290 6068
rect 35332 6028 35372 6068
rect 35414 6028 35454 6068
rect 35496 6028 35536 6068
rect 3688 5272 3728 5312
rect 3770 5272 3810 5312
rect 3852 5272 3892 5312
rect 3934 5272 3974 5312
rect 4016 5272 4056 5312
rect 18808 5272 18848 5312
rect 18890 5272 18930 5312
rect 18972 5272 19012 5312
rect 19054 5272 19094 5312
rect 19136 5272 19176 5312
rect 33928 5272 33968 5312
rect 34010 5272 34050 5312
rect 34092 5272 34132 5312
rect 34174 5272 34214 5312
rect 34256 5272 34296 5312
rect 4928 4516 4968 4556
rect 5010 4516 5050 4556
rect 5092 4516 5132 4556
rect 5174 4516 5214 4556
rect 5256 4516 5296 4556
rect 20048 4516 20088 4556
rect 20130 4516 20170 4556
rect 20212 4516 20252 4556
rect 20294 4516 20334 4556
rect 20376 4516 20416 4556
rect 35168 4516 35208 4556
rect 35250 4516 35290 4556
rect 35332 4516 35372 4556
rect 35414 4516 35454 4556
rect 35496 4516 35536 4556
rect 3688 3760 3728 3800
rect 3770 3760 3810 3800
rect 3852 3760 3892 3800
rect 3934 3760 3974 3800
rect 4016 3760 4056 3800
rect 18808 3760 18848 3800
rect 18890 3760 18930 3800
rect 18972 3760 19012 3800
rect 19054 3760 19094 3800
rect 19136 3760 19176 3800
rect 33928 3760 33968 3800
rect 34010 3760 34050 3800
rect 34092 3760 34132 3800
rect 34174 3760 34214 3800
rect 34256 3760 34296 3800
rect 4928 3004 4968 3044
rect 5010 3004 5050 3044
rect 5092 3004 5132 3044
rect 5174 3004 5214 3044
rect 5256 3004 5296 3044
rect 20048 3004 20088 3044
rect 20130 3004 20170 3044
rect 20212 3004 20252 3044
rect 20294 3004 20334 3044
rect 20376 3004 20416 3044
rect 35168 3004 35208 3044
rect 35250 3004 35290 3044
rect 35332 3004 35372 3044
rect 35414 3004 35454 3044
rect 35496 3004 35536 3044
rect 3688 2248 3728 2288
rect 3770 2248 3810 2288
rect 3852 2248 3892 2288
rect 3934 2248 3974 2288
rect 4016 2248 4056 2288
rect 18808 2248 18848 2288
rect 18890 2248 18930 2288
rect 18972 2248 19012 2288
rect 19054 2248 19094 2288
rect 19136 2248 19176 2288
rect 33928 2248 33968 2288
rect 34010 2248 34050 2288
rect 34092 2248 34132 2288
rect 34174 2248 34214 2288
rect 34256 2248 34296 2288
rect 4928 1492 4968 1532
rect 5010 1492 5050 1532
rect 5092 1492 5132 1532
rect 5174 1492 5214 1532
rect 5256 1492 5296 1532
rect 20048 1492 20088 1532
rect 20130 1492 20170 1532
rect 20212 1492 20252 1532
rect 20294 1492 20334 1532
rect 20376 1492 20416 1532
rect 35168 1492 35208 1532
rect 35250 1492 35290 1532
rect 35332 1492 35372 1532
rect 35414 1492 35454 1532
rect 35496 1492 35536 1532
<< metal5 >>
rect 3652 9848 4092 11844
rect 3652 9808 3688 9848
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 4056 9808 4092 9848
rect 3652 8336 4092 9808
rect 3652 8296 3688 8336
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 4056 8296 4092 8336
rect 3652 6824 4092 8296
rect 3652 6784 3688 6824
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 4056 6784 4092 6824
rect 3652 5312 4092 6784
rect 3652 5272 3688 5312
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 4056 5272 4092 5312
rect 3652 3800 4092 5272
rect 3652 3760 3688 3800
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 4056 3760 4092 3800
rect 3652 2288 4092 3760
rect 3652 2248 3688 2288
rect 3728 2248 3770 2288
rect 3810 2248 3852 2288
rect 3892 2248 3934 2288
rect 3974 2248 4016 2288
rect 4056 2248 4092 2288
rect 3652 0 4092 2248
rect 4892 9092 5332 11844
rect 4892 9052 4928 9092
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 5296 9052 5332 9092
rect 4892 7580 5332 9052
rect 4892 7540 4928 7580
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 5296 7540 5332 7580
rect 4892 6068 5332 7540
rect 4892 6028 4928 6068
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 5296 6028 5332 6068
rect 4892 4556 5332 6028
rect 4892 4516 4928 4556
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 5296 4516 5332 4556
rect 4892 3044 5332 4516
rect 4892 3004 4928 3044
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 5296 3004 5332 3044
rect 4892 1532 5332 3004
rect 4892 1492 4928 1532
rect 4968 1492 5010 1532
rect 5050 1492 5092 1532
rect 5132 1492 5174 1532
rect 5214 1492 5256 1532
rect 5296 1492 5332 1532
rect 4892 0 5332 1492
rect 18772 9848 19212 11844
rect 18772 9808 18808 9848
rect 18848 9808 18890 9848
rect 18930 9808 18972 9848
rect 19012 9808 19054 9848
rect 19094 9808 19136 9848
rect 19176 9808 19212 9848
rect 18772 8336 19212 9808
rect 18772 8296 18808 8336
rect 18848 8296 18890 8336
rect 18930 8296 18972 8336
rect 19012 8296 19054 8336
rect 19094 8296 19136 8336
rect 19176 8296 19212 8336
rect 18772 6824 19212 8296
rect 18772 6784 18808 6824
rect 18848 6784 18890 6824
rect 18930 6784 18972 6824
rect 19012 6784 19054 6824
rect 19094 6784 19136 6824
rect 19176 6784 19212 6824
rect 18772 5312 19212 6784
rect 18772 5272 18808 5312
rect 18848 5272 18890 5312
rect 18930 5272 18972 5312
rect 19012 5272 19054 5312
rect 19094 5272 19136 5312
rect 19176 5272 19212 5312
rect 18772 3800 19212 5272
rect 18772 3760 18808 3800
rect 18848 3760 18890 3800
rect 18930 3760 18972 3800
rect 19012 3760 19054 3800
rect 19094 3760 19136 3800
rect 19176 3760 19212 3800
rect 18772 2288 19212 3760
rect 18772 2248 18808 2288
rect 18848 2248 18890 2288
rect 18930 2248 18972 2288
rect 19012 2248 19054 2288
rect 19094 2248 19136 2288
rect 19176 2248 19212 2288
rect 18772 0 19212 2248
rect 20012 9092 20452 11844
rect 20012 9052 20048 9092
rect 20088 9052 20130 9092
rect 20170 9052 20212 9092
rect 20252 9052 20294 9092
rect 20334 9052 20376 9092
rect 20416 9052 20452 9092
rect 20012 7580 20452 9052
rect 20012 7540 20048 7580
rect 20088 7540 20130 7580
rect 20170 7540 20212 7580
rect 20252 7540 20294 7580
rect 20334 7540 20376 7580
rect 20416 7540 20452 7580
rect 20012 6068 20452 7540
rect 20012 6028 20048 6068
rect 20088 6028 20130 6068
rect 20170 6028 20212 6068
rect 20252 6028 20294 6068
rect 20334 6028 20376 6068
rect 20416 6028 20452 6068
rect 20012 4556 20452 6028
rect 20012 4516 20048 4556
rect 20088 4516 20130 4556
rect 20170 4516 20212 4556
rect 20252 4516 20294 4556
rect 20334 4516 20376 4556
rect 20416 4516 20452 4556
rect 20012 3044 20452 4516
rect 20012 3004 20048 3044
rect 20088 3004 20130 3044
rect 20170 3004 20212 3044
rect 20252 3004 20294 3044
rect 20334 3004 20376 3044
rect 20416 3004 20452 3044
rect 20012 1532 20452 3004
rect 20012 1492 20048 1532
rect 20088 1492 20130 1532
rect 20170 1492 20212 1532
rect 20252 1492 20294 1532
rect 20334 1492 20376 1532
rect 20416 1492 20452 1532
rect 20012 0 20452 1492
rect 33892 9848 34332 11844
rect 33892 9808 33928 9848
rect 33968 9808 34010 9848
rect 34050 9808 34092 9848
rect 34132 9808 34174 9848
rect 34214 9808 34256 9848
rect 34296 9808 34332 9848
rect 33892 8336 34332 9808
rect 33892 8296 33928 8336
rect 33968 8296 34010 8336
rect 34050 8296 34092 8336
rect 34132 8296 34174 8336
rect 34214 8296 34256 8336
rect 34296 8296 34332 8336
rect 33892 6824 34332 8296
rect 33892 6784 33928 6824
rect 33968 6784 34010 6824
rect 34050 6784 34092 6824
rect 34132 6784 34174 6824
rect 34214 6784 34256 6824
rect 34296 6784 34332 6824
rect 33892 5312 34332 6784
rect 33892 5272 33928 5312
rect 33968 5272 34010 5312
rect 34050 5272 34092 5312
rect 34132 5272 34174 5312
rect 34214 5272 34256 5312
rect 34296 5272 34332 5312
rect 33892 3800 34332 5272
rect 33892 3760 33928 3800
rect 33968 3760 34010 3800
rect 34050 3760 34092 3800
rect 34132 3760 34174 3800
rect 34214 3760 34256 3800
rect 34296 3760 34332 3800
rect 33892 2288 34332 3760
rect 33892 2248 33928 2288
rect 33968 2248 34010 2288
rect 34050 2248 34092 2288
rect 34132 2248 34174 2288
rect 34214 2248 34256 2288
rect 34296 2248 34332 2288
rect 33892 0 34332 2248
rect 35132 9092 35572 11844
rect 35132 9052 35168 9092
rect 35208 9052 35250 9092
rect 35290 9052 35332 9092
rect 35372 9052 35414 9092
rect 35454 9052 35496 9092
rect 35536 9052 35572 9092
rect 35132 7580 35572 9052
rect 35132 7540 35168 7580
rect 35208 7540 35250 7580
rect 35290 7540 35332 7580
rect 35372 7540 35414 7580
rect 35454 7540 35496 7580
rect 35536 7540 35572 7580
rect 35132 6068 35572 7540
rect 35132 6028 35168 6068
rect 35208 6028 35250 6068
rect 35290 6028 35332 6068
rect 35372 6028 35414 6068
rect 35454 6028 35496 6068
rect 35536 6028 35572 6068
rect 35132 4556 35572 6028
rect 35132 4516 35168 4556
rect 35208 4516 35250 4556
rect 35290 4516 35332 4556
rect 35372 4516 35414 4556
rect 35454 4516 35496 4556
rect 35536 4516 35572 4556
rect 35132 3044 35572 4516
rect 35132 3004 35168 3044
rect 35208 3004 35250 3044
rect 35290 3004 35332 3044
rect 35372 3004 35414 3044
rect 35454 3004 35496 3044
rect 35536 3004 35572 3044
rect 35132 1532 35572 3004
rect 35132 1492 35168 1532
rect 35208 1492 35250 1532
rect 35290 1492 35332 1532
rect 35372 1492 35414 1532
rect 35454 1492 35496 1532
rect 35536 1492 35572 1532
rect 35132 0 35572 1492
use sg13g2_buf_1  _001_
timestamp 1676381911
transform 1 0 20928 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _002_
timestamp 1676381911
transform 1 0 21312 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _003_
timestamp 1676381911
transform 1 0 21696 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _004_
timestamp 1676381911
transform 1 0 18912 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _005_
timestamp 1676381911
transform 1 0 24384 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _006_
timestamp 1676381911
transform 1 0 23328 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _007_
timestamp 1676381911
transform 1 0 22560 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _008_
timestamp 1676381911
transform 1 0 24768 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _009_
timestamp 1676381911
transform 1 0 19680 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _010_
timestamp 1676381911
transform 1 0 25824 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _011_
timestamp 1676381911
transform 1 0 26688 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _012_
timestamp 1676381911
transform 1 0 27552 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _013_
timestamp 1676381911
transform 1 0 27072 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _014_
timestamp 1676381911
transform 1 0 24000 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _015_
timestamp 1676381911
transform 1 0 27936 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _016_
timestamp 1676381911
transform 1 0 31776 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _017_
timestamp 1676381911
transform 1 0 34368 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _018_
timestamp 1676381911
transform 1 0 31968 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _019_
timestamp 1676381911
transform 1 0 33696 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _020_
timestamp 1676381911
transform 1 0 33216 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _021_
timestamp 1676381911
transform 1 0 32640 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _022_
timestamp 1676381911
transform 1 0 35616 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _023_
timestamp 1676381911
transform 1 0 31776 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _024_
timestamp 1676381911
transform 1 0 36384 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _025_
timestamp 1676381911
transform 1 0 36000 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _026_
timestamp 1676381911
transform 1 0 37440 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _027_
timestamp 1676381911
transform 1 0 34464 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _028_
timestamp 1676381911
transform 1 0 36384 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _029_
timestamp 1676381911
transform 1 0 33792 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _030_
timestamp 1676381911
transform 1 0 37824 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _031_
timestamp 1676381911
transform -1 0 43488 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _032_
timestamp 1676381911
transform 1 0 39456 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _033_
timestamp 1676381911
transform 1 0 7680 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _034_
timestamp 1676381911
transform 1 0 7296 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _035_
timestamp 1676381911
transform 1 0 8448 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _036_
timestamp 1676381911
transform 1 0 11232 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _037_
timestamp 1676381911
transform 1 0 17952 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _038_
timestamp 1676381911
transform 1 0 25728 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _039_
timestamp 1676381911
transform 1 0 26016 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _040_
timestamp 1676381911
transform 1 0 22944 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _041_
timestamp 1676381911
transform 1 0 23712 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _042_
timestamp 1676381911
transform 1 0 27264 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _043_
timestamp 1676381911
transform 1 0 29760 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _044_
timestamp 1676381911
transform 1 0 29376 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _045_
timestamp 1676381911
transform 1 0 30144 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _046_
timestamp 1676381911
transform 1 0 30528 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _047_
timestamp 1676381911
transform 1 0 31584 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _048_
timestamp 1676381911
transform 1 0 31968 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _049_
timestamp 1676381911
transform 1 0 32352 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _050_
timestamp 1676381911
transform 1 0 32928 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _051_
timestamp 1676381911
transform 1 0 33888 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _052_
timestamp 1676381911
transform 1 0 34560 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _053_
timestamp 1676381911
transform 1 0 8736 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _054_
timestamp 1676381911
transform 1 0 9120 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _055_
timestamp 1676381911
transform 1 0 8352 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _056_
timestamp 1676381911
transform 1 0 8256 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _057_
timestamp 1676381911
transform 1 0 10944 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _058_
timestamp 1676381911
transform -1 0 11712 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _059_
timestamp 1676381911
transform 1 0 11712 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _060_
timestamp 1676381911
transform 1 0 10560 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _061_
timestamp 1676381911
transform 1 0 10176 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _062_
timestamp 1676381911
transform 1 0 9792 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _063_
timestamp 1676381911
transform 1 0 9408 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _064_
timestamp 1676381911
transform 1 0 9792 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _065_
timestamp 1676381911
transform -1 0 13920 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _066_
timestamp 1676381911
transform -1 0 15072 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _067_
timestamp 1676381911
transform -1 0 14688 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _068_
timestamp 1676381911
transform -1 0 15456 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _069_
timestamp 1676381911
transform 1 0 13920 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _070_
timestamp 1676381911
transform -1 0 14304 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _071_
timestamp 1676381911
transform 1 0 13152 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _072_
timestamp 1676381911
transform 1 0 13632 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _073_
timestamp 1676381911
transform -1 0 18240 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _074_
timestamp 1676381911
transform -1 0 18624 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _075_
timestamp 1676381911
transform -1 0 19488 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _076_
timestamp 1676381911
transform -1 0 19680 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _077_
timestamp 1676381911
transform -1 0 21696 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _078_
timestamp 1676381911
transform -1 0 19008 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _079_
timestamp 1676381911
transform -1 0 21312 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _080_
timestamp 1676381911
transform -1 0 20544 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _081_
timestamp 1676381911
transform -1 0 20544 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _082_
timestamp 1676381911
transform -1 0 19392 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _083_
timestamp 1676381911
transform -1 0 20160 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _084_
timestamp 1676381911
transform -1 0 20160 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _085_
timestamp 1676381911
transform -1 0 19776 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _086_
timestamp 1676381911
transform -1 0 20928 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _087_
timestamp 1676381911
transform -1 0 20544 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _088_
timestamp 1676381911
transform -1 0 20160 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _089_
timestamp 1676381911
transform -1 0 27552 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _090_
timestamp 1676381911
transform -1 0 26784 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _091_
timestamp 1676381911
transform -1 0 26208 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _092_
timestamp 1676381911
transform -1 0 26688 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _093_
timestamp 1676381911
transform -1 0 25920 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _094_
timestamp 1676381911
transform -1 0 25536 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _095_
timestamp 1676381911
transform -1 0 26304 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _096_
timestamp 1676381911
transform -1 0 26016 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _097_
timestamp 1676381911
transform -1 0 27072 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _098_
timestamp 1676381911
transform -1 0 27456 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _099_
timestamp 1676381911
transform -1 0 27840 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _100_
timestamp 1676381911
transform -1 0 27936 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _101_
timestamp 1676381911
transform -1 0 28320 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _102_
timestamp 1676381911
transform -1 0 28704 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _103_
timestamp 1676381911
transform -1 0 29088 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _104_
timestamp 1676381911
transform -1 0 28320 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _105_
timestamp 1676381911
transform 1 0 9024 0 -1 6048
box -48 -56 432 834
use sg13g2_antennanp  ANTENNA_1
timestamp 1679999689
transform 1 0 34656 0 1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_2
timestamp 1679999689
transform 1 0 35904 0 1 6048
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_3
timestamp 1679999689
transform 1 0 37632 0 1 7560
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_4
timestamp 1679999689
transform 1 0 40224 0 -1 9072
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_5
timestamp 1679999689
transform -1 0 34464 0 1 7560
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_6
timestamp 1679999689
transform -1 0 38496 0 1 7560
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_7
timestamp 1679999689
transform -1 0 34656 0 1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_8
timestamp 1679999689
transform -1 0 35904 0 1 6048
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_9
timestamp 1679999689
transform 1 0 37920 0 1 7560
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_10
timestamp 1679999689
transform 1 0 39648 0 -1 9072
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_11
timestamp 1679999689
transform -1 0 34752 0 1 7560
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_12
timestamp 1679999689
transform 1 0 40704 0 1 9072
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_13
timestamp 1679999689
transform 1 0 39936 0 -1 9072
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_14
timestamp 1679999689
transform 1 0 37344 0 1 7560
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_15
timestamp 1679999689
transform -1 0 38784 0 1 7560
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_16
timestamp 1679999689
transform -1 0 35040 0 1 7560
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_17
timestamp 1679999689
transform 1 0 40416 0 1 9072
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_18
timestamp 1679999689
transform -1 0 36288 0 -1 7560
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_19
timestamp 1679999689
transform -1 0 40416 0 1 9072
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_20
timestamp 1679999689
transform 1 0 37056 0 1 7560
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_21
timestamp 1679999689
transform 1 0 39840 0 1 9072
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_22
timestamp 1679999689
transform 1 0 39264 0 1 9072
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_23
timestamp 1679999689
transform 1 0 39360 0 -1 9072
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_24
timestamp 1679999689
transform -1 0 37056 0 1 7560
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_25
timestamp 1679999689
transform 1 0 39552 0 1 9072
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_26
timestamp 1679999689
transform -1 0 38976 0 1 9072
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_27
timestamp 1679999689
transform 1 0 39072 0 -1 9072
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_28
timestamp 1679999689
transform -1 0 36192 0 1 7560
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_29
timestamp 1679999689
transform 1 0 38976 0 1 9072
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_30
timestamp 1679999689
transform -1 0 38400 0 1 9072
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_31
timestamp 1679999689
transform 1 0 38784 0 -1 9072
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_32
timestamp 1679999689
transform -1 0 35904 0 1 7560
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_33
timestamp 1679999689
transform 1 0 38400 0 1 9072
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_34
timestamp 1679999689
transform -1 0 37824 0 1 9072
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_35
timestamp 1679999689
transform 1 0 38496 0 -1 9072
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_36
timestamp 1679999689
transform -1 0 35616 0 1 7560
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_37
timestamp 1679999689
transform 1 0 37824 0 1 9072
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_38
timestamp 1679999689
transform -1 0 37248 0 1 9072
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_39
timestamp 1679999689
transform 1 0 38208 0 -1 9072
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_40
timestamp 1679999689
transform -1 0 35328 0 1 7560
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_41
timestamp 1679999689
transform 1 0 37248 0 1 9072
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_42
timestamp 1679999689
transform 1 0 35712 0 -1 9072
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_43
timestamp 1679999689
transform 1 0 37152 0 -1 9072
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_44
timestamp 1679999689
transform 1 0 34176 0 -1 9072
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_45
timestamp 1679999689
transform 1 0 36768 0 -1 9072
box -48 -56 336 834
use sg13g2_decap_8  FILLER_0_0
timestamp 1679581782
transform 1 0 1152 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_7
timestamp 1679581782
transform 1 0 1824 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_14
timestamp 1679581782
transform 1 0 2496 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_21
timestamp 1679581782
transform 1 0 3168 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_28
timestamp 1679581782
transform 1 0 3840 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_35
timestamp 1679581782
transform 1 0 4512 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_42
timestamp 1679581782
transform 1 0 5184 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_49
timestamp 1679581782
transform 1 0 5856 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_56
timestamp 1679581782
transform 1 0 6528 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_63
timestamp 1679581782
transform 1 0 7200 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_70
timestamp 1679581782
transform 1 0 7872 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_77
timestamp 1679581782
transform 1 0 8544 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_84
timestamp 1679581782
transform 1 0 9216 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_91
timestamp 1679581782
transform 1 0 9888 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_98
timestamp 1679581782
transform 1 0 10560 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_105
timestamp 1679581782
transform 1 0 11232 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_112
timestamp 1679581782
transform 1 0 11904 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_119
timestamp 1679581782
transform 1 0 12576 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_126
timestamp 1679581782
transform 1 0 13248 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_133
timestamp 1679581782
transform 1 0 13920 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_140
timestamp 1679581782
transform 1 0 14592 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_147
timestamp 1679581782
transform 1 0 15264 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_154
timestamp 1679581782
transform 1 0 15936 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_161
timestamp 1679581782
transform 1 0 16608 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_168
timestamp 1679581782
transform 1 0 17280 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_175
timestamp 1679581782
transform 1 0 17952 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_182
timestamp 1679581782
transform 1 0 18624 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_189
timestamp 1679581782
transform 1 0 19296 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_196
timestamp 1679581782
transform 1 0 19968 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_203
timestamp 1679581782
transform 1 0 20640 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_210
timestamp 1679581782
transform 1 0 21312 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_217
timestamp 1679581782
transform 1 0 21984 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_224
timestamp 1679581782
transform 1 0 22656 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_231
timestamp 1679581782
transform 1 0 23328 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_238
timestamp 1679581782
transform 1 0 24000 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_245
timestamp 1679581782
transform 1 0 24672 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_252
timestamp 1679581782
transform 1 0 25344 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_259
timestamp 1679581782
transform 1 0 26016 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_266
timestamp 1679581782
transform 1 0 26688 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_273
timestamp 1679581782
transform 1 0 27360 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_280
timestamp 1679581782
transform 1 0 28032 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_287
timestamp 1679581782
transform 1 0 28704 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_294
timestamp 1679581782
transform 1 0 29376 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_301
timestamp 1679581782
transform 1 0 30048 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_308
timestamp 1679581782
transform 1 0 30720 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_315
timestamp 1679581782
transform 1 0 31392 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_322
timestamp 1679581782
transform 1 0 32064 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_329
timestamp 1679581782
transform 1 0 32736 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_336
timestamp 1679581782
transform 1 0 33408 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_343
timestamp 1679581782
transform 1 0 34080 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_350
timestamp 1679581782
transform 1 0 34752 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_357
timestamp 1679581782
transform 1 0 35424 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_364
timestamp 1679581782
transform 1 0 36096 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_371
timestamp 1679581782
transform 1 0 36768 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_378
timestamp 1679581782
transform 1 0 37440 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_385
timestamp 1679581782
transform 1 0 38112 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_392
timestamp 1679581782
transform 1 0 38784 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_399
timestamp 1679581782
transform 1 0 39456 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_406
timestamp 1679581782
transform 1 0 40128 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_413
timestamp 1679581782
transform 1 0 40800 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_420
timestamp 1679581782
transform 1 0 41472 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_427
timestamp 1679581782
transform 1 0 42144 0 1 1512
box -48 -56 720 834
use sg13g2_decap_4  FILLER_0_434
timestamp 1679577901
transform 1 0 42816 0 1 1512
box -48 -56 432 834
use sg13g2_fill_1  FILLER_0_438
timestamp 1677579658
transform 1 0 43200 0 1 1512
box -48 -56 144 834
use sg13g2_decap_8  FILLER_1_0
timestamp 1679581782
transform 1 0 1152 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_7
timestamp 1679581782
transform 1 0 1824 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_14
timestamp 1679581782
transform 1 0 2496 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_21
timestamp 1679581782
transform 1 0 3168 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_28
timestamp 1679581782
transform 1 0 3840 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_35
timestamp 1679581782
transform 1 0 4512 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_42
timestamp 1679581782
transform 1 0 5184 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_49
timestamp 1679581782
transform 1 0 5856 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_56
timestamp 1679581782
transform 1 0 6528 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_63
timestamp 1679581782
transform 1 0 7200 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_70
timestamp 1679581782
transform 1 0 7872 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_77
timestamp 1679581782
transform 1 0 8544 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_84
timestamp 1679581782
transform 1 0 9216 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_91
timestamp 1679581782
transform 1 0 9888 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_98
timestamp 1679581782
transform 1 0 10560 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_109
timestamp 1679581782
transform 1 0 11616 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_116
timestamp 1679581782
transform 1 0 12288 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_123
timestamp 1679581782
transform 1 0 12960 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_130
timestamp 1679581782
transform 1 0 13632 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_137
timestamp 1679581782
transform 1 0 14304 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_144
timestamp 1679581782
transform 1 0 14976 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_151
timestamp 1679581782
transform 1 0 15648 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_158
timestamp 1679581782
transform 1 0 16320 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_165
timestamp 1679581782
transform 1 0 16992 0 -1 3024
box -48 -56 720 834
use sg13g2_fill_2  FILLER_1_172
timestamp 1677580104
transform 1 0 17664 0 -1 3024
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_174
timestamp 1677579658
transform 1 0 17856 0 -1 3024
box -48 -56 144 834
use sg13g2_decap_8  FILLER_1_179
timestamp 1679581782
transform 1 0 18336 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_186
timestamp 1679581782
transform 1 0 19008 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_193
timestamp 1679581782
transform 1 0 19680 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_200
timestamp 1679581782
transform 1 0 20352 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_207
timestamp 1679581782
transform 1 0 21024 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_214
timestamp 1679581782
transform 1 0 21696 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_221
timestamp 1679581782
transform 1 0 22368 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_228
timestamp 1679581782
transform 1 0 23040 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_235
timestamp 1679581782
transform 1 0 23712 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_242
timestamp 1679581782
transform 1 0 24384 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_249
timestamp 1679581782
transform 1 0 25056 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_256
timestamp 1679581782
transform 1 0 25728 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_263
timestamp 1679581782
transform 1 0 26400 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_4  FILLER_1_274
timestamp 1679577901
transform 1 0 27456 0 -1 3024
box -48 -56 432 834
use sg13g2_fill_1  FILLER_1_278
timestamp 1677579658
transform 1 0 27840 0 -1 3024
box -48 -56 144 834
use sg13g2_decap_8  FILLER_1_283
timestamp 1679581782
transform 1 0 28320 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_290
timestamp 1679581782
transform 1 0 28992 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_297
timestamp 1679581782
transform 1 0 29664 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_304
timestamp 1679581782
transform 1 0 30336 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_311
timestamp 1679581782
transform 1 0 31008 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_318
timestamp 1679581782
transform 1 0 31680 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_325
timestamp 1679581782
transform 1 0 32352 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_332
timestamp 1679581782
transform 1 0 33024 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_339
timestamp 1679581782
transform 1 0 33696 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_346
timestamp 1679581782
transform 1 0 34368 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_353
timestamp 1679581782
transform 1 0 35040 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_360
timestamp 1679581782
transform 1 0 35712 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_367
timestamp 1679581782
transform 1 0 36384 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_374
timestamp 1679581782
transform 1 0 37056 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_381
timestamp 1679581782
transform 1 0 37728 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_388
timestamp 1679581782
transform 1 0 38400 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_395
timestamp 1679581782
transform 1 0 39072 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_402
timestamp 1679581782
transform 1 0 39744 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_409
timestamp 1679581782
transform 1 0 40416 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_416
timestamp 1679581782
transform 1 0 41088 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_423
timestamp 1679581782
transform 1 0 41760 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_430
timestamp 1679581782
transform 1 0 42432 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_437
timestamp 1679581782
transform 1 0 43104 0 -1 3024
box -48 -56 720 834
use sg13g2_fill_2  FILLER_1_444
timestamp 1677580104
transform 1 0 43776 0 -1 3024
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_446
timestamp 1677579658
transform 1 0 43968 0 -1 3024
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_0
timestamp 1679581782
transform 1 0 1152 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_7
timestamp 1679581782
transform 1 0 1824 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_14
timestamp 1679581782
transform 1 0 2496 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_21
timestamp 1679581782
transform 1 0 3168 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_28
timestamp 1679581782
transform 1 0 3840 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_35
timestamp 1679581782
transform 1 0 4512 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_42
timestamp 1679581782
transform 1 0 5184 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_49
timestamp 1679581782
transform 1 0 5856 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_56
timestamp 1679581782
transform 1 0 6528 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_63
timestamp 1679581782
transform 1 0 7200 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_70
timestamp 1679581782
transform 1 0 7872 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_77
timestamp 1679581782
transform 1 0 8544 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_84
timestamp 1679581782
transform 1 0 9216 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_91
timestamp 1679581782
transform 1 0 9888 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_98
timestamp 1679581782
transform 1 0 10560 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_105
timestamp 1679581782
transform 1 0 11232 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_112
timestamp 1679581782
transform 1 0 11904 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_119
timestamp 1679581782
transform 1 0 12576 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_126
timestamp 1679581782
transform 1 0 13248 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_133
timestamp 1679581782
transform 1 0 13920 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_140
timestamp 1679581782
transform 1 0 14592 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_147
timestamp 1679581782
transform 1 0 15264 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_154
timestamp 1679581782
transform 1 0 15936 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_161
timestamp 1679581782
transform 1 0 16608 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_168
timestamp 1679581782
transform 1 0 17280 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_175
timestamp 1679581782
transform 1 0 17952 0 1 3024
box -48 -56 720 834
use sg13g2_fill_2  FILLER_2_182
timestamp 1677580104
transform 1 0 18624 0 1 3024
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_184
timestamp 1677579658
transform 1 0 18816 0 1 3024
box -48 -56 144 834
use sg13g2_decap_4  FILLER_2_189
timestamp 1679577901
transform 1 0 19296 0 1 3024
box -48 -56 432 834
use sg13g2_decap_8  FILLER_2_197
timestamp 1679581782
transform 1 0 20064 0 1 3024
box -48 -56 720 834
use sg13g2_fill_2  FILLER_2_204
timestamp 1677580104
transform 1 0 20736 0 1 3024
box -48 -56 240 834
use sg13g2_decap_4  FILLER_2_218
timestamp 1679577901
transform 1 0 22080 0 1 3024
box -48 -56 432 834
use sg13g2_fill_1  FILLER_2_222
timestamp 1677579658
transform 1 0 22464 0 1 3024
box -48 -56 144 834
use sg13g2_fill_2  FILLER_2_235
timestamp 1677580104
transform 1 0 23712 0 1 3024
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_237
timestamp 1677579658
transform 1 0 23904 0 1 3024
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_250
timestamp 1679581782
transform 1 0 25152 0 1 3024
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_261
timestamp 1679577901
transform 1 0 26208 0 1 3024
box -48 -56 432 834
use sg13g2_fill_1  FILLER_2_265
timestamp 1677579658
transform 1 0 26592 0 1 3024
box -48 -56 144 834
use sg13g2_decap_4  FILLER_2_270
timestamp 1679577901
transform 1 0 27072 0 1 3024
box -48 -56 432 834
use sg13g2_fill_1  FILLER_2_274
timestamp 1677579658
transform 1 0 27456 0 1 3024
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_279
timestamp 1679581782
transform 1 0 27936 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_286
timestamp 1679581782
transform 1 0 28608 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_293
timestamp 1679581782
transform 1 0 29280 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_300
timestamp 1679581782
transform 1 0 29952 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_307
timestamp 1679581782
transform 1 0 30624 0 1 3024
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_314
timestamp 1679577901
transform 1 0 31296 0 1 3024
box -48 -56 432 834
use sg13g2_fill_1  FILLER_2_318
timestamp 1677579658
transform 1 0 31680 0 1 3024
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_323
timestamp 1679581782
transform 1 0 32160 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_330
timestamp 1679581782
transform 1 0 32832 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_337
timestamp 1679581782
transform 1 0 33504 0 1 3024
box -48 -56 720 834
use sg13g2_fill_2  FILLER_2_344
timestamp 1677580104
transform 1 0 34176 0 1 3024
box -48 -56 240 834
use sg13g2_decap_8  FILLER_2_352
timestamp 1679581782
transform 1 0 34944 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_359
timestamp 1679581782
transform 1 0 35616 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_366
timestamp 1679581782
transform 1 0 36288 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_373
timestamp 1679581782
transform 1 0 36960 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_380
timestamp 1679581782
transform 1 0 37632 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_387
timestamp 1679581782
transform 1 0 38304 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_394
timestamp 1679581782
transform 1 0 38976 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_401
timestamp 1679581782
transform 1 0 39648 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_408
timestamp 1679581782
transform 1 0 40320 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_415
timestamp 1679581782
transform 1 0 40992 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_422
timestamp 1679581782
transform 1 0 41664 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_429
timestamp 1679581782
transform 1 0 42336 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_436
timestamp 1679581782
transform 1 0 43008 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_443
timestamp 1679581782
transform 1 0 43680 0 1 3024
box -48 -56 720 834
use sg13g2_fill_1  FILLER_2_450
timestamp 1677579658
transform 1 0 44352 0 1 3024
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_0
timestamp 1679581782
transform 1 0 1152 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_7
timestamp 1679581782
transform 1 0 1824 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_14
timestamp 1679581782
transform 1 0 2496 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_21
timestamp 1679581782
transform 1 0 3168 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_28
timestamp 1679581782
transform 1 0 3840 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_35
timestamp 1679581782
transform 1 0 4512 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_42
timestamp 1679581782
transform 1 0 5184 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_49
timestamp 1679581782
transform 1 0 5856 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_56
timestamp 1679581782
transform 1 0 6528 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_63
timestamp 1679581782
transform 1 0 7200 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_70
timestamp 1679581782
transform 1 0 7872 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_77
timestamp 1679581782
transform 1 0 8544 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_84
timestamp 1679581782
transform 1 0 9216 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_91
timestamp 1679581782
transform 1 0 9888 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_98
timestamp 1679581782
transform 1 0 10560 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_105
timestamp 1679581782
transform 1 0 11232 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_112
timestamp 1679581782
transform 1 0 11904 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_119
timestamp 1679581782
transform 1 0 12576 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_126
timestamp 1679581782
transform 1 0 13248 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_133
timestamp 1679581782
transform 1 0 13920 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_140
timestamp 1679581782
transform 1 0 14592 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_147
timestamp 1679581782
transform 1 0 15264 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_154
timestamp 1679581782
transform 1 0 15936 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_161
timestamp 1679581782
transform 1 0 16608 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_168
timestamp 1679581782
transform 1 0 17280 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_175
timestamp 1679581782
transform 1 0 17952 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_182
timestamp 1679581782
transform 1 0 18624 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_189
timestamp 1679581782
transform 1 0 19296 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_196
timestamp 1679581782
transform 1 0 19968 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_203
timestamp 1679581782
transform 1 0 20640 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_210
timestamp 1679581782
transform 1 0 21312 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_217
timestamp 1679581782
transform 1 0 21984 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_224
timestamp 1679581782
transform 1 0 22656 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_231
timestamp 1679577901
transform 1 0 23328 0 -1 4536
box -48 -56 432 834
use sg13g2_decap_8  FILLER_3_239
timestamp 1679581782
transform 1 0 24096 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_246
timestamp 1679581782
transform 1 0 24768 0 -1 4536
box -48 -56 720 834
use sg13g2_fill_2  FILLER_3_253
timestamp 1677580104
transform 1 0 25440 0 -1 4536
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_255
timestamp 1677579658
transform 1 0 25632 0 -1 4536
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_260
timestamp 1679581782
transform 1 0 26112 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_267
timestamp 1679581782
transform 1 0 26784 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_274
timestamp 1679581782
transform 1 0 27456 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_281
timestamp 1679581782
transform 1 0 28128 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_288
timestamp 1679581782
transform 1 0 28800 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_295
timestamp 1679581782
transform 1 0 29472 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_302
timestamp 1679581782
transform 1 0 30144 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_309
timestamp 1679581782
transform 1 0 30816 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_316
timestamp 1679581782
transform 1 0 31488 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_323
timestamp 1679581782
transform 1 0 32160 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_330
timestamp 1679581782
transform 1 0 32832 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_337
timestamp 1679581782
transform 1 0 33504 0 -1 4536
box -48 -56 720 834
use sg13g2_fill_2  FILLER_3_344
timestamp 1677580104
transform 1 0 34176 0 -1 4536
box -48 -56 240 834
use sg13g2_decap_8  FILLER_3_350
timestamp 1679581782
transform 1 0 34752 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_357
timestamp 1679581782
transform 1 0 35424 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_364
timestamp 1679581782
transform 1 0 36096 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_371
timestamp 1679581782
transform 1 0 36768 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_378
timestamp 1679581782
transform 1 0 37440 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_385
timestamp 1679581782
transform 1 0 38112 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_392
timestamp 1679581782
transform 1 0 38784 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_399
timestamp 1679581782
transform 1 0 39456 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_406
timestamp 1679581782
transform 1 0 40128 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_413
timestamp 1679581782
transform 1 0 40800 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_420
timestamp 1679581782
transform 1 0 41472 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_427
timestamp 1679581782
transform 1 0 42144 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_434
timestamp 1679581782
transform 1 0 42816 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_441
timestamp 1679581782
transform 1 0 43488 0 -1 4536
box -48 -56 720 834
use sg13g2_fill_2  FILLER_3_448
timestamp 1677580104
transform 1 0 44160 0 -1 4536
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_450
timestamp 1677579658
transform 1 0 44352 0 -1 4536
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_0
timestamp 1679581782
transform 1 0 1152 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_7
timestamp 1679581782
transform 1 0 1824 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_14
timestamp 1679581782
transform 1 0 2496 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_21
timestamp 1679581782
transform 1 0 3168 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_28
timestamp 1679581782
transform 1 0 3840 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_35
timestamp 1679581782
transform 1 0 4512 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_42
timestamp 1679581782
transform 1 0 5184 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_49
timestamp 1679581782
transform 1 0 5856 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_56
timestamp 1679581782
transform 1 0 6528 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_63
timestamp 1679581782
transform 1 0 7200 0 1 4536
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_70
timestamp 1679577901
transform 1 0 7872 0 1 4536
box -48 -56 432 834
use sg13g2_fill_2  FILLER_4_74
timestamp 1677580104
transform 1 0 8256 0 1 4536
box -48 -56 240 834
use sg13g2_decap_8  FILLER_4_80
timestamp 1679581782
transform 1 0 8832 0 1 4536
box -48 -56 720 834
use sg13g2_fill_2  FILLER_4_87
timestamp 1677580104
transform 1 0 9504 0 1 4536
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_89
timestamp 1677579658
transform 1 0 9696 0 1 4536
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_94
timestamp 1679581782
transform 1 0 10176 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_101
timestamp 1679581782
transform 1 0 10848 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_108
timestamp 1679581782
transform 1 0 11520 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_115
timestamp 1679581782
transform 1 0 12192 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_122
timestamp 1679581782
transform 1 0 12864 0 1 4536
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_129
timestamp 1679577901
transform 1 0 13536 0 1 4536
box -48 -56 432 834
use sg13g2_decap_8  FILLER_4_137
timestamp 1679581782
transform 1 0 14304 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_144
timestamp 1679581782
transform 1 0 14976 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_151
timestamp 1679581782
transform 1 0 15648 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_158
timestamp 1679581782
transform 1 0 16320 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_165
timestamp 1679581782
transform 1 0 16992 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_172
timestamp 1679581782
transform 1 0 17664 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_179
timestamp 1679581782
transform 1 0 18336 0 1 4536
box -48 -56 720 834
use sg13g2_fill_2  FILLER_4_186
timestamp 1677580104
transform 1 0 19008 0 1 4536
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_188
timestamp 1677579658
transform 1 0 19200 0 1 4536
box -48 -56 144 834
use sg13g2_fill_1  FILLER_4_193
timestamp 1677579658
transform 1 0 19680 0 1 4536
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_202
timestamp 1679581782
transform 1 0 20544 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_209
timestamp 1679581782
transform 1 0 21216 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_216
timestamp 1679581782
transform 1 0 21888 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_223
timestamp 1679581782
transform 1 0 22560 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_230
timestamp 1679581782
transform 1 0 23232 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_237
timestamp 1679581782
transform 1 0 23904 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_244
timestamp 1679581782
transform 1 0 24576 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_251
timestamp 1679581782
transform 1 0 25248 0 1 4536
box -48 -56 720 834
use sg13g2_fill_1  FILLER_4_258
timestamp 1677579658
transform 1 0 25920 0 1 4536
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_263
timestamp 1679581782
transform 1 0 26400 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_270
timestamp 1679581782
transform 1 0 27072 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_277
timestamp 1679581782
transform 1 0 27744 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_284
timestamp 1679581782
transform 1 0 28416 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_291
timestamp 1679581782
transform 1 0 29088 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_298
timestamp 1679581782
transform 1 0 29760 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_305
timestamp 1679581782
transform 1 0 30432 0 1 4536
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_312
timestamp 1679577901
transform 1 0 31104 0 1 4536
box -48 -56 432 834
use sg13g2_fill_1  FILLER_4_316
timestamp 1677579658
transform 1 0 31488 0 1 4536
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_325
timestamp 1679581782
transform 1 0 32352 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_332
timestamp 1679581782
transform 1 0 33024 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_339
timestamp 1679581782
transform 1 0 33696 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_346
timestamp 1679581782
transform 1 0 34368 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_353
timestamp 1679581782
transform 1 0 35040 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_360
timestamp 1679581782
transform 1 0 35712 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_367
timestamp 1679581782
transform 1 0 36384 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_374
timestamp 1679581782
transform 1 0 37056 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_381
timestamp 1679581782
transform 1 0 37728 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_388
timestamp 1679581782
transform 1 0 38400 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_395
timestamp 1679581782
transform 1 0 39072 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_402
timestamp 1679581782
transform 1 0 39744 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_409
timestamp 1679581782
transform 1 0 40416 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_416
timestamp 1679581782
transform 1 0 41088 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_423
timestamp 1679581782
transform 1 0 41760 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_430
timestamp 1679581782
transform 1 0 42432 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_437
timestamp 1679581782
transform 1 0 43104 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_444
timestamp 1679581782
transform 1 0 43776 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_0
timestamp 1679581782
transform 1 0 1152 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_7
timestamp 1679581782
transform 1 0 1824 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_14
timestamp 1679581782
transform 1 0 2496 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_21
timestamp 1679581782
transform 1 0 3168 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_28
timestamp 1679581782
transform 1 0 3840 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_35
timestamp 1679581782
transform 1 0 4512 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_42
timestamp 1679581782
transform 1 0 5184 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_49
timestamp 1679581782
transform 1 0 5856 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_56
timestamp 1679581782
transform 1 0 6528 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_63
timestamp 1679581782
transform 1 0 7200 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_70
timestamp 1679581782
transform 1 0 7872 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_77
timestamp 1679577901
transform 1 0 8544 0 -1 6048
box -48 -56 432 834
use sg13g2_fill_1  FILLER_5_81
timestamp 1677579658
transform 1 0 8928 0 -1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_114
timestamp 1679581782
transform 1 0 12096 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_121
timestamp 1679577901
transform 1 0 12768 0 -1 6048
box -48 -56 432 834
use sg13g2_decap_8  FILLER_5_149
timestamp 1679581782
transform 1 0 15456 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_156
timestamp 1679581782
transform 1 0 16128 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_163
timestamp 1679581782
transform 1 0 16800 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_170
timestamp 1679577901
transform 1 0 17472 0 -1 6048
box -48 -56 432 834
use sg13g2_decap_8  FILLER_5_214
timestamp 1679581782
transform 1 0 21696 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_221
timestamp 1679581782
transform 1 0 22368 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_228
timestamp 1679581782
transform 1 0 23040 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_235
timestamp 1679581782
transform 1 0 23712 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_242
timestamp 1679581782
transform 1 0 24384 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_249
timestamp 1679581782
transform 1 0 25056 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_256
timestamp 1679581782
transform 1 0 25728 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_263
timestamp 1679581782
transform 1 0 26400 0 -1 6048
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_270
timestamp 1677580104
transform 1 0 27072 0 -1 6048
box -48 -56 240 834
use sg13g2_decap_8  FILLER_5_276
timestamp 1679581782
transform 1 0 27648 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_283
timestamp 1679581782
transform 1 0 28320 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_290
timestamp 1679577901
transform 1 0 28992 0 -1 6048
box -48 -56 432 834
use sg13g2_decap_8  FILLER_5_310
timestamp 1679581782
transform 1 0 30912 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_317
timestamp 1679577901
transform 1 0 31584 0 -1 6048
box -48 -56 432 834
use sg13g2_fill_2  FILLER_5_329
timestamp 1677580104
transform 1 0 32736 0 -1 6048
box -48 -56 240 834
use sg13g2_decap_4  FILLER_5_335
timestamp 1679577901
transform 1 0 33312 0 -1 6048
box -48 -56 432 834
use sg13g2_fill_2  FILLER_5_339
timestamp 1677580104
transform 1 0 33696 0 -1 6048
box -48 -56 240 834
use sg13g2_fill_2  FILLER_5_345
timestamp 1677580104
transform 1 0 34272 0 -1 6048
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_347
timestamp 1677579658
transform 1 0 34464 0 -1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_352
timestamp 1679581782
transform 1 0 34944 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_359
timestamp 1679581782
transform 1 0 35616 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_366
timestamp 1679581782
transform 1 0 36288 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_373
timestamp 1679581782
transform 1 0 36960 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_380
timestamp 1679581782
transform 1 0 37632 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_387
timestamp 1679581782
transform 1 0 38304 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_394
timestamp 1679581782
transform 1 0 38976 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_401
timestamp 1679581782
transform 1 0 39648 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_408
timestamp 1679581782
transform 1 0 40320 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_415
timestamp 1679581782
transform 1 0 40992 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_422
timestamp 1679581782
transform 1 0 41664 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_429
timestamp 1679581782
transform 1 0 42336 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_436
timestamp 1679581782
transform 1 0 43008 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_443
timestamp 1679581782
transform 1 0 43680 0 -1 6048
box -48 -56 720 834
use sg13g2_fill_1  FILLER_5_450
timestamp 1677579658
transform 1 0 44352 0 -1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_0
timestamp 1679581782
transform 1 0 1152 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_7
timestamp 1679581782
transform 1 0 1824 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_14
timestamp 1679581782
transform 1 0 2496 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_21
timestamp 1679581782
transform 1 0 3168 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_28
timestamp 1679581782
transform 1 0 3840 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_35
timestamp 1679581782
transform 1 0 4512 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_42
timestamp 1679581782
transform 1 0 5184 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_49
timestamp 1679581782
transform 1 0 5856 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_56
timestamp 1679581782
transform 1 0 6528 0 1 6048
box -48 -56 720 834
use sg13g2_fill_1  FILLER_6_63
timestamp 1677579658
transform 1 0 7200 0 1 6048
box -48 -56 144 834
use sg13g2_fill_2  FILLER_6_72
timestamp 1677580104
transform 1 0 8064 0 1 6048
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_74
timestamp 1677579658
transform 1 0 8256 0 1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_87
timestamp 1679581782
transform 1 0 9504 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_94
timestamp 1679581782
transform 1 0 10176 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_101
timestamp 1679581782
transform 1 0 10848 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_108
timestamp 1679581782
transform 1 0 11520 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_115
timestamp 1679581782
transform 1 0 12192 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_122
timestamp 1679581782
transform 1 0 12864 0 1 6048
box -48 -56 720 834
use sg13g2_fill_1  FILLER_6_129
timestamp 1677579658
transform 1 0 13536 0 1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_134
timestamp 1679581782
transform 1 0 14016 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_141
timestamp 1679581782
transform 1 0 14688 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_148
timestamp 1679581782
transform 1 0 15360 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_155
timestamp 1679581782
transform 1 0 16032 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_162
timestamp 1679581782
transform 1 0 16704 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_169
timestamp 1679581782
transform 1 0 17376 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_176
timestamp 1679581782
transform 1 0 18048 0 1 6048
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_183
timestamp 1679577901
transform 1 0 18720 0 1 6048
box -48 -56 432 834
use sg13g2_fill_2  FILLER_6_191
timestamp 1677580104
transform 1 0 19488 0 1 6048
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_193
timestamp 1677579658
transform 1 0 19680 0 1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_202
timestamp 1679581782
transform 1 0 20544 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_209
timestamp 1679581782
transform 1 0 21216 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_216
timestamp 1679581782
transform 1 0 21888 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_223
timestamp 1679581782
transform 1 0 22560 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_230
timestamp 1679581782
transform 1 0 23232 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_237
timestamp 1679581782
transform 1 0 23904 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_244
timestamp 1679581782
transform 1 0 24576 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_251
timestamp 1679581782
transform 1 0 25248 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_258
timestamp 1679581782
transform 1 0 25920 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_265
timestamp 1679581782
transform 1 0 26592 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_272
timestamp 1679581782
transform 1 0 27264 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_279
timestamp 1679581782
transform 1 0 27936 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_286
timestamp 1679581782
transform 1 0 28608 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_293
timestamp 1679581782
transform 1 0 29280 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_300
timestamp 1679581782
transform 1 0 29952 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_307
timestamp 1679581782
transform 1 0 30624 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_314
timestamp 1679581782
transform 1 0 31296 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_321
timestamp 1679581782
transform 1 0 31968 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_328
timestamp 1679581782
transform 1 0 32640 0 1 6048
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_335
timestamp 1679577901
transform 1 0 33312 0 1 6048
box -48 -56 432 834
use sg13g2_decap_8  FILLER_6_343
timestamp 1679581782
transform 1 0 34080 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_350
timestamp 1679581782
transform 1 0 34752 0 1 6048
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_357
timestamp 1677580104
transform 1 0 35424 0 1 6048
box -48 -56 240 834
use sg13g2_decap_8  FILLER_6_365
timestamp 1679581782
transform 1 0 36192 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_372
timestamp 1679581782
transform 1 0 36864 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_379
timestamp 1679581782
transform 1 0 37536 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_386
timestamp 1679581782
transform 1 0 38208 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_393
timestamp 1679581782
transform 1 0 38880 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_400
timestamp 1679581782
transform 1 0 39552 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_407
timestamp 1679581782
transform 1 0 40224 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_414
timestamp 1679581782
transform 1 0 40896 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_421
timestamp 1679581782
transform 1 0 41568 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_428
timestamp 1679581782
transform 1 0 42240 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_435
timestamp 1679581782
transform 1 0 42912 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_442
timestamp 1679581782
transform 1 0 43584 0 1 6048
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_449
timestamp 1677580104
transform 1 0 44256 0 1 6048
box -48 -56 240 834
use sg13g2_decap_8  FILLER_7_0
timestamp 1679581782
transform 1 0 1152 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_7
timestamp 1679581782
transform 1 0 1824 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_14
timestamp 1679581782
transform 1 0 2496 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_21
timestamp 1679581782
transform 1 0 3168 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_28
timestamp 1679581782
transform 1 0 3840 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_35
timestamp 1679581782
transform 1 0 4512 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_42
timestamp 1679581782
transform 1 0 5184 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_49
timestamp 1679581782
transform 1 0 5856 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_56
timestamp 1679581782
transform 1 0 6528 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_63
timestamp 1679581782
transform 1 0 7200 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_4  FILLER_7_70
timestamp 1679577901
transform 1 0 7872 0 -1 7560
box -48 -56 432 834
use sg13g2_decap_8  FILLER_7_78
timestamp 1679581782
transform 1 0 8640 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_85
timestamp 1679581782
transform 1 0 9312 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_92
timestamp 1679581782
transform 1 0 9984 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_99
timestamp 1679581782
transform 1 0 10656 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_106
timestamp 1679581782
transform 1 0 11328 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_113
timestamp 1679581782
transform 1 0 12000 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_120
timestamp 1679581782
transform 1 0 12672 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_127
timestamp 1679581782
transform 1 0 13344 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_134
timestamp 1679581782
transform 1 0 14016 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_141
timestamp 1679581782
transform 1 0 14688 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_148
timestamp 1679581782
transform 1 0 15360 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_155
timestamp 1679581782
transform 1 0 16032 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_162
timestamp 1679581782
transform 1 0 16704 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_169
timestamp 1679581782
transform 1 0 17376 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_176
timestamp 1679581782
transform 1 0 18048 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_183
timestamp 1679581782
transform 1 0 18720 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_190
timestamp 1679581782
transform 1 0 19392 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_197
timestamp 1679581782
transform 1 0 20064 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_204
timestamp 1679581782
transform 1 0 20736 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_211
timestamp 1679581782
transform 1 0 21408 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_218
timestamp 1679581782
transform 1 0 22080 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_225
timestamp 1679581782
transform 1 0 22752 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_232
timestamp 1679581782
transform 1 0 23424 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_239
timestamp 1679581782
transform 1 0 24096 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_246
timestamp 1679581782
transform 1 0 24768 0 -1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_7_253
timestamp 1677580104
transform 1 0 25440 0 -1 7560
box -48 -56 240 834
use sg13g2_decap_8  FILLER_7_259
timestamp 1679581782
transform 1 0 26016 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_266
timestamp 1679581782
transform 1 0 26688 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_273
timestamp 1679581782
transform 1 0 27360 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_280
timestamp 1679581782
transform 1 0 28032 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_287
timestamp 1679581782
transform 1 0 28704 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_294
timestamp 1679581782
transform 1 0 29376 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_301
timestamp 1679581782
transform 1 0 30048 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_308
timestamp 1679581782
transform 1 0 30720 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_315
timestamp 1679581782
transform 1 0 31392 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_322
timestamp 1679581782
transform 1 0 32064 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_4  FILLER_7_329
timestamp 1679577901
transform 1 0 32736 0 -1 7560
box -48 -56 432 834
use sg13g2_fill_1  FILLER_7_333
timestamp 1677579658
transform 1 0 33120 0 -1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_338
timestamp 1679581782
transform 1 0 33600 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_345
timestamp 1679581782
transform 1 0 34272 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_352
timestamp 1679581782
transform 1 0 34944 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_366
timestamp 1679581782
transform 1 0 36288 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_373
timestamp 1679581782
transform 1 0 36960 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_380
timestamp 1679581782
transform 1 0 37632 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_387
timestamp 1679581782
transform 1 0 38304 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_394
timestamp 1679581782
transform 1 0 38976 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_401
timestamp 1679581782
transform 1 0 39648 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_408
timestamp 1679581782
transform 1 0 40320 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_415
timestamp 1679581782
transform 1 0 40992 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_422
timestamp 1679581782
transform 1 0 41664 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_429
timestamp 1679581782
transform 1 0 42336 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_436
timestamp 1679581782
transform 1 0 43008 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_443
timestamp 1679581782
transform 1 0 43680 0 -1 7560
box -48 -56 720 834
use sg13g2_fill_1  FILLER_7_450
timestamp 1677579658
transform 1 0 44352 0 -1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_0
timestamp 1679581782
transform 1 0 1152 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_7
timestamp 1679581782
transform 1 0 1824 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_14
timestamp 1679581782
transform 1 0 2496 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_21
timestamp 1679581782
transform 1 0 3168 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_28
timestamp 1679581782
transform 1 0 3840 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_35
timestamp 1679581782
transform 1 0 4512 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_42
timestamp 1679581782
transform 1 0 5184 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_49
timestamp 1679581782
transform 1 0 5856 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_56
timestamp 1679581782
transform 1 0 6528 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_63
timestamp 1679581782
transform 1 0 7200 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_70
timestamp 1679581782
transform 1 0 7872 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_77
timestamp 1679581782
transform 1 0 8544 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_84
timestamp 1679581782
transform 1 0 9216 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_91
timestamp 1679581782
transform 1 0 9888 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_98
timestamp 1679581782
transform 1 0 10560 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_105
timestamp 1679581782
transform 1 0 11232 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_112
timestamp 1679581782
transform 1 0 11904 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_119
timestamp 1679581782
transform 1 0 12576 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_126
timestamp 1679581782
transform 1 0 13248 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_133
timestamp 1679581782
transform 1 0 13920 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_140
timestamp 1679581782
transform 1 0 14592 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_147
timestamp 1679581782
transform 1 0 15264 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_154
timestamp 1679581782
transform 1 0 15936 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_161
timestamp 1679581782
transform 1 0 16608 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_168
timestamp 1679581782
transform 1 0 17280 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_175
timestamp 1679581782
transform 1 0 17952 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_182
timestamp 1679581782
transform 1 0 18624 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_189
timestamp 1679581782
transform 1 0 19296 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_196
timestamp 1679581782
transform 1 0 19968 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_203
timestamp 1679581782
transform 1 0 20640 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_210
timestamp 1679581782
transform 1 0 21312 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_217
timestamp 1679581782
transform 1 0 21984 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_224
timestamp 1679581782
transform 1 0 22656 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_231
timestamp 1679581782
transform 1 0 23328 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_238
timestamp 1679581782
transform 1 0 24000 0 1 7560
box -48 -56 720 834
use sg13g2_decap_4  FILLER_8_245
timestamp 1679577901
transform 1 0 24672 0 1 7560
box -48 -56 432 834
use sg13g2_fill_1  FILLER_8_249
timestamp 1677579658
transform 1 0 25056 0 1 7560
box -48 -56 144 834
use sg13g2_fill_1  FILLER_8_278
timestamp 1677579658
transform 1 0 27840 0 1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_283
timestamp 1679581782
transform 1 0 28320 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_290
timestamp 1679581782
transform 1 0 28992 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_297
timestamp 1679581782
transform 1 0 29664 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_304
timestamp 1679581782
transform 1 0 30336 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_311
timestamp 1679581782
transform 1 0 31008 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_318
timestamp 1679581782
transform 1 0 31680 0 1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_8_325
timestamp 1677580104
transform 1 0 32352 0 1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_327
timestamp 1677579658
transform 1 0 32544 0 1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_332
timestamp 1679581782
transform 1 0 33024 0 1 7560
box -48 -56 720 834
use sg13g2_decap_4  FILLER_8_339
timestamp 1679577901
transform 1 0 33696 0 1 7560
box -48 -56 432 834
use sg13g2_fill_1  FILLER_8_343
timestamp 1677579658
transform 1 0 34080 0 1 7560
box -48 -56 144 834
use sg13g2_fill_2  FILLER_8_365
timestamp 1677580104
transform 1 0 36192 0 1 7560
box -48 -56 240 834
use sg13g2_decap_8  FILLER_8_392
timestamp 1679581782
transform 1 0 38784 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_403
timestamp 1679581782
transform 1 0 39840 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_410
timestamp 1679581782
transform 1 0 40512 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_417
timestamp 1679581782
transform 1 0 41184 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_424
timestamp 1679581782
transform 1 0 41856 0 1 7560
box -48 -56 720 834
use sg13g2_decap_4  FILLER_8_431
timestamp 1679577901
transform 1 0 42528 0 1 7560
box -48 -56 432 834
use sg13g2_fill_2  FILLER_8_435
timestamp 1677580104
transform 1 0 42912 0 1 7560
box -48 -56 240 834
use sg13g2_decap_8  FILLER_8_441
timestamp 1679581782
transform 1 0 43488 0 1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_8_448
timestamp 1677580104
transform 1 0 44160 0 1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_450
timestamp 1677579658
transform 1 0 44352 0 1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_0
timestamp 1679581782
transform 1 0 1152 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_7
timestamp 1679581782
transform 1 0 1824 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_14
timestamp 1679581782
transform 1 0 2496 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_21
timestamp 1679581782
transform 1 0 3168 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_28
timestamp 1679581782
transform 1 0 3840 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_35
timestamp 1679581782
transform 1 0 4512 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_42
timestamp 1679581782
transform 1 0 5184 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_49
timestamp 1679581782
transform 1 0 5856 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_56
timestamp 1679581782
transform 1 0 6528 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_63
timestamp 1679581782
transform 1 0 7200 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_70
timestamp 1679581782
transform 1 0 7872 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_77
timestamp 1679581782
transform 1 0 8544 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_84
timestamp 1679581782
transform 1 0 9216 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_91
timestamp 1679581782
transform 1 0 9888 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_4  FILLER_9_98
timestamp 1679577901
transform 1 0 10560 0 -1 9072
box -48 -56 432 834
use sg13g2_fill_1  FILLER_9_102
timestamp 1677579658
transform 1 0 10944 0 -1 9072
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_199
timestamp 1679581782
transform 1 0 20256 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_206
timestamp 1679581782
transform 1 0 20928 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_213
timestamp 1679581782
transform 1 0 21600 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_220
timestamp 1679581782
transform 1 0 22272 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_227
timestamp 1679581782
transform 1 0 22944 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_234
timestamp 1679581782
transform 1 0 23616 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_241
timestamp 1679581782
transform 1 0 24288 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_248
timestamp 1679581782
transform 1 0 24960 0 -1 9072
box -48 -56 720 834
use sg13g2_fill_2  FILLER_9_255
timestamp 1677580104
transform 1 0 25632 0 -1 9072
box -48 -56 240 834
use sg13g2_fill_2  FILLER_9_261
timestamp 1677580104
transform 1 0 26208 0 -1 9072
box -48 -56 240 834
use sg13g2_decap_4  FILLER_9_267
timestamp 1679577901
transform 1 0 26784 0 -1 9072
box -48 -56 432 834
use sg13g2_decap_8  FILLER_9_291
timestamp 1679581782
transform 1 0 29088 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_298
timestamp 1679581782
transform 1 0 29760 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_305
timestamp 1679581782
transform 1 0 30432 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_312
timestamp 1679581782
transform 1 0 31104 0 -1 9072
box -48 -56 720 834
use sg13g2_fill_1  FILLER_9_339
timestamp 1677579658
transform 1 0 33696 0 -1 9072
box -48 -56 144 834
use sg13g2_fill_1  FILLER_9_359
timestamp 1677579658
transform 1 0 35616 0 -1 9072
box -48 -56 144 834
use sg13g2_fill_1  FILLER_9_374
timestamp 1677579658
transform 1 0 37056 0 -1 9072
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_410
timestamp 1679581782
transform 1 0 40512 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_417
timestamp 1679581782
transform 1 0 41184 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_424
timestamp 1679581782
transform 1 0 41856 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_431
timestamp 1679581782
transform 1 0 42528 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_4  FILLER_9_438
timestamp 1679577901
transform 1 0 43200 0 -1 9072
box -48 -56 432 834
use sg13g2_fill_1  FILLER_9_442
timestamp 1677579658
transform 1 0 43584 0 -1 9072
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_0
timestamp 1679581782
transform 1 0 1152 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_7
timestamp 1679581782
transform 1 0 1824 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_14
timestamp 1679581782
transform 1 0 2496 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_21
timestamp 1679581782
transform 1 0 3168 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_28
timestamp 1679581782
transform 1 0 3840 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_35
timestamp 1679581782
transform 1 0 4512 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_42
timestamp 1679581782
transform 1 0 5184 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_49
timestamp 1679581782
transform 1 0 5856 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_56
timestamp 1679581782
transform 1 0 6528 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_63
timestamp 1679581782
transform 1 0 7200 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_70
timestamp 1679581782
transform 1 0 7872 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_77
timestamp 1679581782
transform 1 0 8544 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_84
timestamp 1679581782
transform 1 0 9216 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_91
timestamp 1679581782
transform 1 0 9888 0 1 9072
box -48 -56 720 834
use sg13g2_fill_1  FILLER_10_98
timestamp 1677579658
transform 1 0 10560 0 1 9072
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_215
timestamp 1679581782
transform 1 0 21792 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_222
timestamp 1679581782
transform 1 0 22464 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_229
timestamp 1679581782
transform 1 0 23136 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_236
timestamp 1679581782
transform 1 0 23808 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_243
timestamp 1679581782
transform 1 0 24480 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_250
timestamp 1679581782
transform 1 0 25152 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_257
timestamp 1679581782
transform 1 0 25824 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_264
timestamp 1679581782
transform 1 0 26496 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_271
timestamp 1679581782
transform 1 0 27168 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_278
timestamp 1679581782
transform 1 0 27840 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_285
timestamp 1679581782
transform 1 0 28512 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_292
timestamp 1679581782
transform 1 0 29184 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_299
timestamp 1679581782
transform 1 0 29856 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_306
timestamp 1679581782
transform 1 0 30528 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_415
timestamp 1679581782
transform 1 0 40992 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_422
timestamp 1679581782
transform 1 0 41664 0 1 9072
box -48 -56 720 834
use sg13g2_decap_4  FILLER_10_429
timestamp 1679577901
transform 1 0 42336 0 1 9072
box -48 -56 432 834
use sg13g2_fill_2  FILLER_10_433
timestamp 1677580104
transform 1 0 42720 0 1 9072
box -48 -56 240 834
use sg13g2_buf_1  output1
timestamp 1676381911
transform 1 0 44064 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output2
timestamp 1676381911
transform 1 0 44448 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output3
timestamp 1676381911
transform 1 0 44832 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output4
timestamp 1676381911
transform 1 0 44448 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output5
timestamp 1676381911
transform 1 0 44832 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output6
timestamp 1676381911
transform 1 0 44448 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output7
timestamp 1676381911
transform 1 0 44832 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output8
timestamp 1676381911
transform 1 0 44448 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  output9
timestamp 1676381911
transform 1 0 44832 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  output10
timestamp 1676381911
transform 1 0 44448 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  output11
timestamp 1676381911
transform 1 0 44832 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  output12
timestamp 1676381911
transform 1 0 43680 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output13
timestamp 1676381911
transform 1 0 44832 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  output14
timestamp 1676381911
transform 1 0 44448 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  output15
timestamp 1676381911
transform 1 0 44832 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output16
timestamp 1676381911
transform 1 0 44448 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output17
timestamp 1676381911
transform 1 0 44832 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output18
timestamp 1676381911
transform 1 0 44448 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output19
timestamp 1676381911
transform 1 0 44064 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output20
timestamp 1676381911
transform 1 0 43680 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output21
timestamp 1676381911
transform 1 0 44064 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output22
timestamp 1676381911
transform 1 0 43296 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output23
timestamp 1676381911
transform 1 0 43296 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output24
timestamp 1676381911
transform 1 0 42912 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output25
timestamp 1676381911
transform 1 0 43680 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output26
timestamp 1676381911
transform 1 0 44448 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output27
timestamp 1676381911
transform 1 0 44064 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output28
timestamp 1676381911
transform 1 0 44832 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output29
timestamp 1676381911
transform 1 0 44448 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output30
timestamp 1676381911
transform 1 0 44832 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output31
timestamp 1676381911
transform 1 0 44448 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output32
timestamp 1676381911
transform 1 0 44832 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output33
timestamp 1676381911
transform -1 0 31968 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output34
timestamp 1676381911
transform -1 0 33696 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output35
timestamp 1676381911
transform -1 0 34656 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output36
timestamp 1676381911
transform -1 0 35040 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output37
timestamp 1676381911
transform -1 0 35424 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output38
timestamp 1676381911
transform -1 0 35808 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output39
timestamp 1676381911
transform -1 0 35232 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output40
timestamp 1676381911
transform -1 0 36192 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output41
timestamp 1676381911
transform -1 0 35616 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output42
timestamp 1676381911
transform -1 0 36576 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output43
timestamp 1676381911
transform -1 0 36960 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output44
timestamp 1676381911
transform -1 0 32352 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output45
timestamp 1676381911
transform -1 0 32736 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output46
timestamp 1676381911
transform -1 0 33120 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output47
timestamp 1676381911
transform -1 0 32544 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output48
timestamp 1676381911
transform -1 0 33504 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output49
timestamp 1676381911
transform -1 0 32928 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output50
timestamp 1676381911
transform -1 0 33888 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output51
timestamp 1676381911
transform -1 0 33312 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output52
timestamp 1676381911
transform -1 0 34272 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output53
timestamp 1676381911
transform -1 0 11424 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output54
timestamp 1676381911
transform 1 0 10656 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output55
timestamp 1676381911
transform -1 0 11808 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output56
timestamp 1676381911
transform 1 0 11040 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output57
timestamp 1676381911
transform -1 0 12192 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output58
timestamp 1676381911
transform 1 0 11424 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output59
timestamp 1676381911
transform -1 0 12576 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output60
timestamp 1676381911
transform 1 0 11808 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output61
timestamp 1676381911
transform -1 0 12960 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output62
timestamp 1676381911
transform 1 0 12192 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output63
timestamp 1676381911
transform -1 0 13344 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output64
timestamp 1676381911
transform 1 0 12576 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output65
timestamp 1676381911
transform -1 0 13728 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output66
timestamp 1676381911
transform 1 0 12960 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output67
timestamp 1676381911
transform -1 0 14112 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output68
timestamp 1676381911
transform 1 0 13344 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output69
timestamp 1676381911
transform -1 0 14496 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output70
timestamp 1676381911
transform 1 0 13728 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output71
timestamp 1676381911
transform -1 0 14880 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output72
timestamp 1676381911
transform 1 0 14112 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output73
timestamp 1676381911
transform -1 0 15264 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output74
timestamp 1676381911
transform -1 0 17184 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output75
timestamp 1676381911
transform 1 0 16416 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output76
timestamp 1676381911
transform -1 0 17568 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output77
timestamp 1676381911
transform 1 0 16800 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output78
timestamp 1676381911
transform -1 0 17952 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output79
timestamp 1676381911
transform 1 0 17184 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output80
timestamp 1676381911
transform 1 0 14496 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output81
timestamp 1676381911
transform -1 0 15648 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output82
timestamp 1676381911
transform 1 0 14880 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output83
timestamp 1676381911
transform -1 0 16032 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output84
timestamp 1676381911
transform 1 0 15264 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output85
timestamp 1676381911
transform -1 0 16416 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output86
timestamp 1676381911
transform 1 0 15648 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output87
timestamp 1676381911
transform -1 0 16800 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output88
timestamp 1676381911
transform 1 0 16032 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output89
timestamp 1676381911
transform -1 0 18336 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output90
timestamp 1676381911
transform -1 0 20256 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output91
timestamp 1676381911
transform 1 0 19488 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output92
timestamp 1676381911
transform 1 0 19872 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output93
timestamp 1676381911
transform -1 0 20640 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output94
timestamp 1676381911
transform -1 0 21024 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output95
timestamp 1676381911
transform -1 0 21792 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output96
timestamp 1676381911
transform 1 0 17568 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output97
timestamp 1676381911
transform -1 0 18720 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output98
timestamp 1676381911
transform 1 0 17952 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output99
timestamp 1676381911
transform -1 0 19104 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output100
timestamp 1676381911
transform 1 0 18336 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output101
timestamp 1676381911
transform -1 0 19488 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output102
timestamp 1676381911
transform 1 0 18720 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output103
timestamp 1676381911
transform -1 0 19872 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output104
timestamp 1676381911
transform 1 0 19104 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output105
timestamp 1676381911
transform -1 0 31584 0 1 9072
box -48 -56 432 834
use sg13g2_tielo  S_term_single_106
timestamp 1680000637
transform -1 0 21408 0 1 9072
box -48 -56 432 834
<< labels >>
flabel metal3 s 20984 11764 21064 11844 0 FreeSans 320 0 0 0 Co
port 0 nsew signal output
flabel metal2 s 0 548 90 628 0 FreeSans 320 0 0 0 FrameData[0]
port 1 nsew signal input
flabel metal2 s 0 3908 90 3988 0 FreeSans 320 0 0 0 FrameData[10]
port 2 nsew signal input
flabel metal2 s 0 4244 90 4324 0 FreeSans 320 0 0 0 FrameData[11]
port 3 nsew signal input
flabel metal2 s 0 4580 90 4660 0 FreeSans 320 0 0 0 FrameData[12]
port 4 nsew signal input
flabel metal2 s 0 4916 90 4996 0 FreeSans 320 0 0 0 FrameData[13]
port 5 nsew signal input
flabel metal2 s 0 5252 90 5332 0 FreeSans 320 0 0 0 FrameData[14]
port 6 nsew signal input
flabel metal2 s 0 5588 90 5668 0 FreeSans 320 0 0 0 FrameData[15]
port 7 nsew signal input
flabel metal2 s 0 5924 90 6004 0 FreeSans 320 0 0 0 FrameData[16]
port 8 nsew signal input
flabel metal2 s 0 6260 90 6340 0 FreeSans 320 0 0 0 FrameData[17]
port 9 nsew signal input
flabel metal2 s 0 6596 90 6676 0 FreeSans 320 0 0 0 FrameData[18]
port 10 nsew signal input
flabel metal2 s 0 6932 90 7012 0 FreeSans 320 0 0 0 FrameData[19]
port 11 nsew signal input
flabel metal2 s 0 884 90 964 0 FreeSans 320 0 0 0 FrameData[1]
port 12 nsew signal input
flabel metal2 s 0 7268 90 7348 0 FreeSans 320 0 0 0 FrameData[20]
port 13 nsew signal input
flabel metal2 s 0 7604 90 7684 0 FreeSans 320 0 0 0 FrameData[21]
port 14 nsew signal input
flabel metal2 s 0 7940 90 8020 0 FreeSans 320 0 0 0 FrameData[22]
port 15 nsew signal input
flabel metal2 s 0 8276 90 8356 0 FreeSans 320 0 0 0 FrameData[23]
port 16 nsew signal input
flabel metal2 s 0 8612 90 8692 0 FreeSans 320 0 0 0 FrameData[24]
port 17 nsew signal input
flabel metal2 s 0 8948 90 9028 0 FreeSans 320 0 0 0 FrameData[25]
port 18 nsew signal input
flabel metal2 s 0 9284 90 9364 0 FreeSans 320 0 0 0 FrameData[26]
port 19 nsew signal input
flabel metal2 s 0 9620 90 9700 0 FreeSans 320 0 0 0 FrameData[27]
port 20 nsew signal input
flabel metal2 s 0 9956 90 10036 0 FreeSans 320 0 0 0 FrameData[28]
port 21 nsew signal input
flabel metal2 s 0 10292 90 10372 0 FreeSans 320 0 0 0 FrameData[29]
port 22 nsew signal input
flabel metal2 s 0 1220 90 1300 0 FreeSans 320 0 0 0 FrameData[2]
port 23 nsew signal input
flabel metal2 s 0 10628 90 10708 0 FreeSans 320 0 0 0 FrameData[30]
port 24 nsew signal input
flabel metal2 s 0 10964 90 11044 0 FreeSans 320 0 0 0 FrameData[31]
port 25 nsew signal input
flabel metal2 s 0 1556 90 1636 0 FreeSans 320 0 0 0 FrameData[3]
port 26 nsew signal input
flabel metal2 s 0 1892 90 1972 0 FreeSans 320 0 0 0 FrameData[4]
port 27 nsew signal input
flabel metal2 s 0 2228 90 2308 0 FreeSans 320 0 0 0 FrameData[5]
port 28 nsew signal input
flabel metal2 s 0 2564 90 2644 0 FreeSans 320 0 0 0 FrameData[6]
port 29 nsew signal input
flabel metal2 s 0 2900 90 2980 0 FreeSans 320 0 0 0 FrameData[7]
port 30 nsew signal input
flabel metal2 s 0 3236 90 3316 0 FreeSans 320 0 0 0 FrameData[8]
port 31 nsew signal input
flabel metal2 s 0 3572 90 3652 0 FreeSans 320 0 0 0 FrameData[9]
port 32 nsew signal input
flabel metal2 s 46278 548 46368 628 0 FreeSans 320 0 0 0 FrameData_O[0]
port 33 nsew signal output
flabel metal2 s 46278 3908 46368 3988 0 FreeSans 320 0 0 0 FrameData_O[10]
port 34 nsew signal output
flabel metal2 s 46278 4244 46368 4324 0 FreeSans 320 0 0 0 FrameData_O[11]
port 35 nsew signal output
flabel metal2 s 46278 4580 46368 4660 0 FreeSans 320 0 0 0 FrameData_O[12]
port 36 nsew signal output
flabel metal2 s 46278 4916 46368 4996 0 FreeSans 320 0 0 0 FrameData_O[13]
port 37 nsew signal output
flabel metal2 s 46278 5252 46368 5332 0 FreeSans 320 0 0 0 FrameData_O[14]
port 38 nsew signal output
flabel metal2 s 46278 5588 46368 5668 0 FreeSans 320 0 0 0 FrameData_O[15]
port 39 nsew signal output
flabel metal2 s 46278 5924 46368 6004 0 FreeSans 320 0 0 0 FrameData_O[16]
port 40 nsew signal output
flabel metal2 s 46278 6260 46368 6340 0 FreeSans 320 0 0 0 FrameData_O[17]
port 41 nsew signal output
flabel metal2 s 46278 6596 46368 6676 0 FreeSans 320 0 0 0 FrameData_O[18]
port 42 nsew signal output
flabel metal2 s 46278 6932 46368 7012 0 FreeSans 320 0 0 0 FrameData_O[19]
port 43 nsew signal output
flabel metal2 s 46278 884 46368 964 0 FreeSans 320 0 0 0 FrameData_O[1]
port 44 nsew signal output
flabel metal2 s 46278 7268 46368 7348 0 FreeSans 320 0 0 0 FrameData_O[20]
port 45 nsew signal output
flabel metal2 s 46278 7604 46368 7684 0 FreeSans 320 0 0 0 FrameData_O[21]
port 46 nsew signal output
flabel metal2 s 46278 7940 46368 8020 0 FreeSans 320 0 0 0 FrameData_O[22]
port 47 nsew signal output
flabel metal2 s 46278 8276 46368 8356 0 FreeSans 320 0 0 0 FrameData_O[23]
port 48 nsew signal output
flabel metal2 s 46278 8612 46368 8692 0 FreeSans 320 0 0 0 FrameData_O[24]
port 49 nsew signal output
flabel metal2 s 46278 8948 46368 9028 0 FreeSans 320 0 0 0 FrameData_O[25]
port 50 nsew signal output
flabel metal2 s 46278 9284 46368 9364 0 FreeSans 320 0 0 0 FrameData_O[26]
port 51 nsew signal output
flabel metal2 s 46278 9620 46368 9700 0 FreeSans 320 0 0 0 FrameData_O[27]
port 52 nsew signal output
flabel metal2 s 46278 9956 46368 10036 0 FreeSans 320 0 0 0 FrameData_O[28]
port 53 nsew signal output
flabel metal2 s 46278 10292 46368 10372 0 FreeSans 320 0 0 0 FrameData_O[29]
port 54 nsew signal output
flabel metal2 s 46278 1220 46368 1300 0 FreeSans 320 0 0 0 FrameData_O[2]
port 55 nsew signal output
flabel metal2 s 46278 10628 46368 10708 0 FreeSans 320 0 0 0 FrameData_O[30]
port 56 nsew signal output
flabel metal2 s 46278 10964 46368 11044 0 FreeSans 320 0 0 0 FrameData_O[31]
port 57 nsew signal output
flabel metal2 s 46278 1556 46368 1636 0 FreeSans 320 0 0 0 FrameData_O[3]
port 58 nsew signal output
flabel metal2 s 46278 1892 46368 1972 0 FreeSans 320 0 0 0 FrameData_O[4]
port 59 nsew signal output
flabel metal2 s 46278 2228 46368 2308 0 FreeSans 320 0 0 0 FrameData_O[5]
port 60 nsew signal output
flabel metal2 s 46278 2564 46368 2644 0 FreeSans 320 0 0 0 FrameData_O[6]
port 61 nsew signal output
flabel metal2 s 46278 2900 46368 2980 0 FreeSans 320 0 0 0 FrameData_O[7]
port 62 nsew signal output
flabel metal2 s 46278 3236 46368 3316 0 FreeSans 320 0 0 0 FrameData_O[8]
port 63 nsew signal output
flabel metal2 s 46278 3572 46368 3652 0 FreeSans 320 0 0 0 FrameData_O[9]
port 64 nsew signal output
flabel metal3 s 4088 0 4168 80 0 FreeSans 320 0 0 0 FrameStrobe[0]
port 65 nsew signal input
flabel metal3 s 25208 0 25288 80 0 FreeSans 320 0 0 0 FrameStrobe[10]
port 66 nsew signal input
flabel metal3 s 27320 0 27400 80 0 FreeSans 320 0 0 0 FrameStrobe[11]
port 67 nsew signal input
flabel metal3 s 29432 0 29512 80 0 FreeSans 320 0 0 0 FrameStrobe[12]
port 68 nsew signal input
flabel metal3 s 31544 0 31624 80 0 FreeSans 320 0 0 0 FrameStrobe[13]
port 69 nsew signal input
flabel metal3 s 33656 0 33736 80 0 FreeSans 320 0 0 0 FrameStrobe[14]
port 70 nsew signal input
flabel metal3 s 35768 0 35848 80 0 FreeSans 320 0 0 0 FrameStrobe[15]
port 71 nsew signal input
flabel metal3 s 37880 0 37960 80 0 FreeSans 320 0 0 0 FrameStrobe[16]
port 72 nsew signal input
flabel metal3 s 39992 0 40072 80 0 FreeSans 320 0 0 0 FrameStrobe[17]
port 73 nsew signal input
flabel metal3 s 42104 0 42184 80 0 FreeSans 320 0 0 0 FrameStrobe[18]
port 74 nsew signal input
flabel metal3 s 44216 0 44296 80 0 FreeSans 320 0 0 0 FrameStrobe[19]
port 75 nsew signal input
flabel metal3 s 6200 0 6280 80 0 FreeSans 320 0 0 0 FrameStrobe[1]
port 76 nsew signal input
flabel metal3 s 8312 0 8392 80 0 FreeSans 320 0 0 0 FrameStrobe[2]
port 77 nsew signal input
flabel metal3 s 10424 0 10504 80 0 FreeSans 320 0 0 0 FrameStrobe[3]
port 78 nsew signal input
flabel metal3 s 12536 0 12616 80 0 FreeSans 320 0 0 0 FrameStrobe[4]
port 79 nsew signal input
flabel metal3 s 14648 0 14728 80 0 FreeSans 320 0 0 0 FrameStrobe[5]
port 80 nsew signal input
flabel metal3 s 16760 0 16840 80 0 FreeSans 320 0 0 0 FrameStrobe[6]
port 81 nsew signal input
flabel metal3 s 18872 0 18952 80 0 FreeSans 320 0 0 0 FrameStrobe[7]
port 82 nsew signal input
flabel metal3 s 20984 0 21064 80 0 FreeSans 320 0 0 0 FrameStrobe[8]
port 83 nsew signal input
flabel metal3 s 23096 0 23176 80 0 FreeSans 320 0 0 0 FrameStrobe[9]
port 84 nsew signal input
flabel metal3 s 31352 11764 31432 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[0]
port 85 nsew signal output
flabel metal3 s 33272 11764 33352 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[10]
port 86 nsew signal output
flabel metal3 s 33464 11764 33544 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[11]
port 87 nsew signal output
flabel metal3 s 33656 11764 33736 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[12]
port 88 nsew signal output
flabel metal3 s 33848 11764 33928 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[13]
port 89 nsew signal output
flabel metal3 s 34040 11764 34120 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[14]
port 90 nsew signal output
flabel metal3 s 34232 11764 34312 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[15]
port 91 nsew signal output
flabel metal3 s 34424 11764 34504 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[16]
port 92 nsew signal output
flabel metal3 s 34616 11764 34696 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[17]
port 93 nsew signal output
flabel metal3 s 34808 11764 34888 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[18]
port 94 nsew signal output
flabel metal3 s 35000 11764 35080 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[19]
port 95 nsew signal output
flabel metal3 s 31544 11764 31624 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[1]
port 96 nsew signal output
flabel metal3 s 31736 11764 31816 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[2]
port 97 nsew signal output
flabel metal3 s 31928 11764 32008 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[3]
port 98 nsew signal output
flabel metal3 s 32120 11764 32200 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[4]
port 99 nsew signal output
flabel metal3 s 32312 11764 32392 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[5]
port 100 nsew signal output
flabel metal3 s 32504 11764 32584 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[6]
port 101 nsew signal output
flabel metal3 s 32696 11764 32776 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[7]
port 102 nsew signal output
flabel metal3 s 32888 11764 32968 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[8]
port 103 nsew signal output
flabel metal3 s 33080 11764 33160 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[9]
port 104 nsew signal output
flabel metal3 s 11000 11764 11080 11844 0 FreeSans 320 0 0 0 N1BEG[0]
port 105 nsew signal output
flabel metal3 s 11192 11764 11272 11844 0 FreeSans 320 0 0 0 N1BEG[1]
port 106 nsew signal output
flabel metal3 s 11384 11764 11464 11844 0 FreeSans 320 0 0 0 N1BEG[2]
port 107 nsew signal output
flabel metal3 s 11576 11764 11656 11844 0 FreeSans 320 0 0 0 N1BEG[3]
port 108 nsew signal output
flabel metal3 s 11768 11764 11848 11844 0 FreeSans 320 0 0 0 N2BEG[0]
port 109 nsew signal output
flabel metal3 s 11960 11764 12040 11844 0 FreeSans 320 0 0 0 N2BEG[1]
port 110 nsew signal output
flabel metal3 s 12152 11764 12232 11844 0 FreeSans 320 0 0 0 N2BEG[2]
port 111 nsew signal output
flabel metal3 s 12344 11764 12424 11844 0 FreeSans 320 0 0 0 N2BEG[3]
port 112 nsew signal output
flabel metal3 s 12536 11764 12616 11844 0 FreeSans 320 0 0 0 N2BEG[4]
port 113 nsew signal output
flabel metal3 s 12728 11764 12808 11844 0 FreeSans 320 0 0 0 N2BEG[5]
port 114 nsew signal output
flabel metal3 s 12920 11764 13000 11844 0 FreeSans 320 0 0 0 N2BEG[6]
port 115 nsew signal output
flabel metal3 s 13112 11764 13192 11844 0 FreeSans 320 0 0 0 N2BEG[7]
port 116 nsew signal output
flabel metal3 s 13304 11764 13384 11844 0 FreeSans 320 0 0 0 N2BEGb[0]
port 117 nsew signal output
flabel metal3 s 13496 11764 13576 11844 0 FreeSans 320 0 0 0 N2BEGb[1]
port 118 nsew signal output
flabel metal3 s 13688 11764 13768 11844 0 FreeSans 320 0 0 0 N2BEGb[2]
port 119 nsew signal output
flabel metal3 s 13880 11764 13960 11844 0 FreeSans 320 0 0 0 N2BEGb[3]
port 120 nsew signal output
flabel metal3 s 14072 11764 14152 11844 0 FreeSans 320 0 0 0 N2BEGb[4]
port 121 nsew signal output
flabel metal3 s 14264 11764 14344 11844 0 FreeSans 320 0 0 0 N2BEGb[5]
port 122 nsew signal output
flabel metal3 s 14456 11764 14536 11844 0 FreeSans 320 0 0 0 N2BEGb[6]
port 123 nsew signal output
flabel metal3 s 14648 11764 14728 11844 0 FreeSans 320 0 0 0 N2BEGb[7]
port 124 nsew signal output
flabel metal3 s 14840 11764 14920 11844 0 FreeSans 320 0 0 0 N4BEG[0]
port 125 nsew signal output
flabel metal3 s 16760 11764 16840 11844 0 FreeSans 320 0 0 0 N4BEG[10]
port 126 nsew signal output
flabel metal3 s 16952 11764 17032 11844 0 FreeSans 320 0 0 0 N4BEG[11]
port 127 nsew signal output
flabel metal3 s 17144 11764 17224 11844 0 FreeSans 320 0 0 0 N4BEG[12]
port 128 nsew signal output
flabel metal3 s 17336 11764 17416 11844 0 FreeSans 320 0 0 0 N4BEG[13]
port 129 nsew signal output
flabel metal3 s 17528 11764 17608 11844 0 FreeSans 320 0 0 0 N4BEG[14]
port 130 nsew signal output
flabel metal3 s 17720 11764 17800 11844 0 FreeSans 320 0 0 0 N4BEG[15]
port 131 nsew signal output
flabel metal3 s 15032 11764 15112 11844 0 FreeSans 320 0 0 0 N4BEG[1]
port 132 nsew signal output
flabel metal3 s 15224 11764 15304 11844 0 FreeSans 320 0 0 0 N4BEG[2]
port 133 nsew signal output
flabel metal3 s 15416 11764 15496 11844 0 FreeSans 320 0 0 0 N4BEG[3]
port 134 nsew signal output
flabel metal3 s 15608 11764 15688 11844 0 FreeSans 320 0 0 0 N4BEG[4]
port 135 nsew signal output
flabel metal3 s 15800 11764 15880 11844 0 FreeSans 320 0 0 0 N4BEG[5]
port 136 nsew signal output
flabel metal3 s 15992 11764 16072 11844 0 FreeSans 320 0 0 0 N4BEG[6]
port 137 nsew signal output
flabel metal3 s 16184 11764 16264 11844 0 FreeSans 320 0 0 0 N4BEG[7]
port 138 nsew signal output
flabel metal3 s 16376 11764 16456 11844 0 FreeSans 320 0 0 0 N4BEG[8]
port 139 nsew signal output
flabel metal3 s 16568 11764 16648 11844 0 FreeSans 320 0 0 0 N4BEG[9]
port 140 nsew signal output
flabel metal3 s 17912 11764 17992 11844 0 FreeSans 320 0 0 0 NN4BEG[0]
port 141 nsew signal output
flabel metal3 s 19832 11764 19912 11844 0 FreeSans 320 0 0 0 NN4BEG[10]
port 142 nsew signal output
flabel metal3 s 20024 11764 20104 11844 0 FreeSans 320 0 0 0 NN4BEG[11]
port 143 nsew signal output
flabel metal3 s 20216 11764 20296 11844 0 FreeSans 320 0 0 0 NN4BEG[12]
port 144 nsew signal output
flabel metal3 s 20408 11764 20488 11844 0 FreeSans 320 0 0 0 NN4BEG[13]
port 145 nsew signal output
flabel metal3 s 20600 11764 20680 11844 0 FreeSans 320 0 0 0 NN4BEG[14]
port 146 nsew signal output
flabel metal3 s 20792 11764 20872 11844 0 FreeSans 320 0 0 0 NN4BEG[15]
port 147 nsew signal output
flabel metal3 s 18104 11764 18184 11844 0 FreeSans 320 0 0 0 NN4BEG[1]
port 148 nsew signal output
flabel metal3 s 18296 11764 18376 11844 0 FreeSans 320 0 0 0 NN4BEG[2]
port 149 nsew signal output
flabel metal3 s 18488 11764 18568 11844 0 FreeSans 320 0 0 0 NN4BEG[3]
port 150 nsew signal output
flabel metal3 s 18680 11764 18760 11844 0 FreeSans 320 0 0 0 NN4BEG[4]
port 151 nsew signal output
flabel metal3 s 18872 11764 18952 11844 0 FreeSans 320 0 0 0 NN4BEG[5]
port 152 nsew signal output
flabel metal3 s 19064 11764 19144 11844 0 FreeSans 320 0 0 0 NN4BEG[6]
port 153 nsew signal output
flabel metal3 s 19256 11764 19336 11844 0 FreeSans 320 0 0 0 NN4BEG[7]
port 154 nsew signal output
flabel metal3 s 19448 11764 19528 11844 0 FreeSans 320 0 0 0 NN4BEG[8]
port 155 nsew signal output
flabel metal3 s 19640 11764 19720 11844 0 FreeSans 320 0 0 0 NN4BEG[9]
port 156 nsew signal output
flabel metal3 s 21176 11764 21256 11844 0 FreeSans 320 0 0 0 S1END[0]
port 157 nsew signal input
flabel metal3 s 21368 11764 21448 11844 0 FreeSans 320 0 0 0 S1END[1]
port 158 nsew signal input
flabel metal3 s 21560 11764 21640 11844 0 FreeSans 320 0 0 0 S1END[2]
port 159 nsew signal input
flabel metal3 s 21752 11764 21832 11844 0 FreeSans 320 0 0 0 S1END[3]
port 160 nsew signal input
flabel metal3 s 23480 11764 23560 11844 0 FreeSans 320 0 0 0 S2END[0]
port 161 nsew signal input
flabel metal3 s 23672 11764 23752 11844 0 FreeSans 320 0 0 0 S2END[1]
port 162 nsew signal input
flabel metal3 s 23864 11764 23944 11844 0 FreeSans 320 0 0 0 S2END[2]
port 163 nsew signal input
flabel metal3 s 24056 11764 24136 11844 0 FreeSans 320 0 0 0 S2END[3]
port 164 nsew signal input
flabel metal3 s 24248 11764 24328 11844 0 FreeSans 320 0 0 0 S2END[4]
port 165 nsew signal input
flabel metal3 s 24440 11764 24520 11844 0 FreeSans 320 0 0 0 S2END[5]
port 166 nsew signal input
flabel metal3 s 24632 11764 24712 11844 0 FreeSans 320 0 0 0 S2END[6]
port 167 nsew signal input
flabel metal3 s 24824 11764 24904 11844 0 FreeSans 320 0 0 0 S2END[7]
port 168 nsew signal input
flabel metal3 s 21944 11764 22024 11844 0 FreeSans 320 0 0 0 S2MID[0]
port 169 nsew signal input
flabel metal3 s 22136 11764 22216 11844 0 FreeSans 320 0 0 0 S2MID[1]
port 170 nsew signal input
flabel metal3 s 22328 11764 22408 11844 0 FreeSans 320 0 0 0 S2MID[2]
port 171 nsew signal input
flabel metal3 s 22520 11764 22600 11844 0 FreeSans 320 0 0 0 S2MID[3]
port 172 nsew signal input
flabel metal3 s 22712 11764 22792 11844 0 FreeSans 320 0 0 0 S2MID[4]
port 173 nsew signal input
flabel metal3 s 22904 11764 22984 11844 0 FreeSans 320 0 0 0 S2MID[5]
port 174 nsew signal input
flabel metal3 s 23096 11764 23176 11844 0 FreeSans 320 0 0 0 S2MID[6]
port 175 nsew signal input
flabel metal3 s 23288 11764 23368 11844 0 FreeSans 320 0 0 0 S2MID[7]
port 176 nsew signal input
flabel metal3 s 25016 11764 25096 11844 0 FreeSans 320 0 0 0 S4END[0]
port 177 nsew signal input
flabel metal3 s 26936 11764 27016 11844 0 FreeSans 320 0 0 0 S4END[10]
port 178 nsew signal input
flabel metal3 s 27128 11764 27208 11844 0 FreeSans 320 0 0 0 S4END[11]
port 179 nsew signal input
flabel metal3 s 27320 11764 27400 11844 0 FreeSans 320 0 0 0 S4END[12]
port 180 nsew signal input
flabel metal3 s 27512 11764 27592 11844 0 FreeSans 320 0 0 0 S4END[13]
port 181 nsew signal input
flabel metal3 s 27704 11764 27784 11844 0 FreeSans 320 0 0 0 S4END[14]
port 182 nsew signal input
flabel metal3 s 27896 11764 27976 11844 0 FreeSans 320 0 0 0 S4END[15]
port 183 nsew signal input
flabel metal3 s 25208 11764 25288 11844 0 FreeSans 320 0 0 0 S4END[1]
port 184 nsew signal input
flabel metal3 s 25400 11764 25480 11844 0 FreeSans 320 0 0 0 S4END[2]
port 185 nsew signal input
flabel metal3 s 25592 11764 25672 11844 0 FreeSans 320 0 0 0 S4END[3]
port 186 nsew signal input
flabel metal3 s 25784 11764 25864 11844 0 FreeSans 320 0 0 0 S4END[4]
port 187 nsew signal input
flabel metal3 s 25976 11764 26056 11844 0 FreeSans 320 0 0 0 S4END[5]
port 188 nsew signal input
flabel metal3 s 26168 11764 26248 11844 0 FreeSans 320 0 0 0 S4END[6]
port 189 nsew signal input
flabel metal3 s 26360 11764 26440 11844 0 FreeSans 320 0 0 0 S4END[7]
port 190 nsew signal input
flabel metal3 s 26552 11764 26632 11844 0 FreeSans 320 0 0 0 S4END[8]
port 191 nsew signal input
flabel metal3 s 26744 11764 26824 11844 0 FreeSans 320 0 0 0 S4END[9]
port 192 nsew signal input
flabel metal3 s 28088 11764 28168 11844 0 FreeSans 320 0 0 0 SS4END[0]
port 193 nsew signal input
flabel metal3 s 30008 11764 30088 11844 0 FreeSans 320 0 0 0 SS4END[10]
port 194 nsew signal input
flabel metal3 s 30200 11764 30280 11844 0 FreeSans 320 0 0 0 SS4END[11]
port 195 nsew signal input
flabel metal3 s 30392 11764 30472 11844 0 FreeSans 320 0 0 0 SS4END[12]
port 196 nsew signal input
flabel metal3 s 30584 11764 30664 11844 0 FreeSans 320 0 0 0 SS4END[13]
port 197 nsew signal input
flabel metal3 s 30776 11764 30856 11844 0 FreeSans 320 0 0 0 SS4END[14]
port 198 nsew signal input
flabel metal3 s 30968 11764 31048 11844 0 FreeSans 320 0 0 0 SS4END[15]
port 199 nsew signal input
flabel metal3 s 28280 11764 28360 11844 0 FreeSans 320 0 0 0 SS4END[1]
port 200 nsew signal input
flabel metal3 s 28472 11764 28552 11844 0 FreeSans 320 0 0 0 SS4END[2]
port 201 nsew signal input
flabel metal3 s 28664 11764 28744 11844 0 FreeSans 320 0 0 0 SS4END[3]
port 202 nsew signal input
flabel metal3 s 28856 11764 28936 11844 0 FreeSans 320 0 0 0 SS4END[4]
port 203 nsew signal input
flabel metal3 s 29048 11764 29128 11844 0 FreeSans 320 0 0 0 SS4END[5]
port 204 nsew signal input
flabel metal3 s 29240 11764 29320 11844 0 FreeSans 320 0 0 0 SS4END[6]
port 205 nsew signal input
flabel metal3 s 29432 11764 29512 11844 0 FreeSans 320 0 0 0 SS4END[7]
port 206 nsew signal input
flabel metal3 s 29624 11764 29704 11844 0 FreeSans 320 0 0 0 SS4END[8]
port 207 nsew signal input
flabel metal3 s 29816 11764 29896 11844 0 FreeSans 320 0 0 0 SS4END[9]
port 208 nsew signal input
flabel metal3 s 1976 0 2056 80 0 FreeSans 320 0 0 0 UserCLK
port 209 nsew signal input
flabel metal3 s 31160 11764 31240 11844 0 FreeSans 320 0 0 0 UserCLKo
port 210 nsew signal output
flabel metal5 s 4892 0 5332 11844 0 FreeSans 2560 90 0 0 VGND
port 211 nsew ground bidirectional
flabel metal5 s 4892 0 5332 40 0 FreeSans 320 0 0 0 VGND
port 211 nsew ground bidirectional
flabel metal5 s 4892 11804 5332 11844 0 FreeSans 320 0 0 0 VGND
port 211 nsew ground bidirectional
flabel metal5 s 20012 0 20452 11844 0 FreeSans 2560 90 0 0 VGND
port 211 nsew ground bidirectional
flabel metal5 s 20012 0 20452 40 0 FreeSans 320 0 0 0 VGND
port 211 nsew ground bidirectional
flabel metal5 s 20012 11804 20452 11844 0 FreeSans 320 0 0 0 VGND
port 211 nsew ground bidirectional
flabel metal5 s 35132 0 35572 11844 0 FreeSans 2560 90 0 0 VGND
port 211 nsew ground bidirectional
flabel metal5 s 35132 0 35572 40 0 FreeSans 320 0 0 0 VGND
port 211 nsew ground bidirectional
flabel metal5 s 35132 11804 35572 11844 0 FreeSans 320 0 0 0 VGND
port 211 nsew ground bidirectional
flabel metal5 s 3652 0 4092 11844 0 FreeSans 2560 90 0 0 VPWR
port 212 nsew power bidirectional
flabel metal5 s 3652 0 4092 40 0 FreeSans 320 0 0 0 VPWR
port 212 nsew power bidirectional
flabel metal5 s 3652 11804 4092 11844 0 FreeSans 320 0 0 0 VPWR
port 212 nsew power bidirectional
flabel metal5 s 18772 0 19212 11844 0 FreeSans 2560 90 0 0 VPWR
port 212 nsew power bidirectional
flabel metal5 s 18772 0 19212 40 0 FreeSans 320 0 0 0 VPWR
port 212 nsew power bidirectional
flabel metal5 s 18772 11804 19212 11844 0 FreeSans 320 0 0 0 VPWR
port 212 nsew power bidirectional
flabel metal5 s 33892 0 34332 11844 0 FreeSans 2560 90 0 0 VPWR
port 212 nsew power bidirectional
flabel metal5 s 33892 0 34332 40 0 FreeSans 320 0 0 0 VPWR
port 212 nsew power bidirectional
flabel metal5 s 33892 11804 34332 11844 0 FreeSans 320 0 0 0 VPWR
port 212 nsew power bidirectional
rlabel metal1 23184 9072 23184 9072 0 VGND
rlabel metal1 23184 9828 23184 9828 0 VPWR
rlabel metal2 9344 588 9344 588 0 FrameData[0]
rlabel metal2 10112 3948 10112 3948 0 FrameData[10]
rlabel metal3 22944 3906 22944 3906 0 FrameData[11]
rlabel metal2 656 4620 656 4620 0 FrameData[12]
rlabel metal2 608 4956 608 4956 0 FrameData[13]
rlabel metal2 368 5292 368 5292 0 FrameData[14]
rlabel metal2 752 5628 752 5628 0 FrameData[15]
rlabel metal3 34464 5040 34464 5040 0 FrameData[16]
rlabel metal2 416 6300 416 6300 0 FrameData[17]
rlabel metal2 1472 6636 1472 6636 0 FrameData[18]
rlabel metal3 33312 6510 33312 6510 0 FrameData[19]
rlabel metal2 9296 924 9296 924 0 FrameData[1]
rlabel metal3 32736 7644 32736 7644 0 FrameData[20]
rlabel metal3 35712 7392 35712 7392 0 FrameData[21]
rlabel metal2 176 7980 176 7980 0 FrameData[22]
rlabel metal2 128 8316 128 8316 0 FrameData[23]
rlabel metal2 752 8652 752 8652 0 FrameData[24]
rlabel metal2 752 8988 752 8988 0 FrameData[25]
rlabel metal2 752 9324 752 9324 0 FrameData[26]
rlabel metal2 752 9660 752 9660 0 FrameData[27]
rlabel metal2 752 9996 752 9996 0 FrameData[28]
rlabel metal2 320 10332 320 10332 0 FrameData[29]
rlabel metal2 752 1260 752 1260 0 FrameData[2]
rlabel metal2 176 10668 176 10668 0 FrameData[30]
rlabel metal2 704 11004 704 11004 0 FrameData[31]
rlabel metal2 9392 1596 9392 1596 0 FrameData[3]
rlabel metal2 704 1932 704 1932 0 FrameData[4]
rlabel metal2 19296 3318 19296 3318 0 FrameData[5]
rlabel metal2 3632 2604 3632 2604 0 FrameData[6]
rlabel metal3 17280 3570 17280 3570 0 FrameData[7]
rlabel metal2 19200 3402 19200 3402 0 FrameData[8]
rlabel metal2 25920 3528 25920 3528 0 FrameData[9]
rlabel metal2 45471 588 45471 588 0 FrameData_O[0]
rlabel metal2 46047 3948 46047 3948 0 FrameData_O[10]
rlabel metal2 45735 4284 45735 4284 0 FrameData_O[11]
rlabel metal2 45951 4620 45951 4620 0 FrameData_O[12]
rlabel metal2 45735 4956 45735 4956 0 FrameData_O[13]
rlabel via2 46287 5292 46287 5292 0 FrameData_O[14]
rlabel metal2 45735 5628 45735 5628 0 FrameData_O[15]
rlabel via2 46287 5964 46287 5964 0 FrameData_O[16]
rlabel metal2 45735 6300 45735 6300 0 FrameData_O[17]
rlabel metal2 45663 6636 45663 6636 0 FrameData_O[18]
rlabel metal2 45735 6972 45735 6972 0 FrameData_O[19]
rlabel metal2 45999 924 45999 924 0 FrameData_O[1]
rlabel metal2 46047 7308 46047 7308 0 FrameData_O[20]
rlabel metal2 45543 7644 45543 7644 0 FrameData_O[21]
rlabel metal2 46047 7980 46047 7980 0 FrameData_O[22]
rlabel metal2 45543 8316 45543 8316 0 FrameData_O[23]
rlabel metal2 46047 8652 46047 8652 0 FrameData_O[24]
rlabel metal2 45951 8988 45951 8988 0 FrameData_O[25]
rlabel metal2 45351 9324 45351 9324 0 FrameData_O[26]
rlabel metal2 45159 9660 45159 9660 0 FrameData_O[27]
rlabel metal2 44424 8904 44424 8904 0 FrameData_O[28]
rlabel metal2 43656 9660 43656 9660 0 FrameData_O[29]
rlabel metal2 45663 1260 45663 1260 0 FrameData_O[2]
rlabel metal2 43320 9660 43320 9660 0 FrameData_O[30]
rlabel metal2 44088 8904 44088 8904 0 FrameData_O[31]
rlabel metal2 45663 1596 45663 1596 0 FrameData_O[3]
rlabel metal2 45663 1932 45663 1932 0 FrameData_O[4]
rlabel metal2 45480 2100 45480 2100 0 FrameData_O[5]
rlabel metal2 46047 2604 46047 2604 0 FrameData_O[6]
rlabel metal2 45336 2856 45336 2856 0 FrameData_O[7]
rlabel metal2 45543 3276 45543 3276 0 FrameData_O[8]
rlabel metal2 45735 3612 45735 3612 0 FrameData_O[9]
rlabel metal2 5952 6384 5952 6384 0 FrameStrobe[0]
rlabel metal2 27552 5292 27552 5292 0 FrameStrobe[10]
rlabel metal3 27312 420 27312 420 0 FrameStrobe[11]
rlabel metal3 29472 324 29472 324 0 FrameStrobe[12]
rlabel metal2 31104 5628 31104 5628 0 FrameStrobe[13]
rlabel metal3 33696 2466 33696 2466 0 FrameStrobe[14]
rlabel metal3 35808 2508 35808 2508 0 FrameStrobe[15]
rlabel metal2 33888 5460 33888 5460 0 FrameStrobe[16]
rlabel metal2 34464 5586 34464 5586 0 FrameStrobe[17]
rlabel metal2 37968 4788 37968 4788 0 FrameStrobe[18]
rlabel metal3 44256 2886 44256 2886 0 FrameStrobe[19]
rlabel metal2 6816 6468 6816 6468 0 FrameStrobe[1]
rlabel metal2 8448 4956 8448 4956 0 FrameStrobe[2]
rlabel metal3 10464 1332 10464 1332 0 FrameStrobe[3]
rlabel metal3 12576 1332 12576 1332 0 FrameStrobe[4]
rlabel metal3 14688 2046 14688 2046 0 FrameStrobe[5]
rlabel metal2 26112 4830 26112 4830 0 FrameStrobe[6]
rlabel metal3 18912 114 18912 114 0 FrameStrobe[7]
rlabel metal2 21984 4200 21984 4200 0 FrameStrobe[8]
rlabel metal3 23136 1470 23136 1470 0 FrameStrobe[9]
rlabel metal2 31512 9576 31512 9576 0 FrameStrobe_O[0]
rlabel metal2 33336 8904 33336 8904 0 FrameStrobe_O[10]
rlabel metal2 33960 9324 33960 9324 0 FrameStrobe_O[11]
rlabel metal2 34200 9660 34200 9660 0 FrameStrobe_O[12]
rlabel metal2 34776 9240 34776 9240 0 FrameStrobe_O[13]
rlabel metal2 35352 9240 35352 9240 0 FrameStrobe_O[14]
rlabel metal2 34632 8904 34632 8904 0 FrameStrobe_O[15]
rlabel metal2 35160 9324 35160 9324 0 FrameStrobe_O[16]
rlabel metal2 34968 8820 34968 8820 0 FrameStrobe_O[17]
rlabel metal2 36024 9660 36024 9660 0 FrameStrobe_O[18]
rlabel metal2 35832 9576 35832 9576 0 FrameStrobe_O[19]
rlabel metal2 31800 9660 31800 9660 0 FrameStrobe_O[1]
rlabel metal2 32088 9576 32088 9576 0 FrameStrobe_O[2]
rlabel metal2 32568 9660 32568 9660 0 FrameStrobe_O[3]
rlabel metal2 32184 8904 32184 8904 0 FrameStrobe_O[4]
rlabel metal2 33144 9660 33144 9660 0 FrameStrobe_O[5]
rlabel metal2 32568 8904 32568 8904 0 FrameStrobe_O[6]
rlabel metal2 33504 9534 33504 9534 0 FrameStrobe_O[7]
rlabel metal2 32952 8904 32952 8904 0 FrameStrobe_O[8]
rlabel metal2 33720 9240 33720 9240 0 FrameStrobe_O[9]
rlabel metal2 11064 8904 11064 8904 0 N1BEG[0]
rlabel metal2 11112 9660 11112 9660 0 N1BEG[1]
rlabel metal2 11448 8904 11448 8904 0 N1BEG[2]
rlabel metal2 11496 9660 11496 9660 0 N1BEG[3]
rlabel metal2 11832 8904 11832 8904 0 N2BEG[0]
rlabel metal2 11880 9660 11880 9660 0 N2BEG[1]
rlabel metal2 12216 8904 12216 8904 0 N2BEG[2]
rlabel metal2 12264 9660 12264 9660 0 N2BEG[3]
rlabel metal2 12600 8904 12600 8904 0 N2BEG[4]
rlabel metal2 12648 9660 12648 9660 0 N2BEG[5]
rlabel metal2 13032 8568 13032 8568 0 N2BEG[6]
rlabel metal3 13152 10722 13152 10722 0 N2BEG[7]
rlabel metal2 13368 8904 13368 8904 0 N2BEGb[0]
rlabel metal2 13416 9660 13416 9660 0 N2BEGb[1]
rlabel metal2 13752 8904 13752 8904 0 N2BEGb[2]
rlabel metal2 13800 9660 13800 9660 0 N2BEGb[3]
rlabel metal2 14136 8904 14136 8904 0 N2BEGb[4]
rlabel metal2 14184 9660 14184 9660 0 N2BEGb[5]
rlabel metal2 14520 8904 14520 8904 0 N2BEGb[6]
rlabel metal2 14568 9660 14568 9660 0 N2BEGb[7]
rlabel metal2 14904 8904 14904 8904 0 N4BEG[0]
rlabel metal2 16824 8904 16824 8904 0 N4BEG[10]
rlabel metal2 16872 9660 16872 9660 0 N4BEG[11]
rlabel metal2 17208 8904 17208 8904 0 N4BEG[12]
rlabel metal2 17256 9660 17256 9660 0 N4BEG[13]
rlabel metal2 17592 8904 17592 8904 0 N4BEG[14]
rlabel metal2 17640 9660 17640 9660 0 N4BEG[15]
rlabel metal2 14952 9660 14952 9660 0 N4BEG[1]
rlabel metal2 15288 8904 15288 8904 0 N4BEG[2]
rlabel metal2 15336 9660 15336 9660 0 N4BEG[3]
rlabel metal2 15672 8904 15672 8904 0 N4BEG[4]
rlabel metal2 15720 9660 15720 9660 0 N4BEG[5]
rlabel metal2 16056 8904 16056 8904 0 N4BEG[6]
rlabel metal2 16104 9660 16104 9660 0 N4BEG[7]
rlabel metal2 16440 8904 16440 8904 0 N4BEG[8]
rlabel metal2 16488 9660 16488 9660 0 N4BEG[9]
rlabel metal2 17976 8904 17976 8904 0 NN4BEG[0]
rlabel metal2 19896 8904 19896 8904 0 NN4BEG[10]
rlabel metal2 19848 9324 19848 9324 0 NN4BEG[11]
rlabel metal2 20232 9660 20232 9660 0 NN4BEG[12]
rlabel metal2 20376 9576 20376 9576 0 NN4BEG[13]
rlabel metal2 20664 9660 20664 9660 0 NN4BEG[14]
rlabel metal2 21288 9660 21288 9660 0 NN4BEG[15]
rlabel metal2 18024 9660 18024 9660 0 NN4BEG[1]
rlabel metal2 18360 8904 18360 8904 0 NN4BEG[2]
rlabel metal2 18408 9660 18408 9660 0 NN4BEG[3]
rlabel metal2 18744 8904 18744 8904 0 NN4BEG[4]
rlabel metal2 18648 9660 18648 9660 0 NN4BEG[5]
rlabel metal2 19224 8904 19224 8904 0 NN4BEG[6]
rlabel metal2 19224 9660 19224 9660 0 NN4BEG[7]
rlabel metal2 19512 8904 19512 8904 0 NN4BEG[8]
rlabel metal2 19560 9576 19560 9576 0 NN4BEG[9]
rlabel metal3 21216 9462 21216 9462 0 S1END[0]
rlabel metal3 21408 9294 21408 9294 0 S1END[1]
rlabel metal3 21600 9252 21600 9252 0 S1END[2]
rlabel metal3 21792 11394 21792 11394 0 S1END[3]
rlabel metal2 19296 6510 19296 6510 0 S2END[0]
rlabel metal3 19584 9492 19584 9492 0 S2END[1]
rlabel metal3 19968 10080 19968 10080 0 S2END[2]
rlabel metal3 15840 6342 15840 6342 0 S2END[3]
rlabel metal2 20544 4578 20544 4578 0 S2END[4]
rlabel metal3 16512 8526 16512 8526 0 S2END[5]
rlabel metal3 14976 6762 14976 6762 0 S2END[6]
rlabel metal3 13728 6762 13728 6762 0 S2END[7]
rlabel metal3 21984 11646 21984 11646 0 S2MID[0]
rlabel via2 22176 11772 22176 11772 0 S2MID[1]
rlabel metal3 22368 11730 22368 11730 0 S2MID[2]
rlabel metal3 22560 10134 22560 10134 0 S2MID[3]
rlabel metal3 22752 10008 22752 10008 0 S2MID[4]
rlabel metal3 22944 11730 22944 11730 0 S2MID[5]
rlabel metal3 16128 5838 16128 5838 0 S2MID[6]
rlabel metal3 13920 4788 13920 4788 0 S2MID[7]
rlabel metal2 19968 5376 19968 5376 0 S4END[0]
rlabel metal3 20064 5544 20064 5544 0 S4END[10]
rlabel metal2 21600 5544 21600 5544 0 S4END[11]
rlabel metal3 19584 4662 19584 4662 0 S4END[12]
rlabel metal3 21984 5964 21984 5964 0 S4END[13]
rlabel metal3 18528 6090 18528 6090 0 S4END[14]
rlabel metal3 18144 6048 18144 6048 0 S4END[15]
rlabel metal2 21792 5670 21792 5670 0 S4END[1]
rlabel metal2 21888 5754 21888 5754 0 S4END[2]
rlabel metal3 22368 4956 22368 4956 0 S4END[3]
rlabel metal2 21600 5040 21600 5040 0 S4END[4]
rlabel metal2 20064 6426 20064 6426 0 S4END[5]
rlabel metal4 20928 4788 20928 4788 0 S4END[6]
rlabel metal3 21600 5040 21600 5040 0 S4END[7]
rlabel metal3 26592 11394 26592 11394 0 S4END[8]
rlabel metal3 21216 5418 21216 5418 0 S4END[9]
rlabel metal3 28128 9882 28128 9882 0 SS4END[0]
rlabel metal3 30048 10848 30048 10848 0 SS4END[10]
rlabel metal3 30240 9672 30240 9672 0 SS4END[11]
rlabel metal3 30432 10092 30432 10092 0 SS4END[12]
rlabel metal3 30624 10470 30624 10470 0 SS4END[13]
rlabel metal3 30816 10428 30816 10428 0 SS4END[14]
rlabel metal3 31008 10386 31008 10386 0 SS4END[15]
rlabel metal3 28320 10302 28320 10302 0 SS4END[1]
rlabel metal3 28512 10218 28512 10218 0 SS4END[2]
rlabel metal3 28704 10260 28704 10260 0 SS4END[3]
rlabel metal3 28896 10344 28896 10344 0 SS4END[4]
rlabel metal3 29088 9840 29088 9840 0 SS4END[5]
rlabel metal4 28272 7980 28272 7980 0 SS4END[6]
rlabel metal3 29472 10050 29472 10050 0 SS4END[7]
rlabel metal3 29664 9462 29664 9462 0 SS4END[8]
rlabel metal3 29856 10134 29856 10134 0 SS4END[9]
rlabel metal3 2016 2844 2016 2844 0 UserCLK
rlabel metal2 31224 9660 31224 9660 0 UserCLKo
rlabel metal2 44160 1974 44160 1974 0 net1
rlabel metal3 44544 6636 44544 6636 0 net10
rlabel metal3 21696 9240 21696 9240 0 net100
rlabel metal2 21216 8694 21216 8694 0 net101
rlabel metal3 18720 7728 18720 7728 0 net102
rlabel metal3 20736 9156 20736 9156 0 net103
rlabel metal2 19488 9828 19488 9828 0 net104
rlabel metal2 17952 5460 17952 5460 0 net105
rlabel metal3 21024 10512 21024 10512 0 net106
rlabel metal2 44928 7098 44928 7098 0 net11
rlabel metal2 41280 1848 41280 1848 0 net12
rlabel metal2 44928 8022 44928 8022 0 net13
rlabel metal2 44064 7980 44064 7980 0 net14
rlabel metal2 44928 8820 44928 8820 0 net15
rlabel metal2 44544 8694 44544 8694 0 net16
rlabel metal2 44928 9534 44928 9534 0 net17
rlabel metal2 44256 9324 44256 9324 0 net18
rlabel metal2 44160 9408 44160 9408 0 net19
rlabel metal2 42432 4116 42432 4116 0 net2
rlabel metal3 43776 9198 43776 9198 0 net20
rlabel metal3 43968 9030 43968 9030 0 net21
rlabel metal3 43392 9156 43392 9156 0 net22
rlabel metal2 40992 1932 40992 1932 0 net23
rlabel metal2 43080 8148 43080 8148 0 net24
rlabel metal2 40152 8148 40152 8148 0 net25
rlabel metal2 44544 2058 44544 2058 0 net26
rlabel metal3 44160 2814 44160 2814 0 net27
rlabel metal3 44640 2562 44640 2562 0 net28
rlabel metal2 41712 2688 41712 2688 0 net29
rlabel metal2 44640 4074 44640 4074 0 net3
rlabel metal2 44928 2772 44928 2772 0 net30
rlabel metal2 44544 3654 44544 3654 0 net31
rlabel metal2 44928 3402 44928 3402 0 net32
rlabel metal3 31680 7896 31680 7896 0 net33
rlabel metal2 33312 8568 33312 8568 0 net34
rlabel metal3 34848 7266 34848 7266 0 net35
rlabel metal2 34368 9870 34368 9870 0 net36
rlabel metal2 34416 9408 34416 9408 0 net37
rlabel metal2 33600 10038 33600 10038 0 net38
rlabel metal3 34752 6888 34752 6888 0 net39
rlabel metal2 34152 2520 34152 2520 0 net4
rlabel metal2 33504 10122 33504 10122 0 net40
rlabel metal2 33336 5628 33336 5628 0 net41
rlabel metal2 34296 5628 34296 5628 0 net42
rlabel metal2 35256 5628 35256 5628 0 net43
rlabel metal2 7848 6636 7848 6636 0 net44
rlabel metal2 9984 4578 9984 4578 0 net45
rlabel metal2 17280 2268 17280 2268 0 net46
rlabel metal2 23592 2856 23592 2856 0 net47
rlabel metal2 33408 9324 33408 9324 0 net48
rlabel metal2 29592 4788 29592 4788 0 net49
rlabel metal2 44928 4914 44928 4914 0 net5
rlabel metal2 33600 9702 33600 9702 0 net50
rlabel metal2 24984 4284 24984 4284 0 net51
rlabel metal3 33216 7098 33216 7098 0 net52
rlabel metal2 9096 6552 9096 6552 0 net53
rlabel metal2 9480 6552 9480 6552 0 net54
rlabel metal2 8712 6552 8712 6552 0 net55
rlabel metal2 8616 7056 8616 7056 0 net56
rlabel metal2 11400 5544 11400 5544 0 net57
rlabel metal2 11352 5628 11352 5628 0 net58
rlabel metal2 12264 5544 12264 5544 0 net59
rlabel metal2 34536 2436 34536 2436 0 net6
rlabel metal2 11064 5460 11064 5460 0 net60
rlabel metal2 10536 5544 10536 5544 0 net61
rlabel metal2 10152 5544 10152 5544 0 net62
rlabel metal2 13104 8652 13104 8652 0 net63
rlabel metal2 10248 5124 10248 5124 0 net64
rlabel metal2 13608 5628 13608 5628 0 net65
rlabel metal2 13992 5460 13992 5460 0 net66
rlabel metal2 14184 5544 14184 5544 0 net67
rlabel metal2 15096 5628 15096 5628 0 net68
rlabel metal2 14328 5628 14328 5628 0 net69
rlabel metal3 43296 4578 43296 4578 0 net7
rlabel metal2 13896 5124 13896 5124 0 net70
rlabel metal2 13512 5544 13512 5544 0 net71
rlabel metal2 14088 6552 14088 6552 0 net72
rlabel metal2 17208 5628 17208 5628 0 net73
rlabel metal2 19752 6468 19752 6468 0 net74
rlabel metal2 19896 5040 19896 5040 0 net75
rlabel metal2 19128 5460 19128 5460 0 net76
rlabel metal2 20520 5460 20520 5460 0 net77
rlabel metal2 20232 5544 20232 5544 0 net78
rlabel metal2 19704 5460 19704 5460 0 net79
rlabel metal2 38232 4284 38232 4284 0 net8
rlabel metal2 18168 5796 18168 5796 0 net80
rlabel metal2 17352 6552 17352 6552 0 net81
rlabel metal2 17208 4788 17208 4788 0 net82
rlabel metal2 21336 5460 21336 5460 0 net83
rlabel metal2 18648 5796 18648 5796 0 net84
rlabel metal2 20856 5460 20856 5460 0 net85
rlabel metal2 17976 6216 17976 6216 0 net86
rlabel metal2 19944 5124 19944 5124 0 net87
rlabel metal2 18936 5796 18936 5796 0 net88
rlabel metal2 21504 9030 21504 9030 0 net89
rlabel metal3 44928 5838 44928 5838 0 net9
rlabel metal3 21696 8736 21696 8736 0 net90
rlabel metal2 19872 9660 19872 9660 0 net91
rlabel metal2 20448 9408 20448 9408 0 net92
rlabel metal2 20544 9450 20544 9450 0 net93
rlabel metal2 20928 9534 20928 9534 0 net94
rlabel metal2 27672 7728 27672 7728 0 net95
rlabel metal2 19392 9954 19392 9954 0 net96
rlabel metal2 21408 8904 21408 8904 0 net97
rlabel metal2 20544 10164 20544 10164 0 net98
rlabel metal2 21312 8778 21312 8778 0 net99
<< properties >>
string FIXED_BBOX 0 0 46368 11844
<< end >>
