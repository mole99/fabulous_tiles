module N_term_DSP (UserCLK,
    UserCLKo,
    FrameData,
    FrameData_O,
    FrameStrobe,
    FrameStrobe_O,
    N1END,
    N2END,
    N2MID,
    N4END,
    NN4END,
    S1BEG,
    S2BEG,
    S2BEGb,
    S4BEG,
    SS4BEG);
 input UserCLK;
 output UserCLKo;
 input [31:0] FrameData;
 output [31:0] FrameData_O;
 input [19:0] FrameStrobe;
 output [19:0] FrameStrobe_O;
 input [3:0] N1END;
 input [7:0] N2END;
 input [7:0] N2MID;
 input [15:0] N4END;
 input [15:0] NN4END;
 output [3:0] S1BEG;
 output [7:0] S2BEG;
 output [7:0] S2BEGb;
 output [15:0] S4BEG;
 output [15:0] SS4BEG;

 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;

 sg13g2_buf_1 _000_ (.A(FrameData[0]),
    .X(net1));
 sg13g2_buf_1 _001_ (.A(FrameData[1]),
    .X(net12));
 sg13g2_buf_1 _002_ (.A(FrameData[2]),
    .X(net23));
 sg13g2_buf_1 _003_ (.A(FrameData[3]),
    .X(net26));
 sg13g2_buf_1 _004_ (.A(FrameData[4]),
    .X(net27));
 sg13g2_buf_1 _005_ (.A(FrameData[5]),
    .X(net28));
 sg13g2_buf_1 _006_ (.A(FrameData[6]),
    .X(net29));
 sg13g2_buf_1 _007_ (.A(FrameData[7]),
    .X(net30));
 sg13g2_buf_1 _008_ (.A(FrameData[8]),
    .X(net31));
 sg13g2_buf_1 _009_ (.A(FrameData[9]),
    .X(net32));
 sg13g2_buf_1 _010_ (.A(FrameData[10]),
    .X(net2));
 sg13g2_buf_1 _011_ (.A(FrameData[11]),
    .X(net3));
 sg13g2_buf_1 _012_ (.A(FrameData[12]),
    .X(net4));
 sg13g2_buf_1 _013_ (.A(FrameData[13]),
    .X(net5));
 sg13g2_buf_1 _014_ (.A(FrameData[14]),
    .X(net6));
 sg13g2_buf_1 _015_ (.A(FrameData[15]),
    .X(net7));
 sg13g2_buf_1 _016_ (.A(FrameData[16]),
    .X(net8));
 sg13g2_buf_1 _017_ (.A(FrameData[17]),
    .X(net9));
 sg13g2_buf_1 _018_ (.A(FrameData[18]),
    .X(net10));
 sg13g2_buf_1 _019_ (.A(FrameData[19]),
    .X(net11));
 sg13g2_buf_1 _020_ (.A(FrameData[20]),
    .X(net13));
 sg13g2_buf_1 _021_ (.A(FrameData[21]),
    .X(net14));
 sg13g2_buf_1 _022_ (.A(FrameData[22]),
    .X(net15));
 sg13g2_buf_1 _023_ (.A(FrameData[23]),
    .X(net16));
 sg13g2_buf_1 _024_ (.A(FrameData[24]),
    .X(net17));
 sg13g2_buf_1 _025_ (.A(FrameData[25]),
    .X(net18));
 sg13g2_buf_1 _026_ (.A(FrameData[26]),
    .X(net19));
 sg13g2_buf_1 _027_ (.A(FrameData[27]),
    .X(net20));
 sg13g2_buf_1 _028_ (.A(FrameData[28]),
    .X(net21));
 sg13g2_buf_1 _029_ (.A(FrameData[29]),
    .X(net22));
 sg13g2_buf_1 _030_ (.A(FrameData[30]),
    .X(net24));
 sg13g2_buf_1 _031_ (.A(FrameData[31]),
    .X(net25));
 sg13g2_buf_1 _032_ (.A(FrameStrobe[0]),
    .X(net33));
 sg13g2_buf_1 _033_ (.A(FrameStrobe[1]),
    .X(net44));
 sg13g2_buf_1 _034_ (.A(FrameStrobe[2]),
    .X(net45));
 sg13g2_buf_1 _035_ (.A(FrameStrobe[3]),
    .X(net46));
 sg13g2_buf_1 _036_ (.A(FrameStrobe[4]),
    .X(net47));
 sg13g2_buf_1 _037_ (.A(FrameStrobe[5]),
    .X(net48));
 sg13g2_buf_1 _038_ (.A(FrameStrobe[6]),
    .X(net49));
 sg13g2_buf_1 _039_ (.A(FrameStrobe[7]),
    .X(net50));
 sg13g2_buf_1 _040_ (.A(FrameStrobe[8]),
    .X(net51));
 sg13g2_buf_1 _041_ (.A(FrameStrobe[9]),
    .X(net52));
 sg13g2_buf_1 _042_ (.A(FrameStrobe[10]),
    .X(net34));
 sg13g2_buf_1 _043_ (.A(FrameStrobe[11]),
    .X(net35));
 sg13g2_buf_1 _044_ (.A(FrameStrobe[12]),
    .X(net36));
 sg13g2_buf_1 _045_ (.A(FrameStrobe[13]),
    .X(net37));
 sg13g2_buf_1 _046_ (.A(FrameStrobe[14]),
    .X(net38));
 sg13g2_buf_1 _047_ (.A(FrameStrobe[15]),
    .X(net39));
 sg13g2_buf_1 _048_ (.A(FrameStrobe[16]),
    .X(net40));
 sg13g2_buf_1 _049_ (.A(FrameStrobe[17]),
    .X(net41));
 sg13g2_buf_1 _050_ (.A(FrameStrobe[18]),
    .X(net42));
 sg13g2_buf_1 _051_ (.A(FrameStrobe[19]),
    .X(net43));
 sg13g2_buf_1 _052_ (.A(N1END[3]),
    .X(net53));
 sg13g2_buf_1 _053_ (.A(N1END[2]),
    .X(net54));
 sg13g2_buf_1 _054_ (.A(N1END[1]),
    .X(net55));
 sg13g2_buf_1 _055_ (.A(N1END[0]),
    .X(net56));
 sg13g2_buf_1 _056_ (.A(N2MID[7]),
    .X(net57));
 sg13g2_buf_1 _057_ (.A(N2MID[6]),
    .X(net58));
 sg13g2_buf_1 _058_ (.A(N2MID[5]),
    .X(net59));
 sg13g2_buf_1 _059_ (.A(N2MID[4]),
    .X(net60));
 sg13g2_buf_1 _060_ (.A(N2MID[3]),
    .X(net61));
 sg13g2_buf_1 _061_ (.A(N2MID[2]),
    .X(net62));
 sg13g2_buf_1 _062_ (.A(N2MID[1]),
    .X(net63));
 sg13g2_buf_1 _063_ (.A(N2MID[0]),
    .X(net64));
 sg13g2_buf_1 _064_ (.A(N2END[7]),
    .X(net65));
 sg13g2_buf_1 _065_ (.A(N2END[6]),
    .X(net66));
 sg13g2_buf_1 _066_ (.A(N2END[5]),
    .X(net67));
 sg13g2_buf_1 _067_ (.A(N2END[4]),
    .X(net68));
 sg13g2_buf_1 _068_ (.A(N2END[3]),
    .X(net69));
 sg13g2_buf_1 _069_ (.A(N2END[2]),
    .X(net70));
 sg13g2_buf_1 _070_ (.A(N2END[1]),
    .X(net71));
 sg13g2_buf_1 _071_ (.A(N2END[0]),
    .X(net72));
 sg13g2_buf_1 _072_ (.A(N4END[15]),
    .X(net73));
 sg13g2_buf_1 _073_ (.A(N4END[14]),
    .X(net80));
 sg13g2_buf_1 _074_ (.A(N4END[13]),
    .X(net81));
 sg13g2_buf_1 _075_ (.A(N4END[12]),
    .X(net82));
 sg13g2_buf_1 _076_ (.A(N4END[11]),
    .X(net83));
 sg13g2_buf_1 _077_ (.A(N4END[10]),
    .X(net84));
 sg13g2_buf_1 _078_ (.A(N4END[9]),
    .X(net85));
 sg13g2_buf_1 _079_ (.A(N4END[8]),
    .X(net86));
 sg13g2_buf_1 _080_ (.A(N4END[7]),
    .X(net87));
 sg13g2_buf_1 _081_ (.A(N4END[6]),
    .X(net88));
 sg13g2_buf_1 _082_ (.A(N4END[5]),
    .X(net74));
 sg13g2_buf_1 _083_ (.A(N4END[4]),
    .X(net75));
 sg13g2_buf_1 _084_ (.A(N4END[3]),
    .X(net76));
 sg13g2_buf_1 _085_ (.A(N4END[2]),
    .X(net77));
 sg13g2_buf_1 _086_ (.A(N4END[1]),
    .X(net78));
 sg13g2_buf_1 _087_ (.A(N4END[0]),
    .X(net79));
 sg13g2_buf_1 _088_ (.A(NN4END[15]),
    .X(net89));
 sg13g2_buf_1 _089_ (.A(NN4END[14]),
    .X(net96));
 sg13g2_buf_1 _090_ (.A(NN4END[13]),
    .X(net97));
 sg13g2_buf_1 _091_ (.A(NN4END[12]),
    .X(net98));
 sg13g2_buf_1 _092_ (.A(NN4END[11]),
    .X(net99));
 sg13g2_buf_1 _093_ (.A(NN4END[10]),
    .X(net100));
 sg13g2_buf_1 _094_ (.A(NN4END[9]),
    .X(net101));
 sg13g2_buf_1 _095_ (.A(NN4END[8]),
    .X(net102));
 sg13g2_buf_1 _096_ (.A(NN4END[7]),
    .X(net103));
 sg13g2_buf_1 _097_ (.A(NN4END[6]),
    .X(net104));
 sg13g2_buf_1 _098_ (.A(NN4END[5]),
    .X(net90));
 sg13g2_buf_1 _099_ (.A(NN4END[4]),
    .X(net91));
 sg13g2_buf_1 _100_ (.A(NN4END[3]),
    .X(net92));
 sg13g2_buf_1 _101_ (.A(NN4END[2]),
    .X(net93));
 sg13g2_buf_1 _102_ (.A(NN4END[1]),
    .X(net94));
 sg13g2_buf_1 _103_ (.A(NN4END[0]),
    .X(net95));
 sg13g2_buf_1 _104_ (.A(UserCLK),
    .X(net105));
 sg13g2_buf_1 output1 (.A(net1),
    .X(FrameData_O[0]));
 sg13g2_buf_1 output2 (.A(net2),
    .X(FrameData_O[10]));
 sg13g2_buf_1 output3 (.A(net3),
    .X(FrameData_O[11]));
 sg13g2_buf_1 output4 (.A(net4),
    .X(FrameData_O[12]));
 sg13g2_buf_1 output5 (.A(net5),
    .X(FrameData_O[13]));
 sg13g2_buf_1 output6 (.A(net6),
    .X(FrameData_O[14]));
 sg13g2_buf_1 output7 (.A(net7),
    .X(FrameData_O[15]));
 sg13g2_buf_1 output8 (.A(net8),
    .X(FrameData_O[16]));
 sg13g2_buf_1 output9 (.A(net9),
    .X(FrameData_O[17]));
 sg13g2_buf_1 output10 (.A(net10),
    .X(FrameData_O[18]));
 sg13g2_buf_1 output11 (.A(net11),
    .X(FrameData_O[19]));
 sg13g2_buf_1 output12 (.A(net12),
    .X(FrameData_O[1]));
 sg13g2_buf_1 output13 (.A(net13),
    .X(FrameData_O[20]));
 sg13g2_buf_1 output14 (.A(net14),
    .X(FrameData_O[21]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(FrameData_O[22]));
 sg13g2_buf_1 output16 (.A(net16),
    .X(FrameData_O[23]));
 sg13g2_buf_1 output17 (.A(net17),
    .X(FrameData_O[24]));
 sg13g2_buf_1 output18 (.A(net18),
    .X(FrameData_O[25]));
 sg13g2_buf_1 output19 (.A(net19),
    .X(FrameData_O[26]));
 sg13g2_buf_1 output20 (.A(net20),
    .X(FrameData_O[27]));
 sg13g2_buf_1 output21 (.A(net21),
    .X(FrameData_O[28]));
 sg13g2_buf_1 output22 (.A(net22),
    .X(FrameData_O[29]));
 sg13g2_buf_1 output23 (.A(net23),
    .X(FrameData_O[2]));
 sg13g2_buf_1 output24 (.A(net24),
    .X(FrameData_O[30]));
 sg13g2_buf_1 output25 (.A(net25),
    .X(FrameData_O[31]));
 sg13g2_buf_1 output26 (.A(net26),
    .X(FrameData_O[3]));
 sg13g2_buf_1 output27 (.A(net27),
    .X(FrameData_O[4]));
 sg13g2_buf_1 output28 (.A(net28),
    .X(FrameData_O[5]));
 sg13g2_buf_1 output29 (.A(net29),
    .X(FrameData_O[6]));
 sg13g2_buf_1 output30 (.A(net30),
    .X(FrameData_O[7]));
 sg13g2_buf_1 output31 (.A(net31),
    .X(FrameData_O[8]));
 sg13g2_buf_1 output32 (.A(net32),
    .X(FrameData_O[9]));
 sg13g2_buf_1 output33 (.A(net33),
    .X(FrameStrobe_O[0]));
 sg13g2_buf_1 output34 (.A(net34),
    .X(FrameStrobe_O[10]));
 sg13g2_buf_1 output35 (.A(net35),
    .X(FrameStrobe_O[11]));
 sg13g2_buf_1 output36 (.A(net36),
    .X(FrameStrobe_O[12]));
 sg13g2_buf_1 output37 (.A(net37),
    .X(FrameStrobe_O[13]));
 sg13g2_buf_1 output38 (.A(net38),
    .X(FrameStrobe_O[14]));
 sg13g2_buf_1 output39 (.A(net39),
    .X(FrameStrobe_O[15]));
 sg13g2_buf_1 output40 (.A(net40),
    .X(FrameStrobe_O[16]));
 sg13g2_buf_1 output41 (.A(net41),
    .X(FrameStrobe_O[17]));
 sg13g2_buf_1 output42 (.A(net42),
    .X(FrameStrobe_O[18]));
 sg13g2_buf_1 output43 (.A(net43),
    .X(FrameStrobe_O[19]));
 sg13g2_buf_1 output44 (.A(net44),
    .X(FrameStrobe_O[1]));
 sg13g2_buf_1 output45 (.A(net45),
    .X(FrameStrobe_O[2]));
 sg13g2_buf_1 output46 (.A(net46),
    .X(FrameStrobe_O[3]));
 sg13g2_buf_1 output47 (.A(net47),
    .X(FrameStrobe_O[4]));
 sg13g2_buf_1 output48 (.A(net48),
    .X(FrameStrobe_O[5]));
 sg13g2_buf_1 output49 (.A(net49),
    .X(FrameStrobe_O[6]));
 sg13g2_buf_1 output50 (.A(net50),
    .X(FrameStrobe_O[7]));
 sg13g2_buf_1 output51 (.A(net51),
    .X(FrameStrobe_O[8]));
 sg13g2_buf_1 output52 (.A(net52),
    .X(FrameStrobe_O[9]));
 sg13g2_buf_1 output53 (.A(net53),
    .X(S1BEG[0]));
 sg13g2_buf_1 output54 (.A(net54),
    .X(S1BEG[1]));
 sg13g2_buf_1 output55 (.A(net55),
    .X(S1BEG[2]));
 sg13g2_buf_1 output56 (.A(net56),
    .X(S1BEG[3]));
 sg13g2_buf_1 output57 (.A(net57),
    .X(S2BEG[0]));
 sg13g2_buf_1 output58 (.A(net58),
    .X(S2BEG[1]));
 sg13g2_buf_1 output59 (.A(net59),
    .X(S2BEG[2]));
 sg13g2_buf_1 output60 (.A(net60),
    .X(S2BEG[3]));
 sg13g2_buf_1 output61 (.A(net61),
    .X(S2BEG[4]));
 sg13g2_buf_1 output62 (.A(net62),
    .X(S2BEG[5]));
 sg13g2_buf_1 output63 (.A(net63),
    .X(S2BEG[6]));
 sg13g2_buf_1 output64 (.A(net64),
    .X(S2BEG[7]));
 sg13g2_buf_1 output65 (.A(net65),
    .X(S2BEGb[0]));
 sg13g2_buf_1 output66 (.A(net66),
    .X(S2BEGb[1]));
 sg13g2_buf_1 output67 (.A(net67),
    .X(S2BEGb[2]));
 sg13g2_buf_1 output68 (.A(net68),
    .X(S2BEGb[3]));
 sg13g2_buf_1 output69 (.A(net69),
    .X(S2BEGb[4]));
 sg13g2_buf_1 output70 (.A(net70),
    .X(S2BEGb[5]));
 sg13g2_buf_1 output71 (.A(net71),
    .X(S2BEGb[6]));
 sg13g2_buf_1 output72 (.A(net72),
    .X(S2BEGb[7]));
 sg13g2_buf_1 output73 (.A(net73),
    .X(S4BEG[0]));
 sg13g2_buf_1 output74 (.A(net74),
    .X(S4BEG[10]));
 sg13g2_buf_1 output75 (.A(net75),
    .X(S4BEG[11]));
 sg13g2_buf_1 output76 (.A(net76),
    .X(S4BEG[12]));
 sg13g2_buf_1 output77 (.A(net77),
    .X(S4BEG[13]));
 sg13g2_buf_1 output78 (.A(net78),
    .X(S4BEG[14]));
 sg13g2_buf_1 output79 (.A(net79),
    .X(S4BEG[15]));
 sg13g2_buf_1 output80 (.A(net80),
    .X(S4BEG[1]));
 sg13g2_buf_1 output81 (.A(net81),
    .X(S4BEG[2]));
 sg13g2_buf_1 output82 (.A(net82),
    .X(S4BEG[3]));
 sg13g2_buf_1 output83 (.A(net83),
    .X(S4BEG[4]));
 sg13g2_buf_1 output84 (.A(net84),
    .X(S4BEG[5]));
 sg13g2_buf_1 output85 (.A(net85),
    .X(S4BEG[6]));
 sg13g2_buf_1 output86 (.A(net86),
    .X(S4BEG[7]));
 sg13g2_buf_1 output87 (.A(net87),
    .X(S4BEG[8]));
 sg13g2_buf_1 output88 (.A(net88),
    .X(S4BEG[9]));
 sg13g2_buf_1 output89 (.A(net89),
    .X(SS4BEG[0]));
 sg13g2_buf_1 output90 (.A(net90),
    .X(SS4BEG[10]));
 sg13g2_buf_1 output91 (.A(net91),
    .X(SS4BEG[11]));
 sg13g2_buf_1 output92 (.A(net92),
    .X(SS4BEG[12]));
 sg13g2_buf_1 output93 (.A(net93),
    .X(SS4BEG[13]));
 sg13g2_buf_1 output94 (.A(net94),
    .X(SS4BEG[14]));
 sg13g2_buf_1 output95 (.A(net95),
    .X(SS4BEG[15]));
 sg13g2_buf_1 output96 (.A(net96),
    .X(SS4BEG[1]));
 sg13g2_buf_1 output97 (.A(net97),
    .X(SS4BEG[2]));
 sg13g2_buf_1 output98 (.A(net98),
    .X(SS4BEG[3]));
 sg13g2_buf_1 output99 (.A(net99),
    .X(SS4BEG[4]));
 sg13g2_buf_1 output100 (.A(net100),
    .X(SS4BEG[5]));
 sg13g2_buf_1 output101 (.A(net101),
    .X(SS4BEG[6]));
 sg13g2_buf_1 output102 (.A(net102),
    .X(SS4BEG[7]));
 sg13g2_buf_1 output103 (.A(net103),
    .X(SS4BEG[8]));
 sg13g2_buf_1 output104 (.A(net104),
    .X(SS4BEG[9]));
 sg13g2_buf_1 output105 (.A(net105),
    .X(UserCLKo));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_4 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_285 ();
 sg13g2_decap_8 FILLER_0_292 ();
 sg13g2_decap_8 FILLER_0_299 ();
 sg13g2_decap_8 FILLER_0_306 ();
 sg13g2_decap_8 FILLER_0_313 ();
 sg13g2_decap_8 FILLER_0_320 ();
 sg13g2_decap_8 FILLER_0_327 ();
 sg13g2_decap_8 FILLER_0_334 ();
 sg13g2_decap_8 FILLER_0_341 ();
 sg13g2_decap_8 FILLER_0_348 ();
 sg13g2_decap_8 FILLER_0_355 ();
 sg13g2_decap_8 FILLER_0_362 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_4 FILLER_1_168 ();
 sg13g2_fill_1 FILLER_1_172 ();
 sg13g2_decap_8 FILLER_1_197 ();
 sg13g2_decap_8 FILLER_1_204 ();
 sg13g2_decap_8 FILLER_1_275 ();
 sg13g2_decap_8 FILLER_1_282 ();
 sg13g2_decap_8 FILLER_1_289 ();
 sg13g2_decap_8 FILLER_1_296 ();
 sg13g2_decap_8 FILLER_1_303 ();
 sg13g2_decap_8 FILLER_1_310 ();
 sg13g2_decap_8 FILLER_1_317 ();
 sg13g2_decap_8 FILLER_1_324 ();
 sg13g2_decap_8 FILLER_1_331 ();
 sg13g2_decap_8 FILLER_1_338 ();
 sg13g2_decap_8 FILLER_1_345 ();
 sg13g2_decap_8 FILLER_1_352 ();
 sg13g2_decap_8 FILLER_1_359 ();
 sg13g2_decap_8 FILLER_1_366 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_4 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_131 ();
 sg13g2_decap_8 FILLER_2_138 ();
 sg13g2_decap_8 FILLER_2_145 ();
 sg13g2_decap_8 FILLER_2_152 ();
 sg13g2_decap_8 FILLER_2_159 ();
 sg13g2_decap_4 FILLER_2_166 ();
 sg13g2_fill_2 FILLER_2_170 ();
 sg13g2_decap_8 FILLER_2_180 ();
 sg13g2_decap_8 FILLER_2_187 ();
 sg13g2_decap_8 FILLER_2_194 ();
 sg13g2_decap_8 FILLER_2_201 ();
 sg13g2_decap_8 FILLER_2_208 ();
 sg13g2_decap_8 FILLER_2_223 ();
 sg13g2_decap_8 FILLER_2_230 ();
 sg13g2_decap_8 FILLER_2_237 ();
 sg13g2_decap_8 FILLER_2_244 ();
 sg13g2_decap_8 FILLER_2_251 ();
 sg13g2_decap_8 FILLER_2_258 ();
 sg13g2_decap_8 FILLER_2_265 ();
 sg13g2_fill_2 FILLER_2_272 ();
 sg13g2_fill_1 FILLER_2_274 ();
 sg13g2_decap_8 FILLER_2_279 ();
 sg13g2_fill_2 FILLER_2_286 ();
 sg13g2_fill_1 FILLER_2_288 ();
 sg13g2_decap_8 FILLER_2_293 ();
 sg13g2_decap_8 FILLER_2_300 ();
 sg13g2_fill_2 FILLER_2_307 ();
 sg13g2_decap_4 FILLER_2_313 ();
 sg13g2_fill_1 FILLER_2_317 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_4 FILLER_2_371 ();
 sg13g2_fill_2 FILLER_2_375 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_fill_2 FILLER_3_70 ();
 sg13g2_fill_1 FILLER_3_72 ();
 sg13g2_decap_8 FILLER_3_81 ();
 sg13g2_fill_2 FILLER_3_88 ();
 sg13g2_fill_1 FILLER_3_90 ();
 sg13g2_decap_8 FILLER_3_99 ();
 sg13g2_decap_4 FILLER_3_106 ();
 sg13g2_fill_1 FILLER_3_110 ();
 sg13g2_fill_2 FILLER_3_135 ();
 sg13g2_decap_8 FILLER_3_141 ();
 sg13g2_decap_8 FILLER_3_148 ();
 sg13g2_fill_2 FILLER_3_191 ();
 sg13g2_decap_8 FILLER_3_197 ();
 sg13g2_fill_2 FILLER_3_204 ();
 sg13g2_fill_1 FILLER_3_206 ();
 sg13g2_decap_8 FILLER_3_243 ();
 sg13g2_decap_8 FILLER_3_250 ();
 sg13g2_decap_8 FILLER_3_261 ();
 sg13g2_fill_2 FILLER_3_268 ();
 sg13g2_fill_1 FILLER_3_270 ();
 sg13g2_decap_8 FILLER_3_275 ();
 sg13g2_fill_1 FILLER_3_282 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_298 ();
 sg13g2_decap_8 FILLER_3_305 ();
 sg13g2_decap_4 FILLER_3_312 ();
 sg13g2_fill_2 FILLER_3_320 ();
 sg13g2_fill_1 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_335 ();
 sg13g2_decap_8 FILLER_3_342 ();
 sg13g2_decap_8 FILLER_3_349 ();
 sg13g2_decap_8 FILLER_3_356 ();
 sg13g2_decap_8 FILLER_3_363 ();
 sg13g2_fill_2 FILLER_3_370 ();
 sg13g2_fill_1 FILLER_3_372 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_fill_1 FILLER_4_71 ();
 sg13g2_fill_1 FILLER_4_88 ();
 sg13g2_decap_8 FILLER_4_97 ();
 sg13g2_decap_8 FILLER_4_104 ();
 sg13g2_decap_8 FILLER_4_111 ();
 sg13g2_decap_4 FILLER_4_118 ();
 sg13g2_fill_2 FILLER_4_122 ();
 sg13g2_decap_8 FILLER_4_128 ();
 sg13g2_decap_8 FILLER_4_135 ();
 sg13g2_decap_8 FILLER_4_142 ();
 sg13g2_decap_4 FILLER_4_149 ();
 sg13g2_fill_1 FILLER_4_153 ();
 sg13g2_decap_8 FILLER_4_158 ();
 sg13g2_fill_2 FILLER_4_169 ();
 sg13g2_decap_8 FILLER_4_179 ();
 sg13g2_decap_8 FILLER_4_186 ();
 sg13g2_decap_8 FILLER_4_193 ();
 sg13g2_decap_8 FILLER_4_200 ();
 sg13g2_decap_8 FILLER_4_207 ();
 sg13g2_fill_2 FILLER_4_214 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_fill_2 FILLER_4_252 ();
 sg13g2_fill_1 FILLER_4_254 ();
 sg13g2_fill_1 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_264 ();
 sg13g2_decap_8 FILLER_4_271 ();
 sg13g2_decap_8 FILLER_4_282 ();
 sg13g2_decap_8 FILLER_4_289 ();
 sg13g2_decap_8 FILLER_4_296 ();
 sg13g2_decap_8 FILLER_4_303 ();
 sg13g2_fill_2 FILLER_4_310 ();
 sg13g2_fill_1 FILLER_4_312 ();
 sg13g2_decap_8 FILLER_4_317 ();
 sg13g2_decap_8 FILLER_4_324 ();
 sg13g2_decap_4 FILLER_4_331 ();
 sg13g2_decap_8 FILLER_4_339 ();
 sg13g2_decap_8 FILLER_4_346 ();
 sg13g2_decap_8 FILLER_4_353 ();
 sg13g2_decap_8 FILLER_4_360 ();
 sg13g2_decap_8 FILLER_4_367 ();
 sg13g2_fill_2 FILLER_4_374 ();
 sg13g2_fill_1 FILLER_4_376 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_fill_1 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_19 ();
 sg13g2_decap_8 FILLER_5_26 ();
 sg13g2_decap_8 FILLER_5_33 ();
 sg13g2_decap_8 FILLER_5_40 ();
 sg13g2_decap_8 FILLER_5_47 ();
 sg13g2_decap_8 FILLER_5_54 ();
 sg13g2_decap_8 FILLER_5_61 ();
 sg13g2_decap_8 FILLER_5_68 ();
 sg13g2_decap_8 FILLER_5_75 ();
 sg13g2_decap_8 FILLER_5_82 ();
 sg13g2_decap_8 FILLER_5_89 ();
 sg13g2_decap_8 FILLER_5_96 ();
 sg13g2_decap_8 FILLER_5_103 ();
 sg13g2_decap_8 FILLER_5_110 ();
 sg13g2_decap_8 FILLER_5_117 ();
 sg13g2_decap_8 FILLER_5_124 ();
 sg13g2_decap_8 FILLER_5_131 ();
 sg13g2_decap_8 FILLER_5_138 ();
 sg13g2_decap_8 FILLER_5_145 ();
 sg13g2_decap_8 FILLER_5_152 ();
 sg13g2_decap_8 FILLER_5_159 ();
 sg13g2_decap_8 FILLER_5_166 ();
 sg13g2_decap_8 FILLER_5_173 ();
 sg13g2_decap_8 FILLER_5_180 ();
 sg13g2_decap_8 FILLER_5_187 ();
 sg13g2_decap_8 FILLER_5_194 ();
 sg13g2_decap_8 FILLER_5_201 ();
 sg13g2_decap_8 FILLER_5_208 ();
 sg13g2_decap_8 FILLER_5_215 ();
 sg13g2_decap_8 FILLER_5_222 ();
 sg13g2_decap_8 FILLER_5_229 ();
 sg13g2_decap_8 FILLER_5_236 ();
 sg13g2_decap_8 FILLER_5_243 ();
 sg13g2_decap_8 FILLER_5_250 ();
 sg13g2_decap_8 FILLER_5_257 ();
 sg13g2_decap_8 FILLER_5_264 ();
 sg13g2_decap_8 FILLER_5_271 ();
 sg13g2_decap_8 FILLER_5_278 ();
 sg13g2_decap_8 FILLER_5_285 ();
 sg13g2_decap_8 FILLER_5_292 ();
 sg13g2_decap_8 FILLER_5_299 ();
 sg13g2_decap_8 FILLER_5_306 ();
 sg13g2_decap_8 FILLER_5_313 ();
 sg13g2_decap_8 FILLER_5_320 ();
 sg13g2_decap_8 FILLER_5_327 ();
 sg13g2_decap_8 FILLER_5_334 ();
 sg13g2_decap_8 FILLER_5_341 ();
 sg13g2_decap_8 FILLER_5_348 ();
 sg13g2_decap_8 FILLER_5_355 ();
 sg13g2_decap_8 FILLER_5_362 ();
 sg13g2_decap_8 FILLER_5_369 ();
 sg13g2_fill_1 FILLER_5_376 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_fill_1 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_19 ();
 sg13g2_decap_8 FILLER_6_26 ();
 sg13g2_decap_8 FILLER_6_33 ();
 sg13g2_decap_8 FILLER_6_40 ();
 sg13g2_decap_8 FILLER_6_47 ();
 sg13g2_decap_8 FILLER_6_54 ();
 sg13g2_decap_8 FILLER_6_61 ();
 sg13g2_decap_8 FILLER_6_68 ();
 sg13g2_decap_8 FILLER_6_75 ();
 sg13g2_decap_8 FILLER_6_82 ();
 sg13g2_decap_8 FILLER_6_89 ();
 sg13g2_decap_8 FILLER_6_96 ();
 sg13g2_decap_8 FILLER_6_103 ();
 sg13g2_decap_8 FILLER_6_110 ();
 sg13g2_decap_8 FILLER_6_117 ();
 sg13g2_decap_8 FILLER_6_124 ();
 sg13g2_decap_8 FILLER_6_131 ();
 sg13g2_decap_8 FILLER_6_138 ();
 sg13g2_decap_8 FILLER_6_145 ();
 sg13g2_decap_8 FILLER_6_152 ();
 sg13g2_decap_8 FILLER_6_159 ();
 sg13g2_decap_8 FILLER_6_166 ();
 sg13g2_decap_8 FILLER_6_173 ();
 sg13g2_decap_8 FILLER_6_180 ();
 sg13g2_decap_8 FILLER_6_187 ();
 sg13g2_decap_8 FILLER_6_194 ();
 sg13g2_decap_8 FILLER_6_201 ();
 sg13g2_decap_8 FILLER_6_208 ();
 sg13g2_decap_8 FILLER_6_215 ();
 sg13g2_decap_8 FILLER_6_222 ();
 sg13g2_decap_8 FILLER_6_229 ();
 sg13g2_decap_8 FILLER_6_236 ();
 sg13g2_decap_8 FILLER_6_243 ();
 sg13g2_decap_8 FILLER_6_250 ();
 sg13g2_decap_8 FILLER_6_257 ();
 sg13g2_decap_8 FILLER_6_264 ();
 sg13g2_fill_2 FILLER_6_271 ();
 sg13g2_fill_1 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_278 ();
 sg13g2_decap_8 FILLER_6_285 ();
 sg13g2_decap_8 FILLER_6_292 ();
 sg13g2_decap_8 FILLER_6_299 ();
 sg13g2_decap_8 FILLER_6_306 ();
 sg13g2_fill_2 FILLER_6_313 ();
 sg13g2_decap_8 FILLER_6_319 ();
 sg13g2_decap_8 FILLER_6_326 ();
 sg13g2_decap_8 FILLER_6_333 ();
 sg13g2_decap_8 FILLER_6_340 ();
 sg13g2_decap_8 FILLER_6_347 ();
 sg13g2_decap_8 FILLER_6_354 ();
 sg13g2_decap_8 FILLER_6_361 ();
 sg13g2_decap_8 FILLER_6_368 ();
 sg13g2_fill_2 FILLER_6_375 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_4 FILLER_7_42 ();
 sg13g2_fill_2 FILLER_7_46 ();
 sg13g2_decap_8 FILLER_7_52 ();
 sg13g2_decap_8 FILLER_7_59 ();
 sg13g2_decap_8 FILLER_7_66 ();
 sg13g2_decap_8 FILLER_7_73 ();
 sg13g2_decap_8 FILLER_7_80 ();
 sg13g2_decap_8 FILLER_7_87 ();
 sg13g2_decap_8 FILLER_7_94 ();
 sg13g2_decap_8 FILLER_7_101 ();
 sg13g2_decap_8 FILLER_7_108 ();
 sg13g2_decap_8 FILLER_7_115 ();
 sg13g2_decap_8 FILLER_7_122 ();
 sg13g2_decap_8 FILLER_7_129 ();
 sg13g2_decap_8 FILLER_7_136 ();
 sg13g2_decap_8 FILLER_7_143 ();
 sg13g2_decap_8 FILLER_7_150 ();
 sg13g2_decap_8 FILLER_7_157 ();
 sg13g2_decap_8 FILLER_7_164 ();
 sg13g2_decap_8 FILLER_7_171 ();
 sg13g2_decap_8 FILLER_7_178 ();
 sg13g2_decap_8 FILLER_7_185 ();
 sg13g2_decap_8 FILLER_7_192 ();
 sg13g2_decap_8 FILLER_7_199 ();
 sg13g2_decap_8 FILLER_7_206 ();
 sg13g2_decap_8 FILLER_7_213 ();
 sg13g2_decap_8 FILLER_7_220 ();
 sg13g2_decap_8 FILLER_7_227 ();
 sg13g2_decap_8 FILLER_7_234 ();
 sg13g2_decap_8 FILLER_7_241 ();
 sg13g2_decap_8 FILLER_7_248 ();
 sg13g2_decap_8 FILLER_7_255 ();
 sg13g2_decap_8 FILLER_7_262 ();
 sg13g2_decap_8 FILLER_7_269 ();
 sg13g2_decap_8 FILLER_7_276 ();
 sg13g2_decap_8 FILLER_7_283 ();
 sg13g2_decap_8 FILLER_7_290 ();
 sg13g2_decap_8 FILLER_7_297 ();
 sg13g2_decap_8 FILLER_7_304 ();
 sg13g2_decap_8 FILLER_7_311 ();
 sg13g2_decap_8 FILLER_7_318 ();
 sg13g2_decap_8 FILLER_7_325 ();
 sg13g2_decap_8 FILLER_7_332 ();
 sg13g2_decap_8 FILLER_7_339 ();
 sg13g2_decap_8 FILLER_7_346 ();
 sg13g2_decap_8 FILLER_7_353 ();
 sg13g2_decap_8 FILLER_7_360 ();
 sg13g2_decap_8 FILLER_7_367 ();
 sg13g2_fill_2 FILLER_7_374 ();
 sg13g2_fill_1 FILLER_7_376 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_4 FILLER_8_91 ();
 sg13g2_fill_1 FILLER_8_95 ();
 sg13g2_fill_2 FILLER_8_100 ();
 sg13g2_fill_1 FILLER_8_102 ();
 sg13g2_decap_8 FILLER_8_111 ();
 sg13g2_decap_8 FILLER_8_118 ();
 sg13g2_decap_8 FILLER_8_125 ();
 sg13g2_decap_8 FILLER_8_132 ();
 sg13g2_decap_8 FILLER_8_139 ();
 sg13g2_decap_8 FILLER_8_146 ();
 sg13g2_decap_8 FILLER_8_153 ();
 sg13g2_decap_8 FILLER_8_160 ();
 sg13g2_decap_8 FILLER_8_167 ();
 sg13g2_decap_8 FILLER_8_174 ();
 sg13g2_decap_8 FILLER_8_181 ();
 sg13g2_decap_8 FILLER_8_188 ();
 sg13g2_decap_8 FILLER_8_195 ();
 sg13g2_decap_8 FILLER_8_202 ();
 sg13g2_decap_8 FILLER_8_209 ();
 sg13g2_decap_8 FILLER_8_216 ();
 sg13g2_decap_8 FILLER_8_223 ();
 sg13g2_decap_8 FILLER_8_230 ();
 sg13g2_decap_8 FILLER_8_237 ();
 sg13g2_decap_8 FILLER_8_244 ();
 sg13g2_decap_8 FILLER_8_251 ();
 sg13g2_decap_8 FILLER_8_258 ();
 sg13g2_decap_8 FILLER_8_265 ();
 sg13g2_decap_8 FILLER_8_272 ();
 sg13g2_decap_8 FILLER_8_279 ();
 sg13g2_decap_4 FILLER_8_286 ();
 sg13g2_fill_2 FILLER_8_290 ();
 sg13g2_decap_8 FILLER_8_296 ();
 sg13g2_decap_8 FILLER_8_303 ();
 sg13g2_decap_8 FILLER_8_310 ();
 sg13g2_decap_8 FILLER_8_317 ();
 sg13g2_decap_8 FILLER_8_324 ();
 sg13g2_decap_8 FILLER_8_331 ();
 sg13g2_decap_8 FILLER_8_338 ();
 sg13g2_decap_8 FILLER_8_345 ();
 sg13g2_decap_8 FILLER_8_352 ();
 sg13g2_decap_8 FILLER_8_359 ();
 sg13g2_decap_8 FILLER_8_366 ();
 sg13g2_decap_4 FILLER_8_373 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_46 ();
 sg13g2_fill_1 FILLER_9_53 ();
 sg13g2_decap_8 FILLER_9_58 ();
 sg13g2_decap_4 FILLER_9_65 ();
 sg13g2_fill_1 FILLER_9_69 ();
 sg13g2_decap_8 FILLER_9_74 ();
 sg13g2_decap_8 FILLER_9_81 ();
 sg13g2_decap_8 FILLER_9_88 ();
 sg13g2_decap_8 FILLER_9_95 ();
 sg13g2_decap_8 FILLER_9_102 ();
 sg13g2_decap_8 FILLER_9_109 ();
 sg13g2_decap_4 FILLER_9_116 ();
 sg13g2_fill_1 FILLER_9_120 ();
 sg13g2_fill_2 FILLER_9_129 ();
 sg13g2_fill_1 FILLER_9_131 ();
 sg13g2_decap_4 FILLER_9_136 ();
 sg13g2_fill_1 FILLER_9_148 ();
 sg13g2_decap_8 FILLER_9_153 ();
 sg13g2_fill_2 FILLER_9_168 ();
 sg13g2_fill_1 FILLER_9_170 ();
 sg13g2_fill_1 FILLER_9_175 ();
 sg13g2_fill_1 FILLER_9_184 ();
 sg13g2_fill_1 FILLER_9_189 ();
 sg13g2_fill_2 FILLER_9_198 ();
 sg13g2_fill_1 FILLER_9_200 ();
 sg13g2_decap_4 FILLER_9_209 ();
 sg13g2_fill_1 FILLER_9_213 ();
 sg13g2_decap_4 FILLER_9_218 ();
 sg13g2_fill_2 FILLER_9_222 ();
 sg13g2_decap_8 FILLER_9_228 ();
 sg13g2_decap_4 FILLER_9_235 ();
 sg13g2_fill_2 FILLER_9_239 ();
 sg13g2_decap_4 FILLER_9_245 ();
 sg13g2_fill_1 FILLER_9_253 ();
 sg13g2_decap_8 FILLER_9_258 ();
 sg13g2_decap_4 FILLER_9_265 ();
 sg13g2_fill_2 FILLER_9_269 ();
 sg13g2_decap_8 FILLER_9_283 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_4 FILLER_9_371 ();
 sg13g2_fill_2 FILLER_9_375 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_4 FILLER_10_364 ();
 sg13g2_fill_1 FILLER_10_368 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_4 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_15 ();
 sg13g2_decap_8 FILLER_11_22 ();
 sg13g2_decap_8 FILLER_11_33 ();
 sg13g2_decap_8 FILLER_11_40 ();
 sg13g2_decap_8 FILLER_11_51 ();
 sg13g2_decap_8 FILLER_11_58 ();
 sg13g2_decap_8 FILLER_11_69 ();
 sg13g2_decap_8 FILLER_11_76 ();
 sg13g2_decap_8 FILLER_11_87 ();
 sg13g2_decap_8 FILLER_11_94 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_123 ();
 sg13g2_decap_8 FILLER_11_130 ();
 sg13g2_decap_8 FILLER_11_141 ();
 sg13g2_decap_8 FILLER_11_148 ();
 sg13g2_decap_8 FILLER_11_159 ();
 sg13g2_decap_8 FILLER_11_166 ();
 sg13g2_decap_8 FILLER_11_177 ();
 sg13g2_decap_8 FILLER_11_184 ();
 sg13g2_decap_8 FILLER_11_195 ();
 sg13g2_decap_8 FILLER_11_202 ();
 sg13g2_decap_8 FILLER_11_213 ();
 sg13g2_decap_8 FILLER_11_220 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_249 ();
 sg13g2_decap_8 FILLER_11_256 ();
 sg13g2_decap_8 FILLER_11_267 ();
 sg13g2_decap_8 FILLER_11_274 ();
 sg13g2_decap_8 FILLER_11_285 ();
 sg13g2_decap_8 FILLER_11_292 ();
 sg13g2_decap_8 FILLER_11_303 ();
 sg13g2_decap_8 FILLER_11_310 ();
 sg13g2_decap_8 FILLER_11_321 ();
 sg13g2_decap_8 FILLER_11_328 ();
 sg13g2_decap_8 FILLER_11_339 ();
 sg13g2_decap_8 FILLER_11_346 ();
 sg13g2_decap_4 FILLER_11_357 ();
 sg13g2_fill_2 FILLER_11_361 ();
 sg13g2_fill_2 FILLER_11_375 ();
endmodule
