magic
tech ihp-sg13g2
magscale 1 2
timestamp 1743691521
<< metal1 >>
rect 1152 10604 20452 10628
rect 1152 10564 4928 10604
rect 4968 10564 5010 10604
rect 5050 10564 5092 10604
rect 5132 10564 5174 10604
rect 5214 10564 5256 10604
rect 5296 10564 20048 10604
rect 20088 10564 20130 10604
rect 20170 10564 20212 10604
rect 20252 10564 20294 10604
rect 20334 10564 20376 10604
rect 20416 10564 20452 10604
rect 1152 10540 20452 10564
rect 1179 10436 1221 10445
rect 1179 10396 1180 10436
rect 1220 10396 1221 10436
rect 1179 10387 1221 10396
rect 2043 10436 2085 10445
rect 2043 10396 2044 10436
rect 2084 10396 2085 10436
rect 2043 10387 2085 10396
rect 3003 10436 3045 10445
rect 3003 10396 3004 10436
rect 3044 10396 3045 10436
rect 3003 10387 3045 10396
rect 3963 10436 4005 10445
rect 3963 10396 3964 10436
rect 4004 10396 4005 10436
rect 3963 10387 4005 10396
rect 4923 10436 4965 10445
rect 4923 10396 4924 10436
rect 4964 10396 4965 10436
rect 4923 10387 4965 10396
rect 5883 10436 5925 10445
rect 5883 10396 5884 10436
rect 5924 10396 5925 10436
rect 5883 10387 5925 10396
rect 6843 10436 6885 10445
rect 6843 10396 6844 10436
rect 6884 10396 6885 10436
rect 6843 10387 6885 10396
rect 7803 10436 7845 10445
rect 7803 10396 7804 10436
rect 7844 10396 7845 10436
rect 7803 10387 7845 10396
rect 8763 10436 8805 10445
rect 8763 10396 8764 10436
rect 8804 10396 8805 10436
rect 8763 10387 8805 10396
rect 9723 10436 9765 10445
rect 9723 10396 9724 10436
rect 9764 10396 9765 10436
rect 9723 10387 9765 10396
rect 10683 10436 10725 10445
rect 10683 10396 10684 10436
rect 10724 10396 10725 10436
rect 10683 10387 10725 10396
rect 11643 10436 11685 10445
rect 11643 10396 11644 10436
rect 11684 10396 11685 10436
rect 11643 10387 11685 10396
rect 12603 10436 12645 10445
rect 12603 10396 12604 10436
rect 12644 10396 12645 10436
rect 12603 10387 12645 10396
rect 13563 10436 13605 10445
rect 13563 10396 13564 10436
rect 13604 10396 13605 10436
rect 13563 10387 13605 10396
rect 14523 10436 14565 10445
rect 14523 10396 14524 10436
rect 14564 10396 14565 10436
rect 14523 10387 14565 10396
rect 15483 10436 15525 10445
rect 15483 10396 15484 10436
rect 15524 10396 15525 10436
rect 15483 10387 15525 10396
rect 16443 10436 16485 10445
rect 16443 10396 16444 10436
rect 16484 10396 16485 10436
rect 16443 10387 16485 10396
rect 17403 10436 17445 10445
rect 17403 10396 17404 10436
rect 17444 10396 17445 10436
rect 17403 10387 17445 10396
rect 18363 10436 18405 10445
rect 18363 10396 18364 10436
rect 18404 10396 18405 10436
rect 18363 10387 18405 10396
rect 19323 10436 19365 10445
rect 19323 10396 19324 10436
rect 19364 10396 19365 10436
rect 19323 10387 19365 10396
rect 18267 10352 18309 10361
rect 18267 10312 18268 10352
rect 18308 10312 18309 10352
rect 18267 10303 18309 10312
rect 1419 10184 1461 10193
rect 1419 10144 1420 10184
rect 1460 10144 1461 10184
rect 1419 10135 1461 10144
rect 2283 10184 2325 10193
rect 2283 10144 2284 10184
rect 2324 10144 2325 10184
rect 2283 10135 2325 10144
rect 3243 10184 3285 10193
rect 3243 10144 3244 10184
rect 3284 10144 3285 10184
rect 3243 10135 3285 10144
rect 4203 10184 4245 10193
rect 4203 10144 4204 10184
rect 4244 10144 4245 10184
rect 4203 10135 4245 10144
rect 5163 10184 5205 10193
rect 5163 10144 5164 10184
rect 5204 10144 5205 10184
rect 5163 10135 5205 10144
rect 6123 10184 6165 10193
rect 6123 10144 6124 10184
rect 6164 10144 6165 10184
rect 6123 10135 6165 10144
rect 7083 10184 7125 10193
rect 7083 10144 7084 10184
rect 7124 10144 7125 10184
rect 7083 10135 7125 10144
rect 8043 10184 8085 10193
rect 8043 10144 8044 10184
rect 8084 10144 8085 10184
rect 8043 10135 8085 10144
rect 9003 10184 9045 10193
rect 9003 10144 9004 10184
rect 9044 10144 9045 10184
rect 9003 10135 9045 10144
rect 9963 10184 10005 10193
rect 9963 10144 9964 10184
rect 10004 10144 10005 10184
rect 9963 10135 10005 10144
rect 10923 10184 10965 10193
rect 10923 10144 10924 10184
rect 10964 10144 10965 10184
rect 10923 10135 10965 10144
rect 11883 10184 11925 10193
rect 11883 10144 11884 10184
rect 11924 10144 11925 10184
rect 11883 10135 11925 10144
rect 12843 10184 12885 10193
rect 12843 10144 12844 10184
rect 12884 10144 12885 10184
rect 12843 10135 12885 10144
rect 13803 10184 13845 10193
rect 13803 10144 13804 10184
rect 13844 10144 13845 10184
rect 13803 10135 13845 10144
rect 14763 10184 14805 10193
rect 14763 10144 14764 10184
rect 14804 10144 14805 10184
rect 14763 10135 14805 10144
rect 15723 10184 15765 10193
rect 15723 10144 15724 10184
rect 15764 10144 15765 10184
rect 15723 10135 15765 10144
rect 16683 10184 16725 10193
rect 16683 10144 16684 10184
rect 16724 10144 16725 10184
rect 16683 10135 16725 10144
rect 17643 10184 17685 10193
rect 17643 10144 17644 10184
rect 17684 10144 17685 10184
rect 17643 10135 17685 10144
rect 18027 10184 18069 10193
rect 18027 10144 18028 10184
rect 18068 10144 18069 10184
rect 18027 10135 18069 10144
rect 18603 10184 18645 10193
rect 18603 10144 18604 10184
rect 18644 10144 18645 10184
rect 18603 10135 18645 10144
rect 18987 10184 19029 10193
rect 18987 10144 18988 10184
rect 19028 10144 19029 10184
rect 18987 10135 19029 10144
rect 19563 10184 19605 10193
rect 19563 10144 19564 10184
rect 19604 10144 19605 10184
rect 19563 10135 19605 10144
rect 19755 10184 19797 10193
rect 19755 10144 19756 10184
rect 19796 10144 19797 10184
rect 19755 10135 19797 10144
rect 20139 10184 20181 10193
rect 20139 10144 20140 10184
rect 20180 10144 20181 10184
rect 20139 10135 20181 10144
rect 19227 10016 19269 10025
rect 19227 9976 19228 10016
rect 19268 9976 19269 10016
rect 19227 9967 19269 9976
rect 19995 10016 20037 10025
rect 19995 9976 19996 10016
rect 20036 9976 20037 10016
rect 19995 9967 20037 9976
rect 20379 10016 20421 10025
rect 20379 9976 20380 10016
rect 20420 9976 20421 10016
rect 20379 9967 20421 9976
rect 1152 9848 20448 9872
rect 1152 9808 3688 9848
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 4056 9808 18808 9848
rect 18848 9808 18890 9848
rect 18930 9808 18972 9848
rect 19012 9808 19054 9848
rect 19094 9808 19136 9848
rect 19176 9808 20448 9848
rect 1152 9784 20448 9808
rect 2331 9680 2373 9689
rect 2331 9640 2332 9680
rect 2372 9640 2373 9680
rect 2331 9631 2373 9640
rect 10875 9680 10917 9689
rect 10875 9640 10876 9680
rect 10916 9640 10917 9680
rect 10875 9631 10917 9640
rect 13755 9680 13797 9689
rect 13755 9640 13756 9680
rect 13796 9640 13797 9680
rect 13755 9631 13797 9640
rect 14811 9680 14853 9689
rect 14811 9640 14812 9680
rect 14852 9640 14853 9680
rect 14811 9631 14853 9640
rect 16635 9680 16677 9689
rect 16635 9640 16636 9680
rect 16676 9640 16677 9680
rect 16635 9631 16677 9640
rect 18747 9680 18789 9689
rect 18747 9640 18748 9680
rect 18788 9640 18789 9680
rect 18747 9631 18789 9640
rect 19131 9680 19173 9689
rect 19131 9640 19132 9680
rect 19172 9640 19173 9680
rect 19131 9631 19173 9640
rect 14139 9596 14181 9605
rect 14139 9556 14140 9596
rect 14180 9556 14181 9596
rect 14139 9547 14181 9556
rect 2571 9512 2613 9521
rect 2571 9472 2572 9512
rect 2612 9472 2613 9512
rect 2571 9463 2613 9472
rect 11115 9512 11157 9521
rect 11115 9472 11116 9512
rect 11156 9472 11157 9512
rect 11115 9463 11157 9472
rect 11307 9512 11349 9521
rect 11307 9472 11308 9512
rect 11348 9472 11349 9512
rect 11307 9463 11349 9472
rect 11547 9512 11589 9521
rect 11547 9472 11548 9512
rect 11588 9472 11589 9512
rect 11547 9463 11589 9472
rect 13995 9512 14037 9521
rect 13995 9472 13996 9512
rect 14036 9472 14037 9512
rect 13995 9463 14037 9472
rect 14379 9512 14421 9521
rect 14379 9472 14380 9512
rect 14420 9472 14421 9512
rect 14379 9463 14421 9472
rect 15051 9512 15093 9521
rect 15051 9472 15052 9512
rect 15092 9472 15093 9512
rect 15051 9463 15093 9472
rect 16395 9512 16437 9521
rect 16395 9472 16396 9512
rect 16436 9472 16437 9512
rect 16395 9463 16437 9472
rect 17547 9512 17589 9521
rect 17547 9472 17548 9512
rect 17588 9472 17589 9512
rect 17547 9463 17589 9472
rect 18123 9512 18165 9521
rect 18123 9472 18124 9512
rect 18164 9472 18165 9512
rect 18123 9463 18165 9472
rect 18507 9512 18549 9521
rect 18507 9472 18508 9512
rect 18548 9472 18549 9512
rect 18507 9463 18549 9472
rect 18891 9512 18933 9521
rect 18891 9472 18892 9512
rect 18932 9472 18933 9512
rect 18891 9463 18933 9472
rect 19467 9512 19509 9521
rect 19467 9472 19468 9512
rect 19508 9472 19509 9512
rect 19467 9463 19509 9472
rect 19851 9512 19893 9521
rect 19851 9472 19852 9512
rect 19892 9472 19893 9512
rect 19851 9463 19893 9472
rect 20139 9512 20181 9521
rect 20139 9472 20140 9512
rect 20180 9472 20181 9512
rect 20139 9463 20181 9472
rect 17787 9260 17829 9269
rect 17787 9220 17788 9260
rect 17828 9220 17829 9260
rect 17787 9211 17829 9220
rect 18363 9260 18405 9269
rect 18363 9220 18364 9260
rect 18404 9220 18405 9260
rect 18363 9211 18405 9220
rect 19227 9260 19269 9269
rect 19227 9220 19228 9260
rect 19268 9220 19269 9260
rect 19227 9211 19269 9220
rect 19611 9260 19653 9269
rect 19611 9220 19612 9260
rect 19652 9220 19653 9260
rect 19611 9211 19653 9220
rect 20379 9260 20421 9269
rect 20379 9220 20380 9260
rect 20420 9220 20421 9260
rect 20379 9211 20421 9220
rect 1152 9092 20452 9116
rect 1152 9052 4928 9092
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 5296 9052 20048 9092
rect 20088 9052 20130 9092
rect 20170 9052 20212 9092
rect 20252 9052 20294 9092
rect 20334 9052 20376 9092
rect 20416 9052 20452 9092
rect 1152 9028 20452 9052
rect 9051 8924 9093 8933
rect 9051 8884 9052 8924
rect 9092 8884 9093 8924
rect 9051 8875 9093 8884
rect 12987 8924 13029 8933
rect 12987 8884 12988 8924
rect 13028 8884 13029 8924
rect 12987 8875 13029 8884
rect 13659 8924 13701 8933
rect 13659 8884 13660 8924
rect 13700 8884 13701 8924
rect 13659 8875 13701 8884
rect 15387 8924 15429 8933
rect 15387 8884 15388 8924
rect 15428 8884 15429 8924
rect 15387 8875 15429 8884
rect 19227 8924 19269 8933
rect 19227 8884 19228 8924
rect 19268 8884 19269 8924
rect 19227 8875 19269 8884
rect 19611 8924 19653 8933
rect 19611 8884 19612 8924
rect 19652 8884 19653 8924
rect 19611 8875 19653 8884
rect 17499 8840 17541 8849
rect 17499 8800 17500 8840
rect 17540 8800 17541 8840
rect 17499 8791 17541 8800
rect 1899 8672 1941 8681
rect 1899 8632 1900 8672
rect 1940 8632 1941 8672
rect 1899 8623 1941 8632
rect 2139 8672 2181 8681
rect 2139 8632 2140 8672
rect 2180 8632 2181 8672
rect 2139 8623 2181 8632
rect 8811 8672 8853 8681
rect 8811 8632 8812 8672
rect 8852 8632 8853 8672
rect 8811 8623 8853 8632
rect 13227 8672 13269 8681
rect 13227 8632 13228 8672
rect 13268 8632 13269 8672
rect 13227 8623 13269 8632
rect 13419 8672 13461 8681
rect 13419 8632 13420 8672
rect 13460 8632 13461 8672
rect 13419 8623 13461 8632
rect 13803 8672 13845 8681
rect 13803 8632 13804 8672
rect 13844 8632 13845 8672
rect 13803 8623 13845 8632
rect 14043 8672 14085 8681
rect 14043 8632 14044 8672
rect 14084 8632 14085 8672
rect 14043 8623 14085 8632
rect 15627 8672 15669 8681
rect 15627 8632 15628 8672
rect 15668 8632 15669 8672
rect 15627 8623 15669 8632
rect 17259 8672 17301 8681
rect 17259 8632 17260 8672
rect 17300 8632 17301 8672
rect 17259 8623 17301 8632
rect 18987 8672 19029 8681
rect 18987 8632 18988 8672
rect 19028 8632 19029 8672
rect 18987 8623 19029 8632
rect 19371 8672 19413 8681
rect 19371 8632 19372 8672
rect 19412 8632 19413 8672
rect 19371 8623 19413 8632
rect 19755 8672 19797 8681
rect 19755 8632 19756 8672
rect 19796 8632 19797 8672
rect 19755 8623 19797 8632
rect 19995 8672 20037 8681
rect 19995 8632 19996 8672
rect 20036 8632 20037 8672
rect 19995 8623 20037 8632
rect 20139 8672 20181 8681
rect 20139 8632 20140 8672
rect 20180 8632 20181 8672
rect 20139 8623 20181 8632
rect 20379 8504 20421 8513
rect 20379 8464 20380 8504
rect 20420 8464 20421 8504
rect 20379 8455 20421 8464
rect 1152 8336 20448 8360
rect 1152 8296 3688 8336
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 4056 8296 18808 8336
rect 18848 8296 18890 8336
rect 18930 8296 18972 8336
rect 19012 8296 19054 8336
rect 19094 8296 19136 8336
rect 19176 8296 20448 8336
rect 1152 8272 20448 8296
rect 1947 8168 1989 8177
rect 1947 8128 1948 8168
rect 1988 8128 1989 8168
rect 1947 8119 1989 8128
rect 6747 8168 6789 8177
rect 6747 8128 6748 8168
rect 6788 8128 6789 8168
rect 6747 8119 6789 8128
rect 8379 8168 8421 8177
rect 8379 8128 8380 8168
rect 8420 8128 8421 8168
rect 8379 8119 8421 8128
rect 15579 8168 15621 8177
rect 15579 8128 15580 8168
rect 15620 8128 15621 8168
rect 15579 8119 15621 8128
rect 15963 8168 16005 8177
rect 15963 8128 15964 8168
rect 16004 8128 16005 8168
rect 15963 8119 16005 8128
rect 7899 8084 7941 8093
rect 7899 8044 7900 8084
rect 7940 8044 7941 8084
rect 7899 8035 7941 8044
rect 2187 8000 2229 8009
rect 2187 7960 2188 8000
rect 2228 7960 2229 8000
rect 2187 7951 2229 7960
rect 4491 8000 4533 8009
rect 4491 7960 4492 8000
rect 4532 7960 4533 8000
rect 4491 7951 4533 7960
rect 6987 8000 7029 8009
rect 6987 7960 6988 8000
rect 7028 7960 7029 8000
rect 6987 7951 7029 7960
rect 7659 8000 7701 8009
rect 7659 7960 7660 8000
rect 7700 7960 7701 8000
rect 7659 7951 7701 7960
rect 8619 8000 8661 8009
rect 8619 7960 8620 8000
rect 8660 7960 8661 8000
rect 8619 7951 8661 7960
rect 9003 8000 9045 8009
rect 9003 7960 9004 8000
rect 9044 7960 9045 8000
rect 9003 7951 9045 7960
rect 9963 8000 10005 8009
rect 9963 7960 9964 8000
rect 10004 7960 10005 8000
rect 9963 7951 10005 7960
rect 15339 8000 15381 8009
rect 15339 7960 15340 8000
rect 15380 7960 15381 8000
rect 15339 7951 15381 7960
rect 15723 8000 15765 8009
rect 15723 7960 15724 8000
rect 15764 7960 15765 8000
rect 15723 7951 15765 7960
rect 17067 8000 17109 8009
rect 17067 7960 17068 8000
rect 17108 7960 17109 8000
rect 17067 7951 17109 7960
rect 17931 8000 17973 8009
rect 17931 7960 17932 8000
rect 17972 7960 17973 8000
rect 17931 7951 17973 7960
rect 19755 8000 19797 8009
rect 19755 7960 19756 8000
rect 19796 7960 19797 8000
rect 19755 7951 19797 7960
rect 20139 8000 20181 8009
rect 20139 7960 20140 8000
rect 20180 7960 20181 8000
rect 20139 7951 20181 7960
rect 9243 7832 9285 7841
rect 9243 7792 9244 7832
rect 9284 7792 9285 7832
rect 9243 7783 9285 7792
rect 17307 7832 17349 7841
rect 17307 7792 17308 7832
rect 17348 7792 17349 7832
rect 17307 7783 17349 7792
rect 19995 7832 20037 7841
rect 19995 7792 19996 7832
rect 20036 7792 20037 7832
rect 19995 7783 20037 7792
rect 4731 7748 4773 7757
rect 4731 7708 4732 7748
rect 4772 7708 4773 7748
rect 4731 7699 4773 7708
rect 10203 7748 10245 7757
rect 10203 7708 10204 7748
rect 10244 7708 10245 7748
rect 10203 7699 10245 7708
rect 18171 7748 18213 7757
rect 18171 7708 18172 7748
rect 18212 7708 18213 7748
rect 18171 7699 18213 7708
rect 20379 7748 20421 7757
rect 20379 7708 20380 7748
rect 20420 7708 20421 7748
rect 20379 7699 20421 7708
rect 1152 7580 20452 7604
rect 1152 7540 4928 7580
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 5296 7540 20048 7580
rect 20088 7540 20130 7580
rect 20170 7540 20212 7580
rect 20252 7540 20294 7580
rect 20334 7540 20376 7580
rect 20416 7540 20452 7580
rect 1152 7516 20452 7540
rect 2091 7160 2133 7169
rect 2091 7120 2092 7160
rect 2132 7120 2133 7160
rect 2091 7111 2133 7120
rect 4875 7160 4917 7169
rect 4875 7120 4876 7160
rect 4916 7120 4917 7160
rect 4875 7111 4917 7120
rect 5115 7160 5157 7169
rect 5115 7120 5116 7160
rect 5156 7120 5157 7160
rect 5115 7111 5157 7120
rect 7371 7160 7413 7169
rect 7371 7120 7372 7160
rect 7412 7120 7413 7160
rect 7371 7111 7413 7120
rect 7755 7160 7797 7169
rect 7755 7120 7756 7160
rect 7796 7120 7797 7160
rect 7755 7111 7797 7120
rect 7995 7160 8037 7169
rect 7995 7120 7996 7160
rect 8036 7120 8037 7160
rect 7995 7111 8037 7120
rect 15243 7160 15285 7169
rect 15243 7120 15244 7160
rect 15284 7120 15285 7160
rect 15243 7111 15285 7120
rect 15483 7160 15525 7169
rect 15483 7120 15484 7160
rect 15524 7120 15525 7160
rect 15483 7111 15525 7120
rect 19083 7160 19125 7169
rect 19083 7120 19084 7160
rect 19124 7120 19125 7160
rect 19083 7111 19125 7120
rect 19467 7160 19509 7169
rect 19467 7120 19468 7160
rect 19508 7120 19509 7160
rect 19467 7111 19509 7120
rect 19851 7160 19893 7169
rect 19851 7120 19852 7160
rect 19892 7120 19893 7160
rect 19851 7111 19893 7120
rect 20091 7160 20133 7169
rect 20091 7120 20092 7160
rect 20132 7120 20133 7160
rect 20091 7111 20133 7120
rect 19323 7076 19365 7085
rect 19323 7036 19324 7076
rect 19364 7036 19365 7076
rect 19323 7027 19365 7036
rect 2331 6992 2373 7001
rect 2331 6952 2332 6992
rect 2372 6952 2373 6992
rect 2331 6943 2373 6952
rect 7611 6992 7653 7001
rect 7611 6952 7612 6992
rect 7652 6952 7653 6992
rect 7611 6943 7653 6952
rect 19707 6992 19749 7001
rect 19707 6952 19708 6992
rect 19748 6952 19749 6992
rect 19707 6943 19749 6952
rect 1152 6824 20448 6848
rect 1152 6784 3688 6824
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 4056 6784 18808 6824
rect 18848 6784 18890 6824
rect 18930 6784 18972 6824
rect 19012 6784 19054 6824
rect 19094 6784 19136 6824
rect 19176 6784 20448 6824
rect 1152 6760 20448 6784
rect 2331 6656 2373 6665
rect 2331 6616 2332 6656
rect 2372 6616 2373 6656
rect 2331 6607 2373 6616
rect 20379 6656 20421 6665
rect 20379 6616 20380 6656
rect 20420 6616 20421 6656
rect 20379 6607 20421 6616
rect 2091 6488 2133 6497
rect 2091 6448 2092 6488
rect 2132 6448 2133 6488
rect 2091 6439 2133 6448
rect 3531 6488 3573 6497
rect 3531 6448 3532 6488
rect 3572 6448 3573 6488
rect 3531 6439 3573 6448
rect 5211 6488 5253 6497
rect 5211 6448 5212 6488
rect 5252 6448 5253 6488
rect 5211 6439 5253 6448
rect 5451 6488 5493 6497
rect 5451 6448 5452 6488
rect 5492 6448 5493 6488
rect 5451 6439 5493 6448
rect 6219 6488 6261 6497
rect 6219 6448 6220 6488
rect 6260 6448 6261 6488
rect 6219 6439 6261 6448
rect 8907 6488 8949 6497
rect 8907 6448 8908 6488
rect 8948 6448 8949 6488
rect 8907 6439 8949 6448
rect 9147 6488 9189 6497
rect 9147 6448 9148 6488
rect 9188 6448 9189 6488
rect 9147 6439 9189 6448
rect 9387 6488 9429 6497
rect 9387 6448 9388 6488
rect 9428 6448 9429 6488
rect 9387 6439 9429 6448
rect 12843 6488 12885 6497
rect 12843 6448 12844 6488
rect 12884 6448 12885 6488
rect 12843 6439 12885 6448
rect 14475 6488 14517 6497
rect 14475 6448 14476 6488
rect 14516 6448 14517 6488
rect 14475 6439 14517 6448
rect 16683 6488 16725 6497
rect 16683 6448 16684 6488
rect 16724 6448 16725 6488
rect 16683 6439 16725 6448
rect 17067 6488 17109 6497
rect 17067 6448 17068 6488
rect 17108 6448 17109 6488
rect 17067 6439 17109 6448
rect 19275 6488 19317 6497
rect 19275 6448 19276 6488
rect 19316 6448 19317 6488
rect 19275 6439 19317 6448
rect 19755 6488 19797 6497
rect 19755 6448 19756 6488
rect 19796 6448 19797 6488
rect 19755 6439 19797 6448
rect 20139 6488 20181 6497
rect 20139 6448 20140 6488
rect 20180 6448 20181 6488
rect 20139 6439 20181 6448
rect 6459 6320 6501 6329
rect 6459 6280 6460 6320
rect 6500 6280 6501 6320
rect 6459 6271 6501 6280
rect 19995 6320 20037 6329
rect 19995 6280 19996 6320
rect 20036 6280 20037 6320
rect 19995 6271 20037 6280
rect 3771 6236 3813 6245
rect 3771 6196 3772 6236
rect 3812 6196 3813 6236
rect 3771 6187 3813 6196
rect 9627 6236 9669 6245
rect 9627 6196 9628 6236
rect 9668 6196 9669 6236
rect 9627 6187 9669 6196
rect 13083 6236 13125 6245
rect 13083 6196 13084 6236
rect 13124 6196 13125 6236
rect 13083 6187 13125 6196
rect 14715 6236 14757 6245
rect 14715 6196 14716 6236
rect 14756 6196 14757 6236
rect 14715 6187 14757 6196
rect 16923 6236 16965 6245
rect 16923 6196 16924 6236
rect 16964 6196 16965 6236
rect 16923 6187 16965 6196
rect 17307 6236 17349 6245
rect 17307 6196 17308 6236
rect 17348 6196 17349 6236
rect 17307 6187 17349 6196
rect 19515 6236 19557 6245
rect 19515 6196 19516 6236
rect 19556 6196 19557 6236
rect 19515 6187 19557 6196
rect 1152 6068 20452 6092
rect 1152 6028 4928 6068
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 5296 6028 20048 6068
rect 20088 6028 20130 6068
rect 20170 6028 20212 6068
rect 20252 6028 20294 6068
rect 20334 6028 20376 6068
rect 20416 6028 20452 6068
rect 1152 6004 20452 6028
rect 20379 5900 20421 5909
rect 20379 5860 20380 5900
rect 20420 5860 20421 5900
rect 20379 5851 20421 5860
rect 19995 5816 20037 5825
rect 19995 5776 19996 5816
rect 20036 5776 20037 5816
rect 19995 5767 20037 5776
rect 1995 5648 2037 5657
rect 1995 5608 1996 5648
rect 2036 5608 2037 5648
rect 1995 5599 2037 5608
rect 2475 5648 2517 5657
rect 2475 5608 2476 5648
rect 2516 5608 2517 5648
rect 2475 5599 2517 5608
rect 2715 5648 2757 5657
rect 2715 5608 2716 5648
rect 2756 5608 2757 5648
rect 2715 5599 2757 5608
rect 4683 5648 4725 5657
rect 4683 5608 4684 5648
rect 4724 5608 4725 5648
rect 4683 5599 4725 5608
rect 9003 5648 9045 5657
rect 9003 5608 9004 5648
rect 9044 5608 9045 5648
rect 9003 5599 9045 5608
rect 15723 5648 15765 5657
rect 15723 5608 15724 5648
rect 15764 5608 15765 5648
rect 15723 5599 15765 5608
rect 16971 5648 17013 5657
rect 16971 5608 16972 5648
rect 17012 5608 17013 5648
rect 16971 5599 17013 5608
rect 18507 5648 18549 5657
rect 18507 5608 18508 5648
rect 18548 5608 18549 5648
rect 18507 5599 18549 5608
rect 18891 5648 18933 5657
rect 18891 5608 18892 5648
rect 18932 5608 18933 5648
rect 18891 5599 18933 5608
rect 19371 5648 19413 5657
rect 19371 5608 19372 5648
rect 19412 5608 19413 5648
rect 19371 5599 19413 5608
rect 19755 5648 19797 5657
rect 19755 5608 19756 5648
rect 19796 5608 19797 5648
rect 19755 5599 19797 5608
rect 20139 5648 20181 5657
rect 20139 5608 20140 5648
rect 20180 5608 20181 5648
rect 20139 5599 20181 5608
rect 4923 5564 4965 5573
rect 4923 5524 4924 5564
rect 4964 5524 4965 5564
rect 4923 5515 4965 5524
rect 2235 5480 2277 5489
rect 2235 5440 2236 5480
rect 2276 5440 2277 5480
rect 2235 5431 2277 5440
rect 9243 5480 9285 5489
rect 9243 5440 9244 5480
rect 9284 5440 9285 5480
rect 9243 5431 9285 5440
rect 15963 5480 16005 5489
rect 15963 5440 15964 5480
rect 16004 5440 16005 5480
rect 15963 5431 16005 5440
rect 17211 5480 17253 5489
rect 17211 5440 17212 5480
rect 17252 5440 17253 5480
rect 17211 5431 17253 5440
rect 18747 5480 18789 5489
rect 18747 5440 18748 5480
rect 18788 5440 18789 5480
rect 18747 5431 18789 5440
rect 19131 5480 19173 5489
rect 19131 5440 19132 5480
rect 19172 5440 19173 5480
rect 19131 5431 19173 5440
rect 19611 5480 19653 5489
rect 19611 5440 19612 5480
rect 19652 5440 19653 5480
rect 19611 5431 19653 5440
rect 1152 5312 20448 5336
rect 1152 5272 3688 5312
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 4056 5272 18808 5312
rect 18848 5272 18890 5312
rect 18930 5272 18972 5312
rect 19012 5272 19054 5312
rect 19094 5272 19136 5312
rect 19176 5272 20448 5312
rect 1152 5248 20448 5272
rect 19323 5060 19365 5069
rect 19323 5020 19324 5060
rect 19364 5020 19365 5060
rect 19323 5011 19365 5020
rect 4971 4976 5013 4985
rect 4971 4936 4972 4976
rect 5012 4936 5013 4976
rect 4971 4927 5013 4936
rect 8715 4976 8757 4985
rect 8715 4936 8716 4976
rect 8756 4936 8757 4976
rect 8715 4927 8757 4936
rect 9099 4976 9141 4985
rect 9099 4936 9100 4976
rect 9140 4936 9141 4976
rect 9099 4927 9141 4936
rect 17067 4976 17109 4985
rect 17067 4936 17068 4976
rect 17108 4936 17109 4976
rect 17067 4927 17109 4936
rect 18730 4976 18788 4977
rect 18730 4936 18739 4976
rect 18779 4936 18788 4976
rect 18730 4935 18788 4936
rect 19083 4976 19125 4985
rect 19083 4936 19084 4976
rect 19124 4936 19125 4976
rect 19083 4927 19125 4936
rect 19467 4976 19509 4985
rect 19467 4936 19468 4976
rect 19508 4936 19509 4976
rect 19467 4927 19509 4936
rect 20139 4976 20181 4985
rect 20139 4936 20140 4976
rect 20180 4936 20181 4976
rect 20139 4927 20181 4936
rect 20379 4976 20421 4985
rect 20379 4936 20380 4976
rect 20420 4936 20421 4976
rect 20379 4927 20421 4936
rect 8955 4808 8997 4817
rect 8955 4768 8956 4808
rect 8996 4768 8997 4808
rect 8955 4759 8997 4768
rect 18939 4808 18981 4817
rect 18939 4768 18940 4808
rect 18980 4768 18981 4808
rect 18939 4759 18981 4768
rect 5211 4724 5253 4733
rect 5211 4684 5212 4724
rect 5252 4684 5253 4724
rect 5211 4675 5253 4684
rect 9339 4724 9381 4733
rect 9339 4684 9340 4724
rect 9380 4684 9381 4724
rect 9339 4675 9381 4684
rect 17307 4724 17349 4733
rect 17307 4684 17308 4724
rect 17348 4684 17349 4724
rect 17307 4675 17349 4684
rect 19707 4724 19749 4733
rect 19707 4684 19708 4724
rect 19748 4684 19749 4724
rect 19707 4675 19749 4684
rect 1152 4556 20452 4580
rect 1152 4516 4928 4556
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 5296 4516 20048 4556
rect 20088 4516 20130 4556
rect 20170 4516 20212 4556
rect 20252 4516 20294 4556
rect 20334 4516 20376 4556
rect 20416 4516 20452 4556
rect 1152 4492 20452 4516
rect 10875 4388 10917 4397
rect 10875 4348 10876 4388
rect 10916 4348 10917 4388
rect 10875 4339 10917 4348
rect 3867 4304 3909 4313
rect 3867 4264 3868 4304
rect 3908 4264 3909 4304
rect 3867 4255 3909 4264
rect 6459 4304 6501 4313
rect 6459 4264 6460 4304
rect 6500 4264 6501 4304
rect 6459 4255 6501 4264
rect 20379 4304 20421 4313
rect 20379 4264 20380 4304
rect 20420 4264 20421 4304
rect 20379 4255 20421 4264
rect 2283 4136 2325 4145
rect 2283 4096 2284 4136
rect 2324 4096 2325 4136
rect 2283 4087 2325 4096
rect 3627 4136 3669 4145
rect 3627 4096 3628 4136
rect 3668 4096 3669 4136
rect 3627 4087 3669 4096
rect 6219 4136 6261 4145
rect 6219 4096 6220 4136
rect 6260 4096 6261 4136
rect 6219 4087 6261 4096
rect 10251 4136 10293 4145
rect 10251 4096 10252 4136
rect 10292 4096 10293 4136
rect 10251 4087 10293 4096
rect 10587 4136 10629 4145
rect 10587 4096 10588 4136
rect 10628 4096 10629 4136
rect 10587 4087 10629 4096
rect 11595 4136 11637 4145
rect 11595 4096 11596 4136
rect 11636 4096 11637 4136
rect 11595 4087 11637 4096
rect 11979 4136 12021 4145
rect 11979 4096 11980 4136
rect 12020 4096 12021 4136
rect 11979 4087 12021 4096
rect 13611 4136 13653 4145
rect 13611 4096 13612 4136
rect 13652 4096 13653 4136
rect 13611 4087 13653 4096
rect 14283 4136 14325 4145
rect 14283 4096 14284 4136
rect 14324 4096 14325 4136
rect 14283 4087 14325 4096
rect 14667 4136 14709 4145
rect 14667 4096 14668 4136
rect 14708 4096 14709 4136
rect 14667 4087 14709 4096
rect 16395 4136 16437 4145
rect 16395 4096 16396 4136
rect 16436 4096 16437 4136
rect 16395 4087 16437 4096
rect 17931 4136 17973 4145
rect 17931 4096 17932 4136
rect 17972 4096 17973 4136
rect 17931 4087 17973 4096
rect 19083 4136 19125 4145
rect 19083 4096 19084 4136
rect 19124 4096 19125 4136
rect 19083 4087 19125 4096
rect 19659 4136 19701 4145
rect 19659 4096 19660 4136
rect 19700 4096 19701 4136
rect 19659 4087 19701 4096
rect 20139 4136 20181 4145
rect 20139 4096 20140 4136
rect 20180 4096 20181 4136
rect 20139 4087 20181 4096
rect 11835 4052 11877 4061
rect 11835 4012 11836 4052
rect 11876 4012 11877 4052
rect 11835 4003 11877 4012
rect 19323 4052 19365 4061
rect 19323 4012 19324 4052
rect 19364 4012 19365 4052
rect 19323 4003 19365 4012
rect 2523 3968 2565 3977
rect 2523 3928 2524 3968
rect 2564 3928 2565 3968
rect 2523 3919 2565 3928
rect 10491 3968 10533 3977
rect 10491 3928 10492 3968
rect 10532 3928 10533 3968
rect 10491 3919 10533 3928
rect 12219 3968 12261 3977
rect 12219 3928 12220 3968
rect 12260 3928 12261 3968
rect 12219 3919 12261 3928
rect 13371 3968 13413 3977
rect 13371 3928 13372 3968
rect 13412 3928 13413 3968
rect 13371 3919 13413 3928
rect 14043 3968 14085 3977
rect 14043 3928 14044 3968
rect 14084 3928 14085 3968
rect 14043 3919 14085 3928
rect 14427 3968 14469 3977
rect 14427 3928 14428 3968
rect 14468 3928 14469 3968
rect 14427 3919 14469 3928
rect 16155 3968 16197 3977
rect 16155 3928 16156 3968
rect 16196 3928 16197 3968
rect 16155 3919 16197 3928
rect 17691 3968 17733 3977
rect 17691 3928 17692 3968
rect 17732 3928 17733 3968
rect 17691 3919 17733 3928
rect 19419 3968 19461 3977
rect 19419 3928 19420 3968
rect 19460 3928 19461 3968
rect 19419 3919 19461 3928
rect 1152 3800 20448 3824
rect 1152 3760 3688 3800
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 4056 3760 18808 3800
rect 18848 3760 18890 3800
rect 18930 3760 18972 3800
rect 19012 3760 19054 3800
rect 19094 3760 19136 3800
rect 19176 3760 20448 3800
rect 1152 3736 20448 3760
rect 20379 3632 20421 3641
rect 20379 3592 20380 3632
rect 20420 3592 20421 3632
rect 20379 3583 20421 3592
rect 6267 3548 6309 3557
rect 6267 3508 6268 3548
rect 6308 3508 6309 3548
rect 6267 3499 6309 3508
rect 19995 3548 20037 3557
rect 19995 3508 19996 3548
rect 20036 3508 20037 3548
rect 19995 3499 20037 3508
rect 2475 3464 2517 3473
rect 2475 3424 2476 3464
rect 2516 3424 2517 3464
rect 2475 3415 2517 3424
rect 6027 3464 6069 3473
rect 6027 3424 6028 3464
rect 6068 3424 6069 3464
rect 6027 3415 6069 3424
rect 15723 3464 15765 3473
rect 15723 3424 15724 3464
rect 15764 3424 15765 3464
rect 15723 3415 15765 3424
rect 17067 3464 17109 3473
rect 17067 3424 17068 3464
rect 17108 3424 17109 3464
rect 17067 3415 17109 3424
rect 18987 3464 19029 3473
rect 18987 3424 18988 3464
rect 19028 3424 19029 3464
rect 18987 3415 19029 3424
rect 19563 3464 19605 3473
rect 19563 3424 19564 3464
rect 19604 3424 19605 3464
rect 19563 3415 19605 3424
rect 19755 3464 19797 3473
rect 19755 3424 19756 3464
rect 19796 3424 19797 3464
rect 19755 3415 19797 3424
rect 20139 3464 20181 3473
rect 20139 3424 20140 3464
rect 20180 3424 20181 3464
rect 20139 3415 20181 3424
rect 19227 3296 19269 3305
rect 19227 3256 19228 3296
rect 19268 3256 19269 3296
rect 19227 3247 19269 3256
rect 2715 3212 2757 3221
rect 2715 3172 2716 3212
rect 2756 3172 2757 3212
rect 2715 3163 2757 3172
rect 15483 3212 15525 3221
rect 15483 3172 15484 3212
rect 15524 3172 15525 3212
rect 15483 3163 15525 3172
rect 16827 3212 16869 3221
rect 16827 3172 16828 3212
rect 16868 3172 16869 3212
rect 16827 3163 16869 3172
rect 19323 3212 19365 3221
rect 19323 3172 19324 3212
rect 19364 3172 19365 3212
rect 19323 3163 19365 3172
rect 1152 3044 20452 3068
rect 1152 3004 4928 3044
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 5296 3004 20048 3044
rect 20088 3004 20130 3044
rect 20170 3004 20212 3044
rect 20252 3004 20294 3044
rect 20334 3004 20376 3044
rect 20416 3004 20452 3044
rect 1152 2980 20452 3004
rect 17211 2876 17253 2885
rect 17211 2836 17212 2876
rect 17252 2836 17253 2876
rect 17211 2827 17253 2836
rect 20379 2876 20421 2885
rect 20379 2836 20380 2876
rect 20420 2836 20421 2876
rect 20379 2827 20421 2836
rect 2331 2792 2373 2801
rect 2331 2752 2332 2792
rect 2372 2752 2373 2792
rect 2331 2743 2373 2752
rect 2091 2624 2133 2633
rect 2091 2584 2092 2624
rect 2132 2584 2133 2624
rect 2091 2575 2133 2584
rect 2475 2624 2517 2633
rect 2475 2584 2476 2624
rect 2516 2584 2517 2624
rect 2475 2575 2517 2584
rect 9195 2624 9237 2633
rect 9195 2584 9196 2624
rect 9236 2584 9237 2624
rect 9195 2575 9237 2584
rect 9579 2624 9621 2633
rect 9579 2584 9580 2624
rect 9620 2584 9621 2624
rect 9579 2575 9621 2584
rect 9963 2624 10005 2633
rect 9963 2584 9964 2624
rect 10004 2584 10005 2624
rect 9963 2575 10005 2584
rect 10347 2624 10389 2633
rect 10347 2584 10348 2624
rect 10388 2584 10389 2624
rect 10347 2575 10389 2584
rect 10731 2624 10773 2633
rect 10731 2584 10732 2624
rect 10772 2584 10773 2624
rect 10731 2575 10773 2584
rect 11115 2624 11157 2633
rect 11115 2584 11116 2624
rect 11156 2584 11157 2624
rect 11115 2575 11157 2584
rect 12843 2624 12885 2633
rect 12843 2584 12844 2624
rect 12884 2584 12885 2624
rect 12843 2575 12885 2584
rect 13227 2624 13269 2633
rect 13227 2584 13228 2624
rect 13268 2584 13269 2624
rect 13227 2575 13269 2584
rect 13611 2624 13653 2633
rect 13611 2584 13612 2624
rect 13652 2584 13653 2624
rect 13611 2575 13653 2584
rect 13995 2624 14037 2633
rect 13995 2584 13996 2624
rect 14036 2584 14037 2624
rect 13995 2575 14037 2584
rect 14379 2624 14421 2633
rect 14379 2584 14380 2624
rect 14420 2584 14421 2624
rect 14379 2575 14421 2584
rect 14763 2624 14805 2633
rect 14763 2584 14764 2624
rect 14804 2584 14805 2624
rect 14763 2575 14805 2584
rect 15147 2624 15189 2633
rect 15147 2584 15148 2624
rect 15188 2584 15189 2624
rect 15147 2575 15189 2584
rect 15627 2624 15669 2633
rect 15627 2584 15628 2624
rect 15668 2584 15669 2624
rect 15627 2575 15669 2584
rect 16011 2624 16053 2633
rect 16011 2584 16012 2624
rect 16052 2584 16053 2624
rect 16011 2575 16053 2584
rect 16779 2624 16821 2633
rect 16779 2584 16780 2624
rect 16820 2584 16821 2624
rect 16779 2575 16821 2584
rect 16971 2624 17013 2633
rect 16971 2584 16972 2624
rect 17012 2584 17013 2624
rect 16971 2575 17013 2584
rect 17355 2624 17397 2633
rect 17355 2584 17356 2624
rect 17396 2584 17397 2624
rect 17355 2575 17397 2584
rect 18891 2624 18933 2633
rect 18891 2584 18892 2624
rect 18932 2584 18933 2624
rect 18891 2575 18933 2584
rect 19467 2624 19509 2633
rect 19467 2584 19468 2624
rect 19508 2584 19509 2624
rect 19467 2575 19509 2584
rect 19851 2624 19893 2633
rect 19851 2584 19852 2624
rect 19892 2584 19893 2624
rect 19851 2575 19893 2584
rect 20139 2624 20181 2633
rect 20139 2584 20140 2624
rect 20180 2584 20181 2624
rect 20139 2575 20181 2584
rect 15387 2540 15429 2549
rect 15387 2500 15388 2540
rect 15428 2500 15429 2540
rect 15387 2491 15429 2500
rect 16539 2540 16581 2549
rect 16539 2500 16540 2540
rect 16580 2500 16581 2540
rect 16539 2491 16581 2500
rect 19131 2540 19173 2549
rect 19131 2500 19132 2540
rect 19172 2500 19173 2540
rect 19131 2491 19173 2500
rect 2715 2456 2757 2465
rect 2715 2416 2716 2456
rect 2756 2416 2757 2456
rect 2715 2407 2757 2416
rect 8955 2456 8997 2465
rect 8955 2416 8956 2456
rect 8996 2416 8997 2456
rect 8955 2407 8997 2416
rect 9339 2456 9381 2465
rect 9339 2416 9340 2456
rect 9380 2416 9381 2456
rect 9339 2407 9381 2416
rect 9723 2456 9765 2465
rect 9723 2416 9724 2456
rect 9764 2416 9765 2456
rect 9723 2407 9765 2416
rect 10107 2456 10149 2465
rect 10107 2416 10108 2456
rect 10148 2416 10149 2456
rect 10107 2407 10149 2416
rect 10491 2456 10533 2465
rect 10491 2416 10492 2456
rect 10532 2416 10533 2456
rect 10491 2407 10533 2416
rect 10875 2456 10917 2465
rect 10875 2416 10876 2456
rect 10916 2416 10917 2456
rect 10875 2407 10917 2416
rect 12603 2456 12645 2465
rect 12603 2416 12604 2456
rect 12644 2416 12645 2456
rect 12603 2407 12645 2416
rect 12987 2456 13029 2465
rect 12987 2416 12988 2456
rect 13028 2416 13029 2456
rect 12987 2407 13029 2416
rect 13371 2456 13413 2465
rect 13371 2416 13372 2456
rect 13412 2416 13413 2456
rect 13371 2407 13413 2416
rect 13755 2456 13797 2465
rect 13755 2416 13756 2456
rect 13796 2416 13797 2456
rect 13755 2407 13797 2416
rect 14139 2456 14181 2465
rect 14139 2416 14140 2456
rect 14180 2416 14181 2456
rect 14139 2407 14181 2416
rect 14523 2456 14565 2465
rect 14523 2416 14524 2456
rect 14564 2416 14565 2456
rect 14523 2407 14565 2416
rect 14907 2456 14949 2465
rect 14907 2416 14908 2456
rect 14948 2416 14949 2456
rect 14907 2407 14949 2416
rect 15771 2456 15813 2465
rect 15771 2416 15772 2456
rect 15812 2416 15813 2456
rect 15771 2407 15813 2416
rect 17595 2456 17637 2465
rect 17595 2416 17596 2456
rect 17636 2416 17637 2456
rect 17595 2407 17637 2416
rect 19227 2456 19269 2465
rect 19227 2416 19228 2456
rect 19268 2416 19269 2456
rect 19227 2407 19269 2416
rect 19611 2456 19653 2465
rect 19611 2416 19612 2456
rect 19652 2416 19653 2456
rect 19611 2407 19653 2416
rect 1152 2288 20448 2312
rect 1152 2248 3688 2288
rect 3728 2248 3770 2288
rect 3810 2248 3852 2288
rect 3892 2248 3934 2288
rect 3974 2248 4016 2288
rect 4056 2248 18808 2288
rect 18848 2248 18890 2288
rect 18930 2248 18972 2288
rect 19012 2248 19054 2288
rect 19094 2248 19136 2288
rect 19176 2248 20448 2288
rect 1152 2224 20448 2248
rect 15099 2120 15141 2129
rect 15099 2080 15100 2120
rect 15140 2080 15141 2120
rect 15099 2071 15141 2080
rect 19995 2120 20037 2129
rect 19995 2080 19996 2120
rect 20036 2080 20037 2120
rect 19995 2071 20037 2080
rect 20379 2036 20421 2045
rect 20379 1996 20380 2036
rect 20420 1996 20421 2036
rect 20379 1987 20421 1996
rect 8235 1952 8277 1961
rect 8235 1912 8236 1952
rect 8276 1912 8277 1952
rect 8235 1903 8277 1912
rect 8619 1952 8661 1961
rect 8619 1912 8620 1952
rect 8660 1912 8661 1952
rect 8619 1903 8661 1912
rect 9003 1952 9045 1961
rect 9003 1912 9004 1952
rect 9044 1912 9045 1952
rect 9003 1903 9045 1912
rect 9387 1952 9429 1961
rect 9387 1912 9388 1952
rect 9428 1912 9429 1952
rect 9387 1903 9429 1912
rect 9771 1952 9813 1961
rect 9771 1912 9772 1952
rect 9812 1912 9813 1952
rect 9771 1903 9813 1912
rect 10155 1952 10197 1961
rect 10155 1912 10156 1952
rect 10196 1912 10197 1952
rect 10155 1903 10197 1912
rect 10539 1952 10581 1961
rect 10539 1912 10540 1952
rect 10580 1912 10581 1952
rect 10539 1903 10581 1912
rect 10923 1952 10965 1961
rect 10923 1912 10924 1952
rect 10964 1912 10965 1952
rect 10923 1903 10965 1912
rect 11259 1952 11301 1961
rect 11259 1912 11260 1952
rect 11300 1912 11301 1952
rect 11259 1903 11301 1912
rect 11883 1952 11925 1961
rect 11883 1912 11884 1952
rect 11924 1912 11925 1952
rect 11883 1903 11925 1912
rect 12267 1952 12309 1961
rect 12267 1912 12268 1952
rect 12308 1912 12309 1952
rect 12267 1903 12309 1912
rect 12651 1952 12693 1961
rect 12651 1912 12652 1952
rect 12692 1912 12693 1952
rect 12651 1903 12693 1912
rect 13035 1952 13077 1961
rect 13035 1912 13036 1952
rect 13076 1912 13077 1952
rect 13035 1903 13077 1912
rect 13419 1952 13461 1961
rect 13419 1912 13420 1952
rect 13460 1912 13461 1952
rect 13419 1903 13461 1912
rect 13803 1952 13845 1961
rect 13803 1912 13804 1952
rect 13844 1912 13845 1952
rect 13803 1903 13845 1912
rect 14187 1952 14229 1961
rect 14187 1912 14188 1952
rect 14228 1912 14229 1952
rect 14187 1903 14229 1912
rect 14571 1952 14613 1961
rect 14571 1912 14572 1952
rect 14612 1912 14613 1952
rect 14571 1903 14613 1912
rect 14955 1952 14997 1961
rect 14955 1912 14956 1952
rect 14996 1912 14997 1952
rect 14955 1903 14997 1912
rect 15339 1952 15381 1961
rect 15339 1912 15340 1952
rect 15380 1912 15381 1952
rect 15339 1903 15381 1912
rect 15771 1952 15813 1961
rect 15771 1912 15772 1952
rect 15812 1912 15813 1952
rect 15771 1903 15813 1912
rect 16107 1952 16149 1961
rect 16107 1912 16108 1952
rect 16148 1912 16149 1952
rect 16107 1903 16149 1912
rect 16491 1952 16533 1961
rect 16491 1912 16492 1952
rect 16532 1912 16533 1952
rect 16491 1903 16533 1912
rect 16875 1952 16917 1961
rect 16875 1912 16876 1952
rect 16916 1912 16917 1952
rect 16875 1903 16917 1912
rect 18219 1952 18261 1961
rect 18219 1912 18220 1952
rect 18260 1912 18261 1952
rect 18219 1903 18261 1912
rect 18603 1952 18645 1961
rect 18603 1912 18604 1952
rect 18644 1912 18645 1952
rect 18603 1903 18645 1912
rect 18987 1952 19029 1961
rect 18987 1912 18988 1952
rect 19028 1912 19029 1952
rect 18987 1903 19029 1912
rect 19371 1952 19413 1961
rect 19371 1912 19372 1952
rect 19412 1912 19413 1952
rect 19371 1903 19413 1912
rect 19755 1952 19797 1961
rect 19755 1912 19756 1952
rect 19796 1912 19797 1952
rect 19755 1903 19797 1912
rect 20139 1952 20181 1961
rect 20139 1912 20140 1952
rect 20180 1912 20181 1952
rect 20139 1903 20181 1912
rect 11547 1784 11589 1793
rect 11547 1744 11548 1784
rect 11588 1744 11589 1784
rect 11547 1735 11589 1744
rect 12411 1784 12453 1793
rect 12411 1744 12412 1784
rect 12452 1744 12453 1784
rect 12411 1735 12453 1744
rect 13563 1784 13605 1793
rect 13563 1744 13564 1784
rect 13604 1744 13605 1784
rect 13563 1735 13605 1744
rect 15483 1784 15525 1793
rect 15483 1744 15484 1784
rect 15524 1744 15525 1784
rect 15483 1735 15525 1744
rect 16635 1784 16677 1793
rect 16635 1744 16636 1784
rect 16676 1744 16677 1784
rect 16635 1735 16677 1744
rect 18843 1784 18885 1793
rect 18843 1744 18844 1784
rect 18884 1744 18885 1784
rect 18843 1735 18885 1744
rect 19611 1784 19653 1793
rect 19611 1744 19612 1784
rect 19652 1744 19653 1784
rect 19611 1735 19653 1744
rect 8475 1700 8517 1709
rect 8475 1660 8476 1700
rect 8516 1660 8517 1700
rect 8475 1651 8517 1660
rect 8859 1700 8901 1709
rect 8859 1660 8860 1700
rect 8900 1660 8901 1700
rect 8859 1651 8901 1660
rect 9243 1700 9285 1709
rect 9243 1660 9244 1700
rect 9284 1660 9285 1700
rect 9243 1651 9285 1660
rect 9627 1700 9669 1709
rect 9627 1660 9628 1700
rect 9668 1660 9669 1700
rect 9627 1651 9669 1660
rect 10011 1700 10053 1709
rect 10011 1660 10012 1700
rect 10052 1660 10053 1700
rect 10011 1651 10053 1660
rect 10395 1700 10437 1709
rect 10395 1660 10396 1700
rect 10436 1660 10437 1700
rect 10395 1651 10437 1660
rect 10779 1700 10821 1709
rect 10779 1660 10780 1700
rect 10820 1660 10821 1700
rect 10779 1651 10821 1660
rect 11163 1700 11205 1709
rect 11163 1660 11164 1700
rect 11204 1660 11205 1700
rect 11163 1651 11205 1660
rect 11643 1700 11685 1709
rect 11643 1660 11644 1700
rect 11684 1660 11685 1700
rect 11643 1651 11685 1660
rect 12027 1700 12069 1709
rect 12027 1660 12028 1700
rect 12068 1660 12069 1700
rect 12027 1651 12069 1660
rect 12795 1700 12837 1709
rect 12795 1660 12796 1700
rect 12836 1660 12837 1700
rect 12795 1651 12837 1660
rect 13179 1700 13221 1709
rect 13179 1660 13180 1700
rect 13220 1660 13221 1700
rect 13179 1651 13221 1660
rect 13947 1700 13989 1709
rect 13947 1660 13948 1700
rect 13988 1660 13989 1700
rect 13947 1651 13989 1660
rect 14331 1700 14373 1709
rect 14331 1660 14332 1700
rect 14372 1660 14373 1700
rect 14331 1651 14373 1660
rect 14715 1700 14757 1709
rect 14715 1660 14716 1700
rect 14756 1660 14757 1700
rect 14715 1651 14757 1660
rect 15867 1700 15909 1709
rect 15867 1660 15868 1700
rect 15908 1660 15909 1700
rect 15867 1651 15909 1660
rect 16251 1700 16293 1709
rect 16251 1660 16252 1700
rect 16292 1660 16293 1700
rect 16251 1651 16293 1660
rect 18459 1700 18501 1709
rect 18459 1660 18460 1700
rect 18500 1660 18501 1700
rect 18459 1651 18501 1660
rect 19227 1700 19269 1709
rect 19227 1660 19228 1700
rect 19268 1660 19269 1700
rect 19227 1651 19269 1660
rect 1152 1532 20452 1556
rect 1152 1492 4928 1532
rect 4968 1492 5010 1532
rect 5050 1492 5092 1532
rect 5132 1492 5174 1532
rect 5214 1492 5256 1532
rect 5296 1492 20048 1532
rect 20088 1492 20130 1532
rect 20170 1492 20212 1532
rect 20252 1492 20294 1532
rect 20334 1492 20376 1532
rect 20416 1492 20452 1532
rect 1152 1468 20452 1492
<< via1 >>
rect 4928 10564 4968 10604
rect 5010 10564 5050 10604
rect 5092 10564 5132 10604
rect 5174 10564 5214 10604
rect 5256 10564 5296 10604
rect 20048 10564 20088 10604
rect 20130 10564 20170 10604
rect 20212 10564 20252 10604
rect 20294 10564 20334 10604
rect 20376 10564 20416 10604
rect 1180 10396 1220 10436
rect 2044 10396 2084 10436
rect 3004 10396 3044 10436
rect 3964 10396 4004 10436
rect 4924 10396 4964 10436
rect 5884 10396 5924 10436
rect 6844 10396 6884 10436
rect 7804 10396 7844 10436
rect 8764 10396 8804 10436
rect 9724 10396 9764 10436
rect 10684 10396 10724 10436
rect 11644 10396 11684 10436
rect 12604 10396 12644 10436
rect 13564 10396 13604 10436
rect 14524 10396 14564 10436
rect 15484 10396 15524 10436
rect 16444 10396 16484 10436
rect 17404 10396 17444 10436
rect 18364 10396 18404 10436
rect 19324 10396 19364 10436
rect 18268 10312 18308 10352
rect 1420 10144 1460 10184
rect 2284 10144 2324 10184
rect 3244 10144 3284 10184
rect 4204 10144 4244 10184
rect 5164 10144 5204 10184
rect 6124 10144 6164 10184
rect 7084 10144 7124 10184
rect 8044 10144 8084 10184
rect 9004 10144 9044 10184
rect 9964 10144 10004 10184
rect 10924 10144 10964 10184
rect 11884 10144 11924 10184
rect 12844 10144 12884 10184
rect 13804 10144 13844 10184
rect 14764 10144 14804 10184
rect 15724 10144 15764 10184
rect 16684 10144 16724 10184
rect 17644 10144 17684 10184
rect 18028 10144 18068 10184
rect 18604 10144 18644 10184
rect 18988 10144 19028 10184
rect 19564 10144 19604 10184
rect 19756 10144 19796 10184
rect 20140 10144 20180 10184
rect 19228 9976 19268 10016
rect 19996 9976 20036 10016
rect 20380 9976 20420 10016
rect 3688 9808 3728 9848
rect 3770 9808 3810 9848
rect 3852 9808 3892 9848
rect 3934 9808 3974 9848
rect 4016 9808 4056 9848
rect 18808 9808 18848 9848
rect 18890 9808 18930 9848
rect 18972 9808 19012 9848
rect 19054 9808 19094 9848
rect 19136 9808 19176 9848
rect 2332 9640 2372 9680
rect 10876 9640 10916 9680
rect 13756 9640 13796 9680
rect 14812 9640 14852 9680
rect 16636 9640 16676 9680
rect 18748 9640 18788 9680
rect 19132 9640 19172 9680
rect 14140 9556 14180 9596
rect 2572 9472 2612 9512
rect 11116 9472 11156 9512
rect 11308 9472 11348 9512
rect 11548 9472 11588 9512
rect 13996 9472 14036 9512
rect 14380 9472 14420 9512
rect 15052 9472 15092 9512
rect 16396 9472 16436 9512
rect 17548 9472 17588 9512
rect 18124 9472 18164 9512
rect 18508 9472 18548 9512
rect 18892 9472 18932 9512
rect 19468 9472 19508 9512
rect 19852 9472 19892 9512
rect 20140 9472 20180 9512
rect 17788 9220 17828 9260
rect 18364 9220 18404 9260
rect 19228 9220 19268 9260
rect 19612 9220 19652 9260
rect 20380 9220 20420 9260
rect 4928 9052 4968 9092
rect 5010 9052 5050 9092
rect 5092 9052 5132 9092
rect 5174 9052 5214 9092
rect 5256 9052 5296 9092
rect 20048 9052 20088 9092
rect 20130 9052 20170 9092
rect 20212 9052 20252 9092
rect 20294 9052 20334 9092
rect 20376 9052 20416 9092
rect 9052 8884 9092 8924
rect 12988 8884 13028 8924
rect 13660 8884 13700 8924
rect 15388 8884 15428 8924
rect 19228 8884 19268 8924
rect 19612 8884 19652 8924
rect 17500 8800 17540 8840
rect 1900 8632 1940 8672
rect 2140 8632 2180 8672
rect 8812 8632 8852 8672
rect 13228 8632 13268 8672
rect 13420 8632 13460 8672
rect 13804 8632 13844 8672
rect 14044 8632 14084 8672
rect 15628 8632 15668 8672
rect 17260 8632 17300 8672
rect 18988 8632 19028 8672
rect 19372 8632 19412 8672
rect 19756 8632 19796 8672
rect 19996 8632 20036 8672
rect 20140 8632 20180 8672
rect 20380 8464 20420 8504
rect 3688 8296 3728 8336
rect 3770 8296 3810 8336
rect 3852 8296 3892 8336
rect 3934 8296 3974 8336
rect 4016 8296 4056 8336
rect 18808 8296 18848 8336
rect 18890 8296 18930 8336
rect 18972 8296 19012 8336
rect 19054 8296 19094 8336
rect 19136 8296 19176 8336
rect 1948 8128 1988 8168
rect 6748 8128 6788 8168
rect 8380 8128 8420 8168
rect 15580 8128 15620 8168
rect 15964 8128 16004 8168
rect 7900 8044 7940 8084
rect 2188 7960 2228 8000
rect 4492 7960 4532 8000
rect 6988 7960 7028 8000
rect 7660 7960 7700 8000
rect 8620 7960 8660 8000
rect 9004 7960 9044 8000
rect 9964 7960 10004 8000
rect 15340 7960 15380 8000
rect 15724 7960 15764 8000
rect 17068 7960 17108 8000
rect 17932 7960 17972 8000
rect 19756 7960 19796 8000
rect 20140 7960 20180 8000
rect 9244 7792 9284 7832
rect 17308 7792 17348 7832
rect 19996 7792 20036 7832
rect 4732 7708 4772 7748
rect 10204 7708 10244 7748
rect 18172 7708 18212 7748
rect 20380 7708 20420 7748
rect 4928 7540 4968 7580
rect 5010 7540 5050 7580
rect 5092 7540 5132 7580
rect 5174 7540 5214 7580
rect 5256 7540 5296 7580
rect 20048 7540 20088 7580
rect 20130 7540 20170 7580
rect 20212 7540 20252 7580
rect 20294 7540 20334 7580
rect 20376 7540 20416 7580
rect 2092 7120 2132 7160
rect 4876 7120 4916 7160
rect 5116 7120 5156 7160
rect 7372 7120 7412 7160
rect 7756 7120 7796 7160
rect 7996 7120 8036 7160
rect 15244 7120 15284 7160
rect 15484 7120 15524 7160
rect 19084 7120 19124 7160
rect 19468 7120 19508 7160
rect 19852 7120 19892 7160
rect 20092 7120 20132 7160
rect 19324 7036 19364 7076
rect 2332 6952 2372 6992
rect 7612 6952 7652 6992
rect 19708 6952 19748 6992
rect 3688 6784 3728 6824
rect 3770 6784 3810 6824
rect 3852 6784 3892 6824
rect 3934 6784 3974 6824
rect 4016 6784 4056 6824
rect 18808 6784 18848 6824
rect 18890 6784 18930 6824
rect 18972 6784 19012 6824
rect 19054 6784 19094 6824
rect 19136 6784 19176 6824
rect 2332 6616 2372 6656
rect 20380 6616 20420 6656
rect 2092 6448 2132 6488
rect 3532 6448 3572 6488
rect 5212 6448 5252 6488
rect 5452 6448 5492 6488
rect 6220 6448 6260 6488
rect 8908 6448 8948 6488
rect 9148 6448 9188 6488
rect 9388 6448 9428 6488
rect 12844 6448 12884 6488
rect 14476 6448 14516 6488
rect 16684 6448 16724 6488
rect 17068 6448 17108 6488
rect 19276 6448 19316 6488
rect 19756 6448 19796 6488
rect 20140 6448 20180 6488
rect 6460 6280 6500 6320
rect 19996 6280 20036 6320
rect 3772 6196 3812 6236
rect 9628 6196 9668 6236
rect 13084 6196 13124 6236
rect 14716 6196 14756 6236
rect 16924 6196 16964 6236
rect 17308 6196 17348 6236
rect 19516 6196 19556 6236
rect 4928 6028 4968 6068
rect 5010 6028 5050 6068
rect 5092 6028 5132 6068
rect 5174 6028 5214 6068
rect 5256 6028 5296 6068
rect 20048 6028 20088 6068
rect 20130 6028 20170 6068
rect 20212 6028 20252 6068
rect 20294 6028 20334 6068
rect 20376 6028 20416 6068
rect 20380 5860 20420 5900
rect 19996 5776 20036 5816
rect 1996 5608 2036 5648
rect 2476 5608 2516 5648
rect 2716 5608 2756 5648
rect 4684 5608 4724 5648
rect 9004 5608 9044 5648
rect 15724 5608 15764 5648
rect 16972 5608 17012 5648
rect 18508 5608 18548 5648
rect 18892 5608 18932 5648
rect 19372 5608 19412 5648
rect 19756 5608 19796 5648
rect 20140 5608 20180 5648
rect 4924 5524 4964 5564
rect 2236 5440 2276 5480
rect 9244 5440 9284 5480
rect 15964 5440 16004 5480
rect 17212 5440 17252 5480
rect 18748 5440 18788 5480
rect 19132 5440 19172 5480
rect 19612 5440 19652 5480
rect 3688 5272 3728 5312
rect 3770 5272 3810 5312
rect 3852 5272 3892 5312
rect 3934 5272 3974 5312
rect 4016 5272 4056 5312
rect 18808 5272 18848 5312
rect 18890 5272 18930 5312
rect 18972 5272 19012 5312
rect 19054 5272 19094 5312
rect 19136 5272 19176 5312
rect 19324 5020 19364 5060
rect 4972 4936 5012 4976
rect 8716 4936 8756 4976
rect 9100 4936 9140 4976
rect 17068 4936 17108 4976
rect 18739 4936 18779 4976
rect 19084 4936 19124 4976
rect 19468 4936 19508 4976
rect 20140 4936 20180 4976
rect 20380 4936 20420 4976
rect 8956 4768 8996 4808
rect 18940 4768 18980 4808
rect 5212 4684 5252 4724
rect 9340 4684 9380 4724
rect 17308 4684 17348 4724
rect 19708 4684 19748 4724
rect 4928 4516 4968 4556
rect 5010 4516 5050 4556
rect 5092 4516 5132 4556
rect 5174 4516 5214 4556
rect 5256 4516 5296 4556
rect 20048 4516 20088 4556
rect 20130 4516 20170 4556
rect 20212 4516 20252 4556
rect 20294 4516 20334 4556
rect 20376 4516 20416 4556
rect 10876 4348 10916 4388
rect 3868 4264 3908 4304
rect 6460 4264 6500 4304
rect 20380 4264 20420 4304
rect 2284 4096 2324 4136
rect 3628 4096 3668 4136
rect 6220 4096 6260 4136
rect 10252 4096 10292 4136
rect 10588 4096 10628 4136
rect 11596 4096 11636 4136
rect 11980 4096 12020 4136
rect 13612 4096 13652 4136
rect 14284 4096 14324 4136
rect 14668 4096 14708 4136
rect 16396 4096 16436 4136
rect 17932 4096 17972 4136
rect 19084 4096 19124 4136
rect 19660 4096 19700 4136
rect 20140 4096 20180 4136
rect 11836 4012 11876 4052
rect 19324 4012 19364 4052
rect 2524 3928 2564 3968
rect 10492 3928 10532 3968
rect 12220 3928 12260 3968
rect 13372 3928 13412 3968
rect 14044 3928 14084 3968
rect 14428 3928 14468 3968
rect 16156 3928 16196 3968
rect 17692 3928 17732 3968
rect 19420 3928 19460 3968
rect 3688 3760 3728 3800
rect 3770 3760 3810 3800
rect 3852 3760 3892 3800
rect 3934 3760 3974 3800
rect 4016 3760 4056 3800
rect 18808 3760 18848 3800
rect 18890 3760 18930 3800
rect 18972 3760 19012 3800
rect 19054 3760 19094 3800
rect 19136 3760 19176 3800
rect 20380 3592 20420 3632
rect 6268 3508 6308 3548
rect 19996 3508 20036 3548
rect 2476 3424 2516 3464
rect 6028 3424 6068 3464
rect 15724 3424 15764 3464
rect 17068 3424 17108 3464
rect 18988 3424 19028 3464
rect 19564 3424 19604 3464
rect 19756 3424 19796 3464
rect 20140 3424 20180 3464
rect 19228 3256 19268 3296
rect 2716 3172 2756 3212
rect 15484 3172 15524 3212
rect 16828 3172 16868 3212
rect 19324 3172 19364 3212
rect 4928 3004 4968 3044
rect 5010 3004 5050 3044
rect 5092 3004 5132 3044
rect 5174 3004 5214 3044
rect 5256 3004 5296 3044
rect 20048 3004 20088 3044
rect 20130 3004 20170 3044
rect 20212 3004 20252 3044
rect 20294 3004 20334 3044
rect 20376 3004 20416 3044
rect 17212 2836 17252 2876
rect 20380 2836 20420 2876
rect 2332 2752 2372 2792
rect 2092 2584 2132 2624
rect 2476 2584 2516 2624
rect 9196 2584 9236 2624
rect 9580 2584 9620 2624
rect 9964 2584 10004 2624
rect 10348 2584 10388 2624
rect 10732 2584 10772 2624
rect 11116 2584 11156 2624
rect 12844 2584 12884 2624
rect 13228 2584 13268 2624
rect 13612 2584 13652 2624
rect 13996 2584 14036 2624
rect 14380 2584 14420 2624
rect 14764 2584 14804 2624
rect 15148 2584 15188 2624
rect 15628 2584 15668 2624
rect 16012 2584 16052 2624
rect 16780 2584 16820 2624
rect 16972 2584 17012 2624
rect 17356 2584 17396 2624
rect 18892 2584 18932 2624
rect 19468 2584 19508 2624
rect 19852 2584 19892 2624
rect 20140 2584 20180 2624
rect 15388 2500 15428 2540
rect 16540 2500 16580 2540
rect 19132 2500 19172 2540
rect 2716 2416 2756 2456
rect 8956 2416 8996 2456
rect 9340 2416 9380 2456
rect 9724 2416 9764 2456
rect 10108 2416 10148 2456
rect 10492 2416 10532 2456
rect 10876 2416 10916 2456
rect 12604 2416 12644 2456
rect 12988 2416 13028 2456
rect 13372 2416 13412 2456
rect 13756 2416 13796 2456
rect 14140 2416 14180 2456
rect 14524 2416 14564 2456
rect 14908 2416 14948 2456
rect 15772 2416 15812 2456
rect 17596 2416 17636 2456
rect 19228 2416 19268 2456
rect 19612 2416 19652 2456
rect 3688 2248 3728 2288
rect 3770 2248 3810 2288
rect 3852 2248 3892 2288
rect 3934 2248 3974 2288
rect 4016 2248 4056 2288
rect 18808 2248 18848 2288
rect 18890 2248 18930 2288
rect 18972 2248 19012 2288
rect 19054 2248 19094 2288
rect 19136 2248 19176 2288
rect 15100 2080 15140 2120
rect 19996 2080 20036 2120
rect 20380 1996 20420 2036
rect 8236 1912 8276 1952
rect 8620 1912 8660 1952
rect 9004 1912 9044 1952
rect 9388 1912 9428 1952
rect 9772 1912 9812 1952
rect 10156 1912 10196 1952
rect 10540 1912 10580 1952
rect 10924 1912 10964 1952
rect 11260 1912 11300 1952
rect 11884 1912 11924 1952
rect 12268 1912 12308 1952
rect 12652 1912 12692 1952
rect 13036 1912 13076 1952
rect 13420 1912 13460 1952
rect 13804 1912 13844 1952
rect 14188 1912 14228 1952
rect 14572 1912 14612 1952
rect 14956 1912 14996 1952
rect 15340 1912 15380 1952
rect 15772 1912 15812 1952
rect 16108 1912 16148 1952
rect 16492 1912 16532 1952
rect 16876 1912 16916 1952
rect 18220 1912 18260 1952
rect 18604 1912 18644 1952
rect 18988 1912 19028 1952
rect 19372 1912 19412 1952
rect 19756 1912 19796 1952
rect 20140 1912 20180 1952
rect 11548 1744 11588 1784
rect 12412 1744 12452 1784
rect 13564 1744 13604 1784
rect 15484 1744 15524 1784
rect 16636 1744 16676 1784
rect 18844 1744 18884 1784
rect 19612 1744 19652 1784
rect 8476 1660 8516 1700
rect 8860 1660 8900 1700
rect 9244 1660 9284 1700
rect 9628 1660 9668 1700
rect 10012 1660 10052 1700
rect 10396 1660 10436 1700
rect 10780 1660 10820 1700
rect 11164 1660 11204 1700
rect 11644 1660 11684 1700
rect 12028 1660 12068 1700
rect 12796 1660 12836 1700
rect 13180 1660 13220 1700
rect 13948 1660 13988 1700
rect 14332 1660 14372 1700
rect 14716 1660 14756 1700
rect 15868 1660 15908 1700
rect 16252 1660 16292 1700
rect 18460 1660 18500 1700
rect 19228 1660 19268 1700
rect 4928 1492 4968 1532
rect 5010 1492 5050 1532
rect 5092 1492 5132 1532
rect 5174 1492 5214 1532
rect 5256 1492 5296 1532
rect 20048 1492 20088 1532
rect 20130 1492 20170 1532
rect 20212 1492 20252 1532
rect 20294 1492 20334 1532
rect 20376 1492 20416 1532
<< metal2 >>
rect 0 11192 90 11212
rect 21510 11192 21600 11212
rect 0 11152 1324 11192
rect 1364 11152 1373 11192
rect 19459 11152 19468 11192
rect 19508 11152 21600 11192
rect 0 11132 90 11152
rect 21510 11132 21600 11152
rect 0 10856 90 10876
rect 21510 10856 21600 10876
rect 0 10816 8620 10856
rect 8660 10816 8669 10856
rect 19363 10816 19372 10856
rect 19412 10816 21600 10856
rect 0 10796 90 10816
rect 21510 10796 21600 10816
rect 4919 10564 4928 10604
rect 4968 10564 5010 10604
rect 5050 10564 5092 10604
rect 5132 10564 5174 10604
rect 5214 10564 5256 10604
rect 5296 10564 5305 10604
rect 20039 10564 20048 10604
rect 20088 10564 20130 10604
rect 20170 10564 20212 10604
rect 20252 10564 20294 10604
rect 20334 10564 20376 10604
rect 20416 10564 20425 10604
rect 0 10520 90 10540
rect 21510 10520 21600 10540
rect 0 10480 172 10520
rect 212 10480 221 10520
rect 2659 10480 2668 10520
rect 2708 10480 18068 10520
rect 0 10460 90 10480
rect 1027 10396 1036 10436
rect 1076 10396 1180 10436
rect 1220 10396 1229 10436
rect 1987 10396 1996 10436
rect 2036 10396 2044 10436
rect 2084 10396 2167 10436
rect 2947 10396 2956 10436
rect 2996 10396 3004 10436
rect 3044 10396 3127 10436
rect 3907 10396 3916 10436
rect 3956 10396 3964 10436
rect 4004 10396 4087 10436
rect 4771 10396 4780 10436
rect 4820 10396 4924 10436
rect 4964 10396 4973 10436
rect 5827 10396 5836 10436
rect 5876 10396 5884 10436
rect 5924 10396 6007 10436
rect 6787 10396 6796 10436
rect 6836 10396 6844 10436
rect 6884 10396 6967 10436
rect 7747 10396 7756 10436
rect 7796 10396 7804 10436
rect 7844 10396 7927 10436
rect 8707 10396 8716 10436
rect 8756 10396 8764 10436
rect 8804 10396 8887 10436
rect 9667 10396 9676 10436
rect 9716 10396 9724 10436
rect 9764 10396 9847 10436
rect 10627 10396 10636 10436
rect 10676 10396 10684 10436
rect 10724 10396 10807 10436
rect 11587 10396 11596 10436
rect 11636 10396 11644 10436
rect 11684 10396 11767 10436
rect 12547 10396 12556 10436
rect 12596 10396 12604 10436
rect 12644 10396 12727 10436
rect 13507 10396 13516 10436
rect 13556 10396 13564 10436
rect 13604 10396 13687 10436
rect 14467 10396 14476 10436
rect 14516 10396 14524 10436
rect 14564 10396 14647 10436
rect 15427 10396 15436 10436
rect 15476 10396 15484 10436
rect 15524 10396 15607 10436
rect 16387 10396 16396 10436
rect 16436 10396 16444 10436
rect 16484 10396 16567 10436
rect 17347 10396 17356 10436
rect 17396 10396 17404 10436
rect 17444 10396 17527 10436
rect 172 10312 13420 10352
rect 13460 10312 13469 10352
rect 0 10184 90 10204
rect 172 10184 212 10312
rect 14371 10228 14380 10268
rect 14420 10228 16820 10268
rect 0 10144 212 10184
rect 1289 10144 1420 10184
rect 1460 10144 1469 10184
rect 1987 10144 1996 10184
rect 2036 10144 2284 10184
rect 2324 10144 2333 10184
rect 3113 10144 3244 10184
rect 3284 10144 3293 10184
rect 4073 10144 4204 10184
rect 4244 10144 4253 10184
rect 5155 10144 5164 10184
rect 5204 10144 5356 10184
rect 5396 10144 5405 10184
rect 5539 10144 5548 10184
rect 5588 10144 6124 10184
rect 6164 10144 6173 10184
rect 6953 10144 7084 10184
rect 7124 10144 7133 10184
rect 7913 10144 8044 10184
rect 8084 10144 8093 10184
rect 8227 10144 8236 10184
rect 8276 10144 9004 10184
rect 9044 10144 9053 10184
rect 9833 10144 9964 10184
rect 10004 10144 10013 10184
rect 10793 10144 10924 10184
rect 10964 10144 10973 10184
rect 11875 10144 11884 10184
rect 11924 10144 11933 10184
rect 12835 10144 12844 10184
rect 12884 10144 13516 10184
rect 13556 10144 13565 10184
rect 13673 10144 13804 10184
rect 13844 10144 13853 10184
rect 14633 10144 14764 10184
rect 14804 10144 14813 10184
rect 15593 10144 15724 10184
rect 15764 10144 15773 10184
rect 16675 10144 16684 10184
rect 16724 10144 16733 10184
rect 0 10124 90 10144
rect 11884 10100 11924 10144
rect 16684 10100 16724 10144
rect 11884 10060 13036 10100
rect 13076 10060 13085 10100
rect 15523 10060 15532 10100
rect 15572 10060 16724 10100
rect 16780 10100 16820 10228
rect 18028 10184 18068 10480
rect 19948 10480 21600 10520
rect 18307 10396 18316 10436
rect 18356 10396 18364 10436
rect 18404 10396 18487 10436
rect 19267 10396 19276 10436
rect 19316 10396 19324 10436
rect 19364 10396 19447 10436
rect 19948 10352 19988 10480
rect 21510 10460 21600 10480
rect 18259 10312 18268 10352
rect 18308 10312 19988 10352
rect 18124 10228 19028 10268
rect 16867 10144 16876 10184
rect 16916 10144 17644 10184
rect 17684 10144 17693 10184
rect 18019 10144 18028 10184
rect 18068 10144 18077 10184
rect 18124 10100 18164 10228
rect 18988 10184 19028 10228
rect 20140 10228 20716 10268
rect 20756 10228 20765 10268
rect 20140 10184 20180 10228
rect 21510 10184 21600 10204
rect 18473 10144 18604 10184
rect 18644 10144 18653 10184
rect 18979 10144 18988 10184
rect 19028 10144 19037 10184
rect 19084 10144 19564 10184
rect 19604 10144 19613 10184
rect 19747 10144 19756 10184
rect 19796 10144 19927 10184
rect 20131 10144 20140 10184
rect 20180 10144 20189 10184
rect 20236 10144 21600 10184
rect 19084 10100 19124 10144
rect 20236 10100 20276 10144
rect 21510 10124 21600 10144
rect 16780 10060 18164 10100
rect 18691 10060 18700 10100
rect 18740 10060 19124 10100
rect 19363 10060 19372 10100
rect 19412 10060 20276 10100
rect 7852 9976 16244 10016
rect 19219 9976 19228 10016
rect 19268 9976 19892 10016
rect 19987 9976 19996 10016
rect 20036 9976 20140 10016
rect 20180 9976 20189 10016
rect 20371 9976 20380 10016
rect 20420 9976 20908 10016
rect 20948 9976 20957 10016
rect 0 9848 90 9868
rect 0 9808 3532 9848
rect 3572 9808 3581 9848
rect 3679 9808 3688 9848
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 4056 9808 4065 9848
rect 0 9788 90 9808
rect 1315 9724 1324 9764
rect 1364 9724 2516 9764
rect 2476 9680 2516 9724
rect 7852 9680 7892 9976
rect 16204 9932 16244 9976
rect 11107 9892 11116 9932
rect 11156 9892 15820 9932
rect 15860 9892 15869 9932
rect 16204 9892 19508 9932
rect 14284 9808 18124 9848
rect 18164 9808 18173 9848
rect 18799 9808 18808 9848
rect 18848 9808 18890 9848
rect 18930 9808 18972 9848
rect 19012 9808 19054 9848
rect 19094 9808 19136 9848
rect 19176 9808 19185 9848
rect 13795 9724 13804 9764
rect 13844 9724 13853 9764
rect 13804 9680 13844 9724
rect 1411 9640 1420 9680
rect 1460 9640 2332 9680
rect 2372 9640 2381 9680
rect 2476 9640 7892 9680
rect 10793 9640 10876 9680
rect 10916 9640 10924 9680
rect 10964 9640 10973 9680
rect 13747 9640 13756 9680
rect 13796 9640 13844 9680
rect 8611 9556 8620 9596
rect 8660 9556 11348 9596
rect 13507 9556 13516 9596
rect 13556 9556 14140 9596
rect 14180 9556 14189 9596
rect 0 9512 90 9532
rect 11308 9512 11348 9556
rect 14284 9512 14324 9808
rect 14380 9724 17932 9764
rect 17972 9724 17981 9764
rect 18988 9724 19276 9764
rect 19316 9724 19325 9764
rect 14380 9512 14420 9724
rect 18988 9680 19028 9724
rect 14755 9640 14764 9680
rect 14804 9640 14812 9680
rect 14852 9640 14935 9680
rect 16627 9640 16636 9680
rect 16676 9640 18604 9680
rect 18644 9640 18653 9680
rect 18739 9640 18748 9680
rect 18788 9640 19028 9680
rect 19123 9640 19132 9680
rect 19172 9640 19372 9680
rect 19412 9640 19421 9680
rect 15052 9556 18028 9596
rect 18068 9556 18077 9596
rect 18124 9556 19180 9596
rect 19220 9556 19229 9596
rect 15052 9512 15092 9556
rect 18124 9512 18164 9556
rect 19468 9512 19508 9892
rect 19852 9848 19892 9976
rect 21510 9848 21600 9868
rect 19852 9808 21600 9848
rect 21510 9788 21600 9808
rect 20131 9556 20140 9596
rect 20180 9556 20852 9596
rect 20812 9512 20852 9556
rect 21510 9512 21600 9532
rect 0 9472 2372 9512
rect 2441 9472 2572 9512
rect 2612 9472 2621 9512
rect 10985 9472 11116 9512
rect 11156 9472 11165 9512
rect 11299 9472 11308 9512
rect 11348 9472 11357 9512
rect 11539 9472 11548 9512
rect 11588 9472 13804 9512
rect 13844 9472 13853 9512
rect 13987 9472 13996 9512
rect 14036 9472 14324 9512
rect 14371 9472 14380 9512
rect 14420 9472 14429 9512
rect 15043 9472 15052 9512
rect 15092 9472 15101 9512
rect 16387 9472 16396 9512
rect 16436 9472 17260 9512
rect 17300 9472 17309 9512
rect 17417 9472 17548 9512
rect 17588 9472 17597 9512
rect 18115 9472 18124 9512
rect 18164 9472 18173 9512
rect 18377 9472 18508 9512
rect 18548 9472 18557 9512
rect 18761 9472 18892 9512
rect 18932 9472 18941 9512
rect 19459 9472 19468 9512
rect 19508 9472 19517 9512
rect 19651 9472 19660 9512
rect 19700 9472 19852 9512
rect 19892 9472 19901 9512
rect 20131 9472 20140 9512
rect 20180 9472 20524 9512
rect 20564 9472 20573 9512
rect 20812 9472 21600 9512
rect 0 9452 90 9472
rect 2332 9428 2372 9472
rect 21510 9452 21600 9472
rect 2332 9388 10060 9428
rect 10100 9388 10109 9428
rect 3523 9304 3532 9344
rect 3572 9304 13804 9344
rect 13844 9304 13853 9344
rect 18988 9304 20428 9344
rect 20468 9304 20477 9344
rect 18988 9260 19028 9304
rect 15811 9220 15820 9260
rect 15860 9220 17452 9260
rect 17492 9220 17501 9260
rect 17779 9220 17788 9260
rect 17828 9220 18260 9260
rect 18355 9220 18364 9260
rect 18404 9220 19028 9260
rect 19084 9220 19228 9260
rect 19268 9220 19277 9260
rect 19372 9220 19612 9260
rect 19652 9220 19661 9260
rect 20371 9220 20380 9260
rect 20420 9220 21004 9260
rect 21044 9220 21053 9260
rect 0 9176 90 9196
rect 18220 9176 18260 9220
rect 0 9136 15340 9176
rect 15380 9136 15389 9176
rect 18220 9136 18700 9176
rect 18740 9136 18749 9176
rect 0 9116 90 9136
rect 4919 9052 4928 9092
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 5296 9052 5305 9092
rect 12940 9052 15380 9092
rect 15619 9052 15628 9092
rect 15668 9052 18892 9092
rect 18932 9052 18941 9092
rect 12940 9008 12980 9052
rect 1219 8968 1228 9008
rect 1268 8968 12980 9008
rect 15340 9008 15380 9052
rect 15340 8968 17300 9008
rect 17539 8968 17548 9008
rect 17588 8968 18988 9008
rect 19028 8968 19037 9008
rect 9043 8884 9052 8924
rect 9092 8884 9964 8924
rect 10004 8884 10013 8924
rect 12979 8884 12988 8924
rect 13028 8884 13036 8924
rect 13076 8884 13159 8924
rect 13651 8884 13660 8924
rect 13700 8884 15244 8924
rect 15284 8884 15293 8924
rect 15379 8884 15388 8924
rect 15428 8884 15724 8924
rect 15764 8884 15773 8924
rect 0 8840 90 8860
rect 0 8800 4588 8840
rect 4628 8800 4637 8840
rect 6499 8800 6508 8840
rect 6548 8800 17204 8840
rect 0 8780 90 8800
rect 1900 8716 3340 8756
rect 3380 8716 3389 8756
rect 13228 8716 17068 8756
rect 17108 8716 17117 8756
rect 1900 8672 1940 8716
rect 13228 8672 13268 8716
rect 1891 8632 1900 8672
rect 1940 8632 1949 8672
rect 2131 8632 2140 8672
rect 2180 8632 2284 8672
rect 2324 8632 2333 8672
rect 8681 8632 8716 8672
rect 8756 8632 8812 8672
rect 8852 8632 8861 8672
rect 13219 8632 13228 8672
rect 13268 8632 13277 8672
rect 13411 8632 13420 8672
rect 13460 8632 13591 8672
rect 13673 8632 13804 8672
rect 13844 8632 13853 8672
rect 14035 8632 14044 8672
rect 14084 8632 14380 8672
rect 14420 8632 14429 8672
rect 15619 8632 15628 8672
rect 15668 8632 17108 8672
rect 0 8504 90 8524
rect 17068 8504 17108 8632
rect 17164 8588 17204 8800
rect 17260 8672 17300 8968
rect 17347 8884 17356 8924
rect 17396 8884 19028 8924
rect 18988 8840 19028 8884
rect 17491 8800 17500 8840
rect 17540 8800 18604 8840
rect 18644 8800 18653 8840
rect 18979 8800 18988 8840
rect 19028 8800 19037 8840
rect 17347 8716 17356 8756
rect 17396 8716 17740 8756
rect 17780 8716 17789 8756
rect 18019 8716 18028 8756
rect 18068 8716 18316 8756
rect 18356 8716 18365 8756
rect 19084 8672 19124 9220
rect 19372 9176 19412 9220
rect 21510 9176 21600 9196
rect 19171 9136 19180 9176
rect 19220 9136 19412 9176
rect 20899 9136 20908 9176
rect 20948 9136 21600 9176
rect 21510 9116 21600 9136
rect 20039 9052 20048 9092
rect 20088 9052 20130 9092
rect 20170 9052 20212 9092
rect 20252 9052 20294 9092
rect 20334 9052 20376 9092
rect 20416 9052 20425 9092
rect 19219 8884 19228 8924
rect 19268 8884 19468 8924
rect 19508 8884 19517 8924
rect 19603 8884 19612 8924
rect 19652 8884 19756 8924
rect 19796 8884 19805 8924
rect 21510 8840 21600 8860
rect 19171 8800 19180 8840
rect 19220 8800 19564 8840
rect 19604 8800 19613 8840
rect 20995 8800 21004 8840
rect 21044 8800 21600 8840
rect 21510 8780 21600 8800
rect 17251 8632 17260 8672
rect 17300 8632 17309 8672
rect 17356 8632 18932 8672
rect 18979 8632 18988 8672
rect 19028 8632 19124 8672
rect 19241 8632 19372 8672
rect 19412 8632 19421 8672
rect 19468 8632 19756 8672
rect 19796 8632 19805 8672
rect 19987 8632 19996 8672
rect 20036 8632 20084 8672
rect 20131 8632 20140 8672
rect 20180 8632 20620 8672
rect 20660 8632 20669 8672
rect 17356 8588 17396 8632
rect 17164 8548 17396 8588
rect 18892 8588 18932 8632
rect 19468 8588 19508 8632
rect 18892 8548 19508 8588
rect 20044 8588 20084 8632
rect 20044 8548 20852 8588
rect 20812 8504 20852 8548
rect 21510 8504 21600 8524
rect 0 8464 4108 8504
rect 4148 8464 4157 8504
rect 17068 8464 18412 8504
rect 18452 8464 18461 8504
rect 20371 8464 20380 8504
rect 20420 8464 20429 8504
rect 20812 8464 21600 8504
rect 0 8444 90 8464
rect 20380 8336 20420 8464
rect 21510 8444 21600 8464
rect 3679 8296 3688 8336
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 4056 8296 4065 8336
rect 8620 8296 16780 8336
rect 16820 8296 16829 8336
rect 18799 8296 18808 8336
rect 18848 8296 18890 8336
rect 18930 8296 18972 8336
rect 19012 8296 19054 8336
rect 19094 8296 19136 8336
rect 19176 8296 19185 8336
rect 20380 8296 21044 8336
rect 0 8168 90 8188
rect 0 8128 1708 8168
rect 1748 8128 1757 8168
rect 1865 8128 1948 8168
rect 1988 8128 1996 8168
rect 2036 8128 2045 8168
rect 6739 8128 6748 8168
rect 6788 8128 7084 8168
rect 7124 8128 7133 8168
rect 8035 8128 8044 8168
rect 8084 8128 8380 8168
rect 8420 8128 8429 8168
rect 0 8108 90 8128
rect 7891 8044 7900 8084
rect 7940 8044 8236 8084
rect 8276 8044 8285 8084
rect 8620 8000 8660 8296
rect 15820 8212 20716 8252
rect 20756 8212 20765 8252
rect 15820 8168 15860 8212
rect 21004 8168 21044 8296
rect 21510 8168 21600 8188
rect 15571 8128 15580 8168
rect 15620 8128 15860 8168
rect 15955 8128 15964 8168
rect 16004 8128 16876 8168
rect 16916 8128 16925 8168
rect 17251 8128 17260 8168
rect 17300 8128 20180 8168
rect 21004 8128 21600 8168
rect 15052 8044 19796 8084
rect 2179 7960 2188 8000
rect 2228 7960 2764 8000
rect 2804 7960 2813 8000
rect 4291 7960 4300 8000
rect 4340 7960 4492 8000
rect 4532 7960 4541 8000
rect 6857 7960 6892 8000
rect 6932 7960 6988 8000
rect 7028 7960 7037 8000
rect 7529 7960 7660 8000
rect 7700 7960 7709 8000
rect 8611 7960 8620 8000
rect 8660 7960 8669 8000
rect 8995 7960 9004 8000
rect 9044 7960 9053 8000
rect 9100 7960 9964 8000
rect 10004 7960 10013 8000
rect 9004 7916 9044 7960
rect 4483 7876 4492 7916
rect 4532 7876 9044 7916
rect 0 7832 90 7852
rect 9100 7832 9140 7960
rect 0 7792 3052 7832
rect 3092 7792 3101 7832
rect 4675 7792 4684 7832
rect 4724 7792 9140 7832
rect 9235 7792 9244 7832
rect 9284 7792 12076 7832
rect 12116 7792 12125 7832
rect 0 7772 90 7792
rect 4723 7708 4732 7748
rect 4772 7708 7796 7748
rect 10195 7708 10204 7748
rect 10244 7708 11500 7748
rect 11540 7708 11549 7748
rect 7756 7664 7796 7708
rect 7756 7624 13132 7664
rect 13172 7624 13181 7664
rect 15052 7580 15092 8044
rect 19756 8000 19796 8044
rect 20140 8000 20180 8128
rect 21510 8108 21600 8128
rect 15209 7960 15340 8000
rect 15380 7960 15389 8000
rect 15715 7960 15724 8000
rect 15764 7960 15773 8000
rect 16937 7960 17068 8000
rect 17108 7960 17117 8000
rect 17347 7960 17356 8000
rect 17396 7960 17932 8000
rect 17972 7960 17981 8000
rect 19747 7960 19756 8000
rect 19796 7960 19805 8000
rect 20131 7960 20140 8000
rect 20180 7960 20189 8000
rect 15724 7664 15764 7960
rect 21510 7832 21600 7852
rect 17299 7792 17308 7832
rect 17348 7792 19756 7832
rect 19796 7792 19805 7832
rect 19987 7792 19996 7832
rect 20036 7792 21600 7832
rect 21510 7772 21600 7792
rect 18163 7708 18172 7748
rect 18212 7708 18700 7748
rect 18740 7708 18749 7748
rect 20371 7708 20380 7748
rect 20420 7708 20429 7748
rect 20380 7664 20420 7708
rect 15724 7624 19468 7664
rect 19508 7624 19517 7664
rect 20380 7624 21044 7664
rect 4919 7540 4928 7580
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 5296 7540 5305 7580
rect 6307 7540 6316 7580
rect 6356 7540 15092 7580
rect 20039 7540 20048 7580
rect 20088 7540 20130 7580
rect 20170 7540 20212 7580
rect 20252 7540 20294 7580
rect 20334 7540 20376 7580
rect 20416 7540 20425 7580
rect 0 7496 90 7516
rect 21004 7496 21044 7624
rect 21510 7496 21600 7516
rect 0 7456 12844 7496
rect 12884 7456 12893 7496
rect 21004 7456 21600 7496
rect 0 7436 90 7456
rect 21510 7436 21600 7456
rect 931 7288 940 7328
rect 980 7288 17356 7328
rect 17396 7288 17405 7328
rect 3244 7204 3572 7244
rect 0 7160 90 7180
rect 0 7120 2036 7160
rect 2083 7120 2092 7160
rect 2132 7120 2956 7160
rect 2996 7120 3005 7160
rect 0 7100 90 7120
rect 1996 7076 2036 7120
rect 3244 7076 3284 7204
rect 1996 7036 3284 7076
rect 3532 7076 3572 7204
rect 4588 7204 5780 7244
rect 7651 7204 7660 7244
rect 7700 7204 16972 7244
rect 17012 7204 17021 7244
rect 4588 7160 4628 7204
rect 5740 7160 5780 7204
rect 21510 7160 21600 7180
rect 3619 7120 3628 7160
rect 3668 7120 4628 7160
rect 4745 7120 4876 7160
rect 4916 7120 4925 7160
rect 5107 7120 5116 7160
rect 5156 7120 5548 7160
rect 5588 7120 5597 7160
rect 5740 7120 7372 7160
rect 7412 7120 7421 7160
rect 7625 7120 7756 7160
rect 7796 7120 7805 7160
rect 7987 7120 7996 7160
rect 8036 7120 9004 7160
rect 9044 7120 9053 7160
rect 15113 7120 15244 7160
rect 15284 7120 15293 7160
rect 15401 7120 15484 7160
rect 15524 7120 15532 7160
rect 15572 7120 15581 7160
rect 19075 7120 19084 7160
rect 19124 7120 19133 7160
rect 19180 7120 19468 7160
rect 19508 7120 19517 7160
rect 19721 7120 19852 7160
rect 19892 7120 19901 7160
rect 20083 7120 20092 7160
rect 20132 7120 20524 7160
rect 20564 7120 20573 7160
rect 20803 7120 20812 7160
rect 20852 7120 21600 7160
rect 19084 7076 19124 7120
rect 3532 7036 5452 7076
rect 5492 7036 5501 7076
rect 7468 7036 8180 7076
rect 9187 7036 9196 7076
rect 9236 7036 19124 7076
rect 7468 6992 7508 7036
rect 8140 6992 8180 7036
rect 2323 6952 2332 6992
rect 2372 6952 2381 6992
rect 5731 6952 5740 6992
rect 5780 6952 7508 6992
rect 7603 6952 7612 6992
rect 7652 6952 8084 6992
rect 8140 6952 12980 6992
rect 0 6824 90 6844
rect 0 6784 76 6824
rect 116 6784 125 6824
rect 0 6764 90 6784
rect 2332 6740 2372 6952
rect 8044 6908 8084 6952
rect 12940 6908 12980 6952
rect 19180 6908 19220 7120
rect 21510 7100 21600 7120
rect 19315 7036 19324 7076
rect 19364 7036 20420 7076
rect 19699 6952 19708 6992
rect 19748 6952 19988 6992
rect 8044 6868 9964 6908
rect 10004 6868 10013 6908
rect 10060 6868 10964 6908
rect 12940 6868 19220 6908
rect 10060 6824 10100 6868
rect 3148 6784 3572 6824
rect 3679 6784 3688 6824
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 4056 6784 4065 6824
rect 4579 6784 4588 6824
rect 4628 6784 10100 6824
rect 10924 6824 10964 6868
rect 10924 6784 12980 6824
rect 18799 6784 18808 6824
rect 18848 6784 18890 6824
rect 18930 6784 18972 6824
rect 19012 6784 19054 6824
rect 19094 6784 19136 6824
rect 19176 6784 19185 6824
rect 3148 6740 3188 6784
rect 2332 6700 3188 6740
rect 3532 6656 3572 6784
rect 12940 6740 12980 6784
rect 12940 6700 19852 6740
rect 19892 6700 19901 6740
rect 2323 6616 2332 6656
rect 2372 6616 3244 6656
rect 3284 6616 3293 6656
rect 3532 6616 10732 6656
rect 10772 6616 10781 6656
rect 9091 6532 9100 6572
rect 9140 6532 10636 6572
rect 10676 6532 10685 6572
rect 16396 6532 18796 6572
rect 18836 6532 18845 6572
rect 0 6488 90 6508
rect 16396 6488 16436 6532
rect 19948 6488 19988 6952
rect 20380 6824 20420 7036
rect 21510 6824 21600 6844
rect 20380 6784 21600 6824
rect 21510 6764 21600 6784
rect 20371 6616 20380 6656
rect 20420 6616 20812 6656
rect 20852 6616 20861 6656
rect 21510 6488 21600 6508
rect 0 6448 76 6488
rect 116 6448 125 6488
rect 1961 6448 2092 6488
rect 2132 6448 2141 6488
rect 3139 6448 3148 6488
rect 3188 6448 3532 6488
rect 3572 6448 3581 6488
rect 5081 6448 5164 6488
rect 5204 6448 5212 6488
rect 5252 6448 5261 6488
rect 5321 6448 5452 6488
rect 5492 6448 5501 6488
rect 6211 6448 6220 6488
rect 6260 6448 6269 6488
rect 8777 6448 8908 6488
rect 8948 6448 8957 6488
rect 9139 6448 9148 6488
rect 9188 6448 9196 6488
rect 9236 6448 9319 6488
rect 9379 6448 9388 6488
rect 9428 6448 9559 6488
rect 12713 6448 12844 6488
rect 12884 6448 12893 6488
rect 12940 6448 14476 6488
rect 14516 6448 14525 6488
rect 15235 6448 15244 6488
rect 15284 6448 16436 6488
rect 16553 6448 16684 6488
rect 16724 6448 16733 6488
rect 17059 6448 17068 6488
rect 17108 6448 17117 6488
rect 17347 6448 17356 6488
rect 17396 6448 19276 6488
rect 19316 6448 19325 6488
rect 19625 6448 19756 6488
rect 19796 6448 19805 6488
rect 19948 6448 20140 6488
rect 20180 6448 20189 6488
rect 21292 6448 21600 6488
rect 0 6428 90 6448
rect 6220 6404 6260 6448
rect 12940 6404 12980 6448
rect 3427 6364 3436 6404
rect 3476 6364 6260 6404
rect 11587 6364 11596 6404
rect 11636 6364 12980 6404
rect 17068 6320 17108 6448
rect 21292 6320 21332 6448
rect 21510 6428 21600 6448
rect 6451 6280 6460 6320
rect 6500 6280 7852 6320
rect 7892 6280 7901 6320
rect 10051 6280 10060 6320
rect 10100 6280 17108 6320
rect 19987 6280 19996 6320
rect 20036 6280 21332 6320
rect 3763 6196 3772 6236
rect 3812 6196 7948 6236
rect 7988 6196 7997 6236
rect 9619 6196 9628 6236
rect 9668 6196 11404 6236
rect 11444 6196 11453 6236
rect 13075 6196 13084 6236
rect 13124 6196 14612 6236
rect 14707 6196 14716 6236
rect 14756 6196 16780 6236
rect 16820 6196 16829 6236
rect 16915 6196 16924 6236
rect 16964 6196 17252 6236
rect 17299 6196 17308 6236
rect 17348 6196 19412 6236
rect 19507 6196 19516 6236
rect 19556 6196 20620 6236
rect 20660 6196 20669 6236
rect 0 6152 90 6172
rect 14572 6152 14612 6196
rect 0 6112 1228 6152
rect 1268 6112 1277 6152
rect 14572 6112 17068 6152
rect 17108 6112 17117 6152
rect 0 6092 90 6112
rect 4919 6028 4928 6068
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 5296 6028 5305 6068
rect 9475 6028 9484 6068
rect 9524 6028 16588 6068
rect 16628 6028 16637 6068
rect 3619 5944 3628 5984
rect 3668 5944 7756 5984
rect 7796 5944 7805 5984
rect 7939 5944 7948 5984
rect 7988 5944 9772 5984
rect 9812 5944 9821 5984
rect 5443 5860 5452 5900
rect 5492 5860 16300 5900
rect 16340 5860 16349 5900
rect 0 5816 90 5836
rect 17212 5816 17252 6196
rect 19372 6152 19412 6196
rect 21510 6152 21600 6172
rect 19372 6112 20524 6152
rect 20564 6112 20573 6152
rect 21004 6112 21600 6152
rect 20039 6028 20048 6068
rect 20088 6028 20130 6068
rect 20170 6028 20212 6068
rect 20252 6028 20294 6068
rect 20334 6028 20376 6068
rect 20416 6028 20425 6068
rect 21004 5900 21044 6112
rect 21510 6092 21600 6112
rect 18595 5860 18604 5900
rect 18644 5860 19604 5900
rect 20371 5860 20380 5900
rect 20420 5860 21044 5900
rect 0 5776 16684 5816
rect 16724 5776 16733 5816
rect 17212 5776 19508 5816
rect 0 5756 90 5776
rect 172 5692 11596 5732
rect 11636 5692 11645 5732
rect 13891 5692 13900 5732
rect 13940 5692 17012 5732
rect 18691 5692 18700 5732
rect 18740 5692 19412 5732
rect 172 5648 212 5692
rect 16972 5648 17012 5692
rect 19372 5648 19412 5692
rect 19468 5648 19508 5776
rect 19564 5732 19604 5860
rect 21510 5816 21600 5836
rect 19987 5776 19996 5816
rect 20036 5776 21600 5816
rect 21510 5756 21600 5776
rect 19564 5692 20180 5732
rect 20140 5648 20180 5692
rect 67 5608 76 5648
rect 116 5608 212 5648
rect 1987 5608 1996 5648
rect 2036 5608 2188 5648
rect 2228 5608 2237 5648
rect 2467 5608 2476 5648
rect 2516 5608 2525 5648
rect 2659 5608 2668 5648
rect 2708 5608 2716 5648
rect 2756 5608 2839 5648
rect 3331 5608 3340 5648
rect 3380 5608 4684 5648
rect 4724 5608 4733 5648
rect 4780 5608 9004 5648
rect 9044 5608 9053 5648
rect 13699 5608 13708 5648
rect 13748 5608 15724 5648
rect 15764 5608 15773 5648
rect 16963 5608 16972 5648
rect 17012 5608 17021 5648
rect 18377 5608 18508 5648
rect 18548 5608 18557 5648
rect 18883 5608 18892 5648
rect 18932 5608 19063 5648
rect 19363 5608 19372 5648
rect 19412 5608 19421 5648
rect 19468 5608 19756 5648
rect 19796 5608 19805 5648
rect 20131 5608 20140 5648
rect 20180 5608 20189 5648
rect 2476 5564 2516 5608
rect 4780 5564 4820 5608
rect 163 5524 172 5564
rect 212 5524 2516 5564
rect 4771 5524 4780 5564
rect 4820 5524 4829 5564
rect 4915 5524 4924 5564
rect 4964 5524 9484 5564
rect 9524 5524 9533 5564
rect 0 5480 90 5500
rect 21510 5480 21600 5500
rect 0 5440 76 5480
rect 116 5440 125 5480
rect 2227 5440 2236 5480
rect 2276 5440 2900 5480
rect 9235 5440 9244 5480
rect 9284 5440 11212 5480
rect 11252 5440 11261 5480
rect 15955 5440 15964 5480
rect 16004 5440 17108 5480
rect 17203 5440 17212 5480
rect 17252 5440 18220 5480
rect 18260 5440 18269 5480
rect 18700 5440 18748 5480
rect 18788 5440 18797 5480
rect 19123 5440 19132 5480
rect 19172 5440 19276 5480
rect 19316 5440 19325 5480
rect 19603 5440 19612 5480
rect 19652 5440 20564 5480
rect 21475 5440 21484 5480
rect 21524 5440 21600 5480
rect 0 5420 90 5440
rect 2860 5396 2900 5440
rect 17068 5396 17108 5440
rect 2860 5356 9196 5396
rect 9236 5356 9245 5396
rect 17068 5356 18604 5396
rect 18644 5356 18653 5396
rect 3679 5272 3688 5312
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 4056 5272 4065 5312
rect 7939 5272 7948 5312
rect 7988 5272 10060 5312
rect 10100 5272 10109 5312
rect 1123 5188 1132 5228
rect 1172 5188 14476 5228
rect 14516 5188 14525 5228
rect 0 5144 90 5164
rect 0 5104 940 5144
rect 980 5104 989 5144
rect 5443 5104 5452 5144
rect 5492 5104 8852 5144
rect 0 5084 90 5104
rect 5347 5020 5356 5060
rect 5396 5020 8756 5060
rect 8716 4976 8756 5020
rect 8812 4976 8852 5104
rect 18700 4976 18740 5440
rect 18799 5272 18808 5312
rect 18848 5272 18890 5312
rect 18930 5272 18972 5312
rect 19012 5272 19054 5312
rect 19094 5272 19136 5312
rect 19176 5272 19185 5312
rect 20524 5144 20564 5440
rect 21510 5420 21600 5440
rect 21510 5144 21600 5164
rect 20524 5104 21600 5144
rect 21510 5084 21600 5104
rect 19315 5020 19324 5060
rect 19364 5020 20620 5060
rect 20660 5020 20669 5060
rect 2371 4936 2380 4976
rect 2420 4936 4972 4976
rect 5012 4936 5021 4976
rect 7756 4936 7988 4976
rect 8707 4936 8716 4976
rect 8756 4936 8765 4976
rect 8812 4936 9100 4976
rect 9140 4936 9149 4976
rect 14371 4936 14380 4976
rect 14420 4936 17068 4976
rect 17108 4936 17117 4976
rect 18700 4936 18739 4976
rect 18779 4936 18788 4976
rect 18953 4936 19084 4976
rect 19124 4936 19133 4976
rect 19459 4936 19468 4976
rect 19508 4936 19517 4976
rect 19843 4936 19852 4976
rect 19892 4936 20140 4976
rect 20180 4936 20189 4976
rect 20371 4936 20380 4976
rect 20420 4936 21484 4976
rect 21524 4936 21533 4976
rect 7756 4892 7796 4936
rect 1411 4852 1420 4892
rect 1460 4852 7796 4892
rect 7948 4892 7988 4936
rect 19468 4892 19508 4936
rect 7948 4852 19508 4892
rect 0 4808 90 4828
rect 21510 4808 21600 4828
rect 0 4768 7948 4808
rect 7988 4768 7997 4808
rect 8947 4768 8956 4808
rect 8996 4768 10924 4808
rect 10964 4768 10973 4808
rect 18931 4768 18940 4808
rect 18980 4768 20564 4808
rect 21283 4768 21292 4808
rect 21332 4768 21600 4808
rect 0 4748 90 4768
rect 5203 4684 5212 4724
rect 5252 4684 8236 4724
rect 8276 4684 8285 4724
rect 9331 4684 9340 4724
rect 9380 4684 10540 4724
rect 10580 4684 10589 4724
rect 17299 4684 17308 4724
rect 17348 4684 18796 4724
rect 18836 4684 18845 4724
rect 19699 4684 19708 4724
rect 19748 4684 19988 4724
rect 1315 4600 1324 4640
rect 1364 4600 19084 4640
rect 19124 4600 19133 4640
rect 4919 4516 4928 4556
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 5296 4516 5305 4556
rect 16771 4516 16780 4556
rect 16820 4516 19852 4556
rect 19892 4516 19901 4556
rect 0 4472 90 4492
rect 0 4432 18508 4472
rect 18548 4432 18557 4472
rect 0 4412 90 4432
rect 19948 4388 19988 4684
rect 20039 4516 20048 4556
rect 20088 4516 20130 4556
rect 20170 4516 20212 4556
rect 20252 4516 20294 4556
rect 20334 4516 20376 4556
rect 20416 4516 20425 4556
rect 20524 4472 20564 4768
rect 21510 4748 21600 4768
rect 21510 4472 21600 4492
rect 20524 4432 21600 4472
rect 21510 4412 21600 4432
rect 10867 4348 10876 4388
rect 10916 4348 14668 4388
rect 14708 4348 14717 4388
rect 18211 4348 18220 4388
rect 18260 4348 19852 4388
rect 19892 4348 19901 4388
rect 19948 4348 20140 4388
rect 20180 4348 20189 4388
rect 3859 4264 3868 4304
rect 3908 4264 4204 4304
rect 4244 4264 4253 4304
rect 6377 4264 6460 4304
rect 6500 4264 6508 4304
rect 6548 4264 6557 4304
rect 7363 4264 7372 4304
rect 7412 4264 10820 4304
rect 20371 4264 20380 4304
rect 20420 4264 21292 4304
rect 21332 4264 21341 4304
rect 3628 4180 10156 4220
rect 10196 4180 10205 4220
rect 0 4136 90 4156
rect 3628 4136 3668 4180
rect 10780 4136 10820 4264
rect 12931 4180 12940 4220
rect 12980 4180 19700 4220
rect 19660 4136 19700 4180
rect 20140 4180 20524 4220
rect 20564 4180 20573 4220
rect 20140 4136 20180 4180
rect 21510 4136 21600 4156
rect 0 4096 1420 4136
rect 1460 4096 1469 4136
rect 2275 4096 2284 4136
rect 2324 4096 2764 4136
rect 2804 4096 2813 4136
rect 3619 4096 3628 4136
rect 3668 4096 3677 4136
rect 4099 4096 4108 4136
rect 4148 4096 6220 4136
rect 6260 4096 6269 4136
rect 7747 4096 7756 4136
rect 7796 4096 10252 4136
rect 10292 4096 10301 4136
rect 10444 4096 10588 4136
rect 10628 4096 10637 4136
rect 10780 4096 11596 4136
rect 11636 4096 11645 4136
rect 11849 4096 11980 4136
rect 12020 4096 12029 4136
rect 12163 4096 12172 4136
rect 12212 4096 13612 4136
rect 13652 4096 13661 4136
rect 14153 4096 14284 4136
rect 14324 4096 14333 4136
rect 14659 4096 14668 4136
rect 14708 4096 14717 4136
rect 16387 4096 16396 4136
rect 16436 4096 16492 4136
rect 16532 4096 16567 4136
rect 16675 4096 16684 4136
rect 16724 4096 17932 4136
rect 17972 4096 17981 4136
rect 18787 4096 18796 4136
rect 18836 4096 19084 4136
rect 19124 4096 19133 4136
rect 19651 4096 19660 4136
rect 19700 4096 19709 4136
rect 20131 4096 20140 4136
rect 20180 4096 20189 4136
rect 20419 4096 20428 4136
rect 20468 4096 21600 4136
rect 0 4076 90 4096
rect 10444 4052 10484 4096
rect 5827 4012 5836 4052
rect 5876 4012 6644 4052
rect 7555 4012 7564 4052
rect 7604 4012 10484 4052
rect 11827 4012 11836 4052
rect 11876 4012 13996 4052
rect 14036 4012 14045 4052
rect 6604 3968 6644 4012
rect 2515 3928 2524 3968
rect 2564 3928 2900 3968
rect 6604 3928 10348 3968
rect 10388 3928 10397 3968
rect 10483 3928 10492 3968
rect 10532 3928 10772 3968
rect 12211 3928 12220 3968
rect 12260 3928 13036 3968
rect 13076 3928 13085 3968
rect 13219 3928 13228 3968
rect 13268 3928 13372 3968
rect 13412 3928 13421 3968
rect 13795 3928 13804 3968
rect 13844 3928 14044 3968
rect 14084 3928 14093 3968
rect 14179 3928 14188 3968
rect 14228 3928 14428 3968
rect 14468 3928 14477 3968
rect 2860 3884 2900 3928
rect 10732 3884 10772 3928
rect 2860 3844 8620 3884
rect 8660 3844 8669 3884
rect 10732 3844 13612 3884
rect 13652 3844 13661 3884
rect 0 3800 90 3820
rect 14668 3800 14708 4096
rect 21510 4076 21600 4096
rect 19315 4012 19324 4052
rect 19364 4012 20468 4052
rect 15811 3928 15820 3968
rect 15860 3928 16156 3968
rect 16196 3928 16205 3968
rect 17347 3928 17356 3968
rect 17396 3928 17692 3968
rect 17732 3928 17741 3968
rect 18211 3928 18220 3968
rect 18260 3928 19420 3968
rect 19460 3928 19469 3968
rect 20428 3800 20468 4012
rect 21510 3800 21600 3820
rect 0 3760 2900 3800
rect 3679 3760 3688 3800
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 4056 3760 4065 3800
rect 8515 3760 8524 3800
rect 8564 3760 14708 3800
rect 18799 3760 18808 3800
rect 18848 3760 18890 3800
rect 18930 3760 18972 3800
rect 19012 3760 19054 3800
rect 19094 3760 19136 3800
rect 19176 3760 19185 3800
rect 20428 3760 21600 3800
rect 0 3740 90 3760
rect 2860 3716 2900 3760
rect 21510 3740 21600 3760
rect 2860 3676 14380 3716
rect 14420 3676 14429 3716
rect 2860 3592 13708 3632
rect 13748 3592 13757 3632
rect 20297 3592 20380 3632
rect 20420 3592 20428 3632
rect 20468 3592 20477 3632
rect 2860 3548 2900 3592
rect 2188 3508 2900 3548
rect 6185 3508 6268 3548
rect 6308 3508 6316 3548
rect 6356 3508 6365 3548
rect 7939 3508 7948 3548
rect 7988 3508 11980 3548
rect 12020 3508 12029 3548
rect 12940 3508 19604 3548
rect 19987 3508 19996 3548
rect 20036 3508 20852 3548
rect 0 3464 90 3484
rect 2188 3464 2228 3508
rect 12940 3464 12980 3508
rect 19564 3464 19604 3508
rect 20812 3464 20852 3508
rect 21510 3464 21600 3484
rect 0 3424 2228 3464
rect 2345 3424 2476 3464
rect 2516 3424 2525 3464
rect 3043 3424 3052 3464
rect 3092 3424 6028 3464
rect 6068 3424 6077 3464
rect 6124 3424 12980 3464
rect 15715 3424 15724 3464
rect 15764 3424 15773 3464
rect 16937 3424 17068 3464
rect 17108 3424 17117 3464
rect 18979 3424 18988 3464
rect 19028 3424 19276 3464
rect 19316 3424 19325 3464
rect 19555 3424 19564 3464
rect 19604 3424 19613 3464
rect 19747 3424 19756 3464
rect 19796 3424 19805 3464
rect 20009 3424 20140 3464
rect 20180 3424 20189 3464
rect 20812 3424 21600 3464
rect 0 3404 90 3424
rect 6124 3380 6164 3424
rect 5635 3340 5644 3380
rect 5684 3340 6164 3380
rect 6211 3340 6220 3380
rect 6260 3340 10060 3380
rect 10100 3340 10109 3380
rect 15724 3296 15764 3424
rect 19756 3380 19796 3424
rect 21510 3404 21600 3424
rect 18595 3340 18604 3380
rect 18644 3340 19796 3380
rect 6979 3256 6988 3296
rect 7028 3256 15764 3296
rect 19219 3256 19228 3296
rect 19268 3256 21004 3296
rect 21044 3256 21053 3296
rect 2707 3172 2716 3212
rect 2756 3172 7180 3212
rect 7220 3172 7229 3212
rect 8131 3172 8140 3212
rect 8180 3172 12172 3212
rect 12212 3172 12221 3212
rect 14371 3172 14380 3212
rect 14420 3172 15484 3212
rect 15524 3172 15533 3212
rect 15907 3172 15916 3212
rect 15956 3172 16828 3212
rect 16868 3172 16877 3212
rect 17443 3172 17452 3212
rect 17492 3172 19324 3212
rect 19364 3172 19373 3212
rect 0 3128 90 3148
rect 21510 3128 21600 3148
rect 0 3088 13900 3128
rect 13940 3088 13949 3128
rect 21004 3088 21600 3128
rect 0 3068 90 3088
rect 4919 3004 4928 3044
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 5296 3004 5305 3044
rect 6019 3004 6028 3044
rect 6068 3004 7316 3044
rect 8419 3004 8428 3044
rect 8468 3004 14284 3044
rect 14324 3004 14333 3044
rect 20039 3004 20048 3044
rect 20088 3004 20130 3044
rect 20170 3004 20212 3044
rect 20252 3004 20294 3044
rect 20334 3004 20376 3044
rect 20416 3004 20425 3044
rect 7276 2960 7316 3004
rect 7084 2920 7180 2960
rect 7220 2920 7229 2960
rect 7276 2920 16684 2960
rect 16724 2920 16733 2960
rect 7084 2876 7124 2920
rect 21004 2876 21044 3088
rect 21510 3068 21600 3088
rect 7084 2836 11156 2876
rect 17203 2836 17212 2876
rect 17252 2836 18604 2876
rect 18644 2836 18653 2876
rect 20371 2836 20380 2876
rect 20420 2836 21044 2876
rect 0 2792 90 2812
rect 0 2752 1132 2792
rect 1172 2752 1181 2792
rect 2323 2752 2332 2792
rect 2372 2752 9100 2792
rect 9140 2752 9149 2792
rect 0 2732 90 2752
rect 2275 2668 2284 2708
rect 2324 2668 7220 2708
rect 9475 2668 9484 2708
rect 9524 2668 10388 2708
rect 7180 2624 7220 2668
rect 10348 2624 10388 2668
rect 11116 2624 11156 2836
rect 21510 2792 21600 2812
rect 17251 2752 17260 2792
rect 17300 2752 19892 2792
rect 20995 2752 21004 2792
rect 21044 2752 21600 2792
rect 12844 2668 14188 2708
rect 14228 2668 14237 2708
rect 15148 2668 15916 2708
rect 15956 2668 15965 2708
rect 12844 2624 12884 2668
rect 15148 2624 15188 2668
rect 19852 2624 19892 2752
rect 21510 2732 21600 2752
rect 19939 2668 19948 2708
rect 19988 2668 19997 2708
rect 19948 2624 19988 2668
rect 1795 2584 1804 2624
rect 1844 2584 2092 2624
rect 2132 2584 2141 2624
rect 2467 2584 2476 2624
rect 2516 2584 2525 2624
rect 7180 2584 8812 2624
rect 8852 2584 8861 2624
rect 9065 2584 9196 2624
rect 9236 2584 9245 2624
rect 9449 2584 9580 2624
rect 9620 2584 9629 2624
rect 9833 2584 9964 2624
rect 10004 2584 10013 2624
rect 10339 2584 10348 2624
rect 10388 2584 10397 2624
rect 10601 2584 10732 2624
rect 10772 2584 10781 2624
rect 11107 2584 11116 2624
rect 11156 2584 11165 2624
rect 12835 2584 12844 2624
rect 12884 2584 12893 2624
rect 13097 2584 13228 2624
rect 13268 2584 13277 2624
rect 13481 2584 13612 2624
rect 13652 2584 13661 2624
rect 13865 2584 13996 2624
rect 14036 2584 14045 2624
rect 14249 2584 14380 2624
rect 14420 2584 14429 2624
rect 14755 2584 14764 2624
rect 14804 2584 14813 2624
rect 15139 2584 15148 2624
rect 15188 2584 15197 2624
rect 15427 2584 15436 2624
rect 15476 2584 15628 2624
rect 15668 2584 15677 2624
rect 15881 2584 16012 2624
rect 16052 2584 16061 2624
rect 16649 2584 16780 2624
rect 16820 2584 16829 2624
rect 16963 2584 16972 2624
rect 17012 2584 17021 2624
rect 17347 2584 17356 2624
rect 17396 2584 17405 2624
rect 18761 2584 18892 2624
rect 18932 2584 18941 2624
rect 19337 2584 19372 2624
rect 19412 2584 19468 2624
rect 19508 2584 19517 2624
rect 19843 2584 19852 2624
rect 19892 2584 19901 2624
rect 19948 2584 20140 2624
rect 20180 2584 20189 2624
rect 2476 2540 2516 2584
rect 14764 2540 14804 2584
rect 1987 2500 1996 2540
rect 2036 2500 2516 2540
rect 7651 2500 7660 2540
rect 7700 2500 11692 2540
rect 11732 2500 11741 2540
rect 11875 2500 11884 2540
rect 11924 2500 14708 2540
rect 14764 2500 15388 2540
rect 15428 2500 15437 2540
rect 15619 2500 15628 2540
rect 15668 2500 16540 2540
rect 16580 2500 16589 2540
rect 0 2456 90 2476
rect 0 2416 1324 2456
rect 1364 2416 1373 2456
rect 2707 2416 2716 2456
rect 2756 2416 8044 2456
rect 8084 2416 8093 2456
rect 8825 2416 8908 2456
rect 8948 2416 8956 2456
rect 8996 2416 9005 2456
rect 9209 2416 9292 2456
rect 9332 2416 9340 2456
rect 9380 2416 9389 2456
rect 9593 2416 9676 2456
rect 9716 2416 9724 2456
rect 9764 2416 9773 2456
rect 9977 2416 10060 2456
rect 10100 2416 10108 2456
rect 10148 2416 10157 2456
rect 10361 2416 10444 2456
rect 10484 2416 10492 2456
rect 10532 2416 10541 2456
rect 10745 2416 10828 2456
rect 10868 2416 10876 2456
rect 10916 2416 10925 2456
rect 12473 2416 12556 2456
rect 12596 2416 12604 2456
rect 12644 2416 12653 2456
rect 12979 2416 12988 2456
rect 13028 2416 13036 2456
rect 13076 2416 13159 2456
rect 13241 2416 13324 2456
rect 13364 2416 13372 2456
rect 13412 2416 13421 2456
rect 13625 2416 13708 2456
rect 13748 2416 13756 2456
rect 13796 2416 13805 2456
rect 14009 2416 14092 2456
rect 14132 2416 14140 2456
rect 14180 2416 14189 2456
rect 14393 2416 14476 2456
rect 14516 2416 14524 2456
rect 14564 2416 14573 2456
rect 0 2396 90 2416
rect 14668 2372 14708 2500
rect 16972 2456 17012 2584
rect 14777 2416 14860 2456
rect 14900 2416 14908 2456
rect 14948 2416 14957 2456
rect 15641 2416 15724 2456
rect 15764 2416 15772 2456
rect 15812 2416 15821 2456
rect 15907 2416 15916 2456
rect 15956 2416 17012 2456
rect 1411 2332 1420 2372
rect 1460 2332 8332 2372
rect 8372 2332 8381 2372
rect 8620 2332 11980 2372
rect 12020 2332 12029 2372
rect 12163 2332 12172 2372
rect 12212 2332 14572 2372
rect 14612 2332 14621 2372
rect 14668 2332 15340 2372
rect 15380 2332 15389 2372
rect 8620 2288 8660 2332
rect 3679 2248 3688 2288
rect 3728 2248 3770 2288
rect 3810 2248 3852 2288
rect 3892 2248 3934 2288
rect 3974 2248 4016 2288
rect 4056 2248 4065 2288
rect 6787 2248 6796 2288
rect 6836 2248 8660 2288
rect 8812 2248 15436 2288
rect 15476 2248 15485 2288
rect 8812 2204 8852 2248
rect 17356 2204 17396 2584
rect 19123 2500 19132 2540
rect 19172 2500 19796 2540
rect 17587 2416 17596 2456
rect 17636 2416 18548 2456
rect 19219 2416 19228 2456
rect 19268 2416 19277 2456
rect 19468 2416 19612 2456
rect 19652 2416 19661 2456
rect 6595 2164 6604 2204
rect 6644 2164 8852 2204
rect 9091 2164 9100 2204
rect 9140 2164 17396 2204
rect 0 2120 90 2140
rect 0 2080 7660 2120
rect 7700 2080 7709 2120
rect 8803 2080 8812 2120
rect 8852 2080 13460 2120
rect 14371 2080 14380 2120
rect 14420 2080 15100 2120
rect 15140 2080 15149 2120
rect 15331 2080 15340 2120
rect 15380 2080 17260 2120
rect 17300 2080 17309 2120
rect 0 2060 90 2080
rect 7843 1996 7852 2036
rect 7892 1996 9428 2036
rect 11491 1996 11500 2036
rect 11540 1996 12692 2036
rect 9388 1952 9428 1996
rect 12652 1952 12692 1996
rect 13420 1952 13460 2080
rect 13507 1996 13516 2036
rect 13556 1996 14228 2036
rect 15715 1996 15724 2036
rect 15764 1996 15773 2036
rect 16108 1996 17356 2036
rect 17396 1996 17405 2036
rect 18124 1996 18220 2036
rect 18260 1996 18269 2036
rect 14188 1952 14228 1996
rect 15724 1952 15764 1996
rect 16108 1952 16148 1996
rect 8105 1912 8236 1952
rect 8276 1912 8285 1952
rect 8419 1912 8428 1952
rect 8468 1912 8620 1952
rect 8660 1912 8669 1952
rect 8873 1912 9004 1952
rect 9044 1912 9053 1952
rect 9379 1912 9388 1952
rect 9428 1912 9437 1952
rect 9641 1912 9772 1952
rect 9812 1912 9821 1952
rect 10147 1912 10156 1952
rect 10196 1912 10205 1952
rect 10409 1912 10540 1952
rect 10580 1912 10589 1952
rect 10793 1912 10924 1952
rect 10964 1912 10973 1952
rect 11129 1912 11212 1952
rect 11252 1912 11260 1952
rect 11300 1912 11309 1952
rect 11395 1912 11404 1952
rect 11444 1912 11884 1952
rect 11924 1912 11933 1952
rect 12067 1912 12076 1952
rect 12116 1912 12268 1952
rect 12308 1912 12317 1952
rect 12643 1912 12652 1952
rect 12692 1912 12701 1952
rect 13027 1912 13036 1952
rect 13076 1912 13132 1952
rect 13172 1912 13207 1952
rect 13411 1912 13420 1952
rect 13460 1912 13469 1952
rect 13673 1912 13804 1952
rect 13844 1912 13853 1952
rect 14179 1912 14188 1952
rect 14228 1912 14237 1952
rect 14537 1912 14572 1952
rect 14612 1912 14668 1952
rect 14708 1912 14717 1952
rect 14947 1912 14956 1952
rect 14996 1912 15005 1952
rect 15331 1912 15340 1952
rect 15380 1912 15628 1952
rect 15668 1912 15677 1952
rect 15724 1912 15772 1952
rect 15812 1912 15821 1952
rect 16099 1912 16108 1952
rect 16148 1912 16157 1952
rect 16483 1912 16492 1952
rect 16532 1912 16541 1952
rect 16867 1912 16876 1952
rect 16916 1912 17452 1952
rect 17492 1912 17501 1952
rect 10156 1868 10196 1912
rect 14956 1868 14996 1912
rect 16492 1868 16532 1912
rect 18124 1868 18164 1996
rect 18508 1952 18548 2416
rect 18799 2248 18808 2288
rect 18848 2248 18890 2288
rect 18930 2248 18972 2288
rect 19012 2248 19054 2288
rect 19094 2248 19136 2288
rect 19176 2248 19185 2288
rect 19228 2120 19268 2416
rect 19084 2080 19268 2120
rect 18595 1996 18604 2036
rect 18644 1996 19028 2036
rect 18988 1952 19028 1996
rect 18211 1912 18220 1952
rect 18260 1912 18269 1952
rect 18508 1912 18604 1952
rect 18644 1912 18653 1952
rect 18979 1912 18988 1952
rect 19028 1912 19037 1952
rect 6403 1828 6412 1868
rect 6452 1828 8564 1868
rect 8611 1828 8620 1868
rect 8660 1828 10196 1868
rect 10252 1828 12172 1868
rect 12212 1828 12221 1868
rect 14956 1828 15820 1868
rect 15860 1828 15869 1868
rect 16492 1828 18164 1868
rect 18220 1868 18260 1912
rect 19084 1868 19124 2080
rect 19468 1952 19508 2416
rect 19756 1952 19796 2500
rect 21510 2456 21600 2476
rect 20419 2416 20428 2456
rect 20468 2416 21600 2456
rect 21510 2396 21600 2416
rect 21510 2120 21600 2140
rect 19987 2080 19996 2120
rect 20036 2080 21600 2120
rect 21510 2060 21600 2080
rect 20297 1996 20380 2036
rect 20420 1996 20428 2036
rect 20468 1996 20477 2036
rect 19363 1912 19372 1952
rect 19412 1912 19508 1952
rect 19747 1912 19756 1952
rect 19796 1912 19805 1952
rect 20131 1912 20140 1952
rect 20180 1912 20620 1952
rect 20660 1912 20669 1952
rect 18220 1828 19124 1868
rect 0 1784 90 1804
rect 8524 1784 8564 1828
rect 10252 1784 10292 1828
rect 21510 1784 21600 1804
rect 0 1744 8372 1784
rect 8524 1744 10292 1784
rect 11395 1744 11404 1784
rect 11444 1744 11548 1784
rect 11588 1744 11597 1784
rect 11779 1744 11788 1784
rect 11828 1744 12412 1784
rect 12452 1744 12461 1784
rect 12739 1744 12748 1784
rect 12788 1744 13564 1784
rect 13604 1744 13613 1784
rect 14659 1744 14668 1784
rect 14708 1744 15484 1784
rect 15524 1744 15533 1784
rect 15619 1744 15628 1784
rect 15668 1744 16636 1784
rect 16676 1744 16685 1784
rect 18835 1744 18844 1784
rect 18884 1744 19180 1784
rect 19220 1744 19229 1784
rect 19603 1744 19612 1784
rect 19652 1744 21600 1784
rect 0 1724 90 1744
rect 8332 1616 8372 1744
rect 21510 1724 21600 1744
rect 8467 1660 8476 1700
rect 8516 1660 8716 1700
rect 8756 1660 8765 1700
rect 8851 1660 8860 1700
rect 8900 1660 9100 1700
rect 9140 1660 9149 1700
rect 9235 1660 9244 1700
rect 9284 1660 9484 1700
rect 9524 1660 9533 1700
rect 9619 1660 9628 1700
rect 9668 1660 9868 1700
rect 9908 1660 9917 1700
rect 10003 1660 10012 1700
rect 10052 1660 10252 1700
rect 10292 1660 10301 1700
rect 10387 1660 10396 1700
rect 10436 1660 10636 1700
rect 10676 1660 10685 1700
rect 10771 1660 10780 1700
rect 10820 1660 11020 1700
rect 11060 1660 11069 1700
rect 11155 1660 11164 1700
rect 11204 1660 11212 1700
rect 11252 1660 11335 1700
rect 11513 1660 11596 1700
rect 11636 1660 11644 1700
rect 11684 1660 11693 1700
rect 11897 1660 11980 1700
rect 12020 1660 12028 1700
rect 12068 1660 12077 1700
rect 12163 1660 12172 1700
rect 12212 1660 12796 1700
rect 12836 1660 12845 1700
rect 12940 1660 13180 1700
rect 13220 1660 13229 1700
rect 13324 1660 13948 1700
rect 13988 1660 13997 1700
rect 14092 1660 14332 1700
rect 14372 1660 14381 1700
rect 14476 1660 14716 1700
rect 14756 1660 14765 1700
rect 15244 1660 15868 1700
rect 15908 1660 15917 1700
rect 16012 1660 16252 1700
rect 16292 1660 16301 1700
rect 18451 1660 18460 1700
rect 18500 1660 19124 1700
rect 19219 1660 19228 1700
rect 19268 1660 20524 1700
rect 20564 1660 20573 1700
rect 12940 1616 12980 1660
rect 13324 1616 13364 1660
rect 14092 1616 14132 1660
rect 67 1576 76 1616
rect 116 1576 7220 1616
rect 8332 1576 11884 1616
rect 11924 1576 11933 1616
rect 12355 1576 12364 1616
rect 12404 1576 12980 1616
rect 13123 1576 13132 1616
rect 13172 1576 13364 1616
rect 13507 1576 13516 1616
rect 13556 1576 14132 1616
rect 7180 1532 7220 1576
rect 14476 1532 14516 1660
rect 15244 1616 15284 1660
rect 15043 1576 15052 1616
rect 15092 1576 15284 1616
rect 16012 1532 16052 1660
rect 19084 1616 19124 1660
rect 19084 1576 21484 1616
rect 21524 1576 21533 1616
rect 4919 1492 4928 1532
rect 4968 1492 5010 1532
rect 5050 1492 5092 1532
rect 5132 1492 5174 1532
rect 5214 1492 5256 1532
rect 5296 1492 5305 1532
rect 7180 1492 13844 1532
rect 13891 1492 13900 1532
rect 13940 1492 14516 1532
rect 15235 1492 15244 1532
rect 15284 1492 16052 1532
rect 16108 1492 19372 1532
rect 19412 1492 19421 1532
rect 20039 1492 20048 1532
rect 20088 1492 20130 1532
rect 20170 1492 20212 1532
rect 20252 1492 20294 1532
rect 20334 1492 20376 1532
rect 20416 1492 20425 1532
rect 0 1448 90 1468
rect 13804 1448 13844 1492
rect 16108 1448 16148 1492
rect 21510 1448 21600 1468
rect 0 1408 76 1448
rect 116 1408 125 1448
rect 13804 1408 16148 1448
rect 21475 1408 21484 1448
rect 21524 1408 21600 1448
rect 0 1388 90 1408
rect 21510 1388 21600 1408
rect 0 1112 90 1132
rect 21510 1112 21600 1132
rect 0 1072 1420 1112
rect 1460 1072 1469 1112
rect 19171 1072 19180 1112
rect 19220 1072 21600 1112
rect 0 1052 90 1072
rect 21510 1052 21600 1072
rect 0 776 90 796
rect 21510 776 21600 796
rect 0 736 15916 776
rect 15956 736 15965 776
rect 20515 736 20524 776
rect 20564 736 21600 776
rect 0 716 90 736
rect 21510 716 21600 736
rect 8803 148 8812 188
rect 8852 148 8861 188
rect 8812 104 8852 148
rect 8812 64 17356 104
rect 17396 64 17405 104
<< via2 >>
rect 1324 11152 1364 11192
rect 19468 11152 19508 11192
rect 8620 10816 8660 10856
rect 19372 10816 19412 10856
rect 4928 10564 4968 10604
rect 5010 10564 5050 10604
rect 5092 10564 5132 10604
rect 5174 10564 5214 10604
rect 5256 10564 5296 10604
rect 20048 10564 20088 10604
rect 20130 10564 20170 10604
rect 20212 10564 20252 10604
rect 20294 10564 20334 10604
rect 20376 10564 20416 10604
rect 172 10480 212 10520
rect 2668 10480 2708 10520
rect 1036 10396 1076 10436
rect 1996 10396 2036 10436
rect 2956 10396 2996 10436
rect 3916 10396 3956 10436
rect 4780 10396 4820 10436
rect 5836 10396 5876 10436
rect 6796 10396 6836 10436
rect 7756 10396 7796 10436
rect 8716 10396 8756 10436
rect 9676 10396 9716 10436
rect 10636 10396 10676 10436
rect 11596 10396 11636 10436
rect 12556 10396 12596 10436
rect 13516 10396 13556 10436
rect 14476 10396 14516 10436
rect 15436 10396 15476 10436
rect 16396 10396 16436 10436
rect 17356 10396 17396 10436
rect 13420 10312 13460 10352
rect 14380 10228 14420 10268
rect 1420 10144 1460 10184
rect 1996 10144 2036 10184
rect 3244 10144 3284 10184
rect 4204 10144 4244 10184
rect 5356 10144 5396 10184
rect 5548 10144 5588 10184
rect 7084 10144 7124 10184
rect 8044 10144 8084 10184
rect 8236 10144 8276 10184
rect 9964 10144 10004 10184
rect 10924 10144 10964 10184
rect 13516 10144 13556 10184
rect 13804 10144 13844 10184
rect 14764 10144 14804 10184
rect 15724 10144 15764 10184
rect 13036 10060 13076 10100
rect 15532 10060 15572 10100
rect 18316 10396 18356 10436
rect 19276 10396 19316 10436
rect 16876 10144 16916 10184
rect 20716 10228 20756 10268
rect 18604 10144 18644 10184
rect 19756 10144 19796 10184
rect 18700 10060 18740 10100
rect 19372 10060 19412 10100
rect 20140 9976 20180 10016
rect 20908 9976 20948 10016
rect 3532 9808 3572 9848
rect 3688 9808 3728 9848
rect 3770 9808 3810 9848
rect 3852 9808 3892 9848
rect 3934 9808 3974 9848
rect 4016 9808 4056 9848
rect 1324 9724 1364 9764
rect 11116 9892 11156 9932
rect 15820 9892 15860 9932
rect 18124 9808 18164 9848
rect 18808 9808 18848 9848
rect 18890 9808 18930 9848
rect 18972 9808 19012 9848
rect 19054 9808 19094 9848
rect 19136 9808 19176 9848
rect 13804 9724 13844 9764
rect 1420 9640 1460 9680
rect 10924 9640 10964 9680
rect 8620 9556 8660 9596
rect 13516 9556 13556 9596
rect 17932 9724 17972 9764
rect 19276 9724 19316 9764
rect 14764 9640 14804 9680
rect 18604 9640 18644 9680
rect 19372 9640 19412 9680
rect 18028 9556 18068 9596
rect 19180 9556 19220 9596
rect 20140 9556 20180 9596
rect 2572 9472 2612 9512
rect 11116 9472 11156 9512
rect 13804 9472 13844 9512
rect 17260 9472 17300 9512
rect 17548 9472 17588 9512
rect 18508 9472 18548 9512
rect 18892 9472 18932 9512
rect 19660 9472 19700 9512
rect 20524 9472 20564 9512
rect 10060 9388 10100 9428
rect 3532 9304 3572 9344
rect 13804 9304 13844 9344
rect 20428 9304 20468 9344
rect 15820 9220 15860 9260
rect 17452 9220 17492 9260
rect 21004 9220 21044 9260
rect 15340 9136 15380 9176
rect 18700 9136 18740 9176
rect 4928 9052 4968 9092
rect 5010 9052 5050 9092
rect 5092 9052 5132 9092
rect 5174 9052 5214 9092
rect 5256 9052 5296 9092
rect 15628 9052 15668 9092
rect 18892 9052 18932 9092
rect 1228 8968 1268 9008
rect 17548 8968 17588 9008
rect 18988 8968 19028 9008
rect 9964 8884 10004 8924
rect 13036 8884 13076 8924
rect 15244 8884 15284 8924
rect 15724 8884 15764 8924
rect 4588 8800 4628 8840
rect 6508 8800 6548 8840
rect 3340 8716 3380 8756
rect 17068 8716 17108 8756
rect 2284 8632 2324 8672
rect 8716 8632 8756 8672
rect 13420 8632 13460 8672
rect 13804 8632 13844 8672
rect 14380 8632 14420 8672
rect 17356 8884 17396 8924
rect 18604 8800 18644 8840
rect 18988 8800 19028 8840
rect 17356 8716 17396 8756
rect 17740 8716 17780 8756
rect 18028 8716 18068 8756
rect 18316 8716 18356 8756
rect 19180 9136 19220 9176
rect 20908 9136 20948 9176
rect 20048 9052 20088 9092
rect 20130 9052 20170 9092
rect 20212 9052 20252 9092
rect 20294 9052 20334 9092
rect 20376 9052 20416 9092
rect 19468 8884 19508 8924
rect 19756 8884 19796 8924
rect 19180 8800 19220 8840
rect 19564 8800 19604 8840
rect 21004 8800 21044 8840
rect 19372 8632 19412 8672
rect 20620 8632 20660 8672
rect 4108 8464 4148 8504
rect 18412 8464 18452 8504
rect 3688 8296 3728 8336
rect 3770 8296 3810 8336
rect 3852 8296 3892 8336
rect 3934 8296 3974 8336
rect 4016 8296 4056 8336
rect 16780 8296 16820 8336
rect 18808 8296 18848 8336
rect 18890 8296 18930 8336
rect 18972 8296 19012 8336
rect 19054 8296 19094 8336
rect 19136 8296 19176 8336
rect 1708 8128 1748 8168
rect 1996 8128 2036 8168
rect 7084 8128 7124 8168
rect 8044 8128 8084 8168
rect 8236 8044 8276 8084
rect 20716 8212 20756 8252
rect 16876 8128 16916 8168
rect 17260 8128 17300 8168
rect 2764 7960 2804 8000
rect 4300 7960 4340 8000
rect 6892 7960 6932 8000
rect 7660 7960 7700 8000
rect 4492 7876 4532 7916
rect 3052 7792 3092 7832
rect 4684 7792 4724 7832
rect 12076 7792 12116 7832
rect 11500 7708 11540 7748
rect 13132 7624 13172 7664
rect 15340 7960 15380 8000
rect 17068 7960 17108 8000
rect 17356 7960 17396 8000
rect 19756 7792 19796 7832
rect 18700 7708 18740 7748
rect 19468 7624 19508 7664
rect 4928 7540 4968 7580
rect 5010 7540 5050 7580
rect 5092 7540 5132 7580
rect 5174 7540 5214 7580
rect 5256 7540 5296 7580
rect 6316 7540 6356 7580
rect 20048 7540 20088 7580
rect 20130 7540 20170 7580
rect 20212 7540 20252 7580
rect 20294 7540 20334 7580
rect 20376 7540 20416 7580
rect 12844 7456 12884 7496
rect 940 7288 980 7328
rect 17356 7288 17396 7328
rect 2956 7120 2996 7160
rect 7660 7204 7700 7244
rect 16972 7204 17012 7244
rect 3628 7120 3668 7160
rect 4876 7120 4916 7160
rect 5548 7120 5588 7160
rect 7756 7120 7796 7160
rect 9004 7120 9044 7160
rect 15244 7120 15284 7160
rect 15532 7120 15572 7160
rect 19852 7120 19892 7160
rect 20524 7120 20564 7160
rect 20812 7120 20852 7160
rect 5452 7036 5492 7076
rect 9196 7036 9236 7076
rect 5740 6952 5780 6992
rect 76 6784 116 6824
rect 9964 6868 10004 6908
rect 3688 6784 3728 6824
rect 3770 6784 3810 6824
rect 3852 6784 3892 6824
rect 3934 6784 3974 6824
rect 4016 6784 4056 6824
rect 4588 6784 4628 6824
rect 18808 6784 18848 6824
rect 18890 6784 18930 6824
rect 18972 6784 19012 6824
rect 19054 6784 19094 6824
rect 19136 6784 19176 6824
rect 19852 6700 19892 6740
rect 3244 6616 3284 6656
rect 10732 6616 10772 6656
rect 9100 6532 9140 6572
rect 10636 6532 10676 6572
rect 18796 6532 18836 6572
rect 20812 6616 20852 6656
rect 76 6448 116 6488
rect 2092 6448 2132 6488
rect 3148 6448 3188 6488
rect 5164 6448 5204 6488
rect 5452 6448 5492 6488
rect 8908 6448 8948 6488
rect 9196 6448 9236 6488
rect 9388 6448 9428 6488
rect 12844 6448 12884 6488
rect 15244 6448 15284 6488
rect 16684 6448 16724 6488
rect 17356 6448 17396 6488
rect 19756 6448 19796 6488
rect 3436 6364 3476 6404
rect 11596 6364 11636 6404
rect 7852 6280 7892 6320
rect 10060 6280 10100 6320
rect 7948 6196 7988 6236
rect 11404 6196 11444 6236
rect 16780 6196 16820 6236
rect 20620 6196 20660 6236
rect 1228 6112 1268 6152
rect 17068 6112 17108 6152
rect 4928 6028 4968 6068
rect 5010 6028 5050 6068
rect 5092 6028 5132 6068
rect 5174 6028 5214 6068
rect 5256 6028 5296 6068
rect 9484 6028 9524 6068
rect 16588 6028 16628 6068
rect 3628 5944 3668 5984
rect 7756 5944 7796 5984
rect 7948 5944 7988 5984
rect 9772 5944 9812 5984
rect 5452 5860 5492 5900
rect 16300 5860 16340 5900
rect 20524 6112 20564 6152
rect 20048 6028 20088 6068
rect 20130 6028 20170 6068
rect 20212 6028 20252 6068
rect 20294 6028 20334 6068
rect 20376 6028 20416 6068
rect 18604 5860 18644 5900
rect 16684 5776 16724 5816
rect 11596 5692 11636 5732
rect 13900 5692 13940 5732
rect 18700 5692 18740 5732
rect 76 5608 116 5648
rect 2188 5608 2228 5648
rect 2668 5608 2708 5648
rect 3340 5608 3380 5648
rect 13708 5608 13748 5648
rect 18508 5608 18548 5648
rect 18892 5608 18932 5648
rect 172 5524 212 5564
rect 4780 5524 4820 5564
rect 9484 5524 9524 5564
rect 76 5440 116 5480
rect 11212 5440 11252 5480
rect 18220 5440 18260 5480
rect 19276 5440 19316 5480
rect 21484 5440 21524 5480
rect 9196 5356 9236 5396
rect 18604 5356 18644 5396
rect 3688 5272 3728 5312
rect 3770 5272 3810 5312
rect 3852 5272 3892 5312
rect 3934 5272 3974 5312
rect 4016 5272 4056 5312
rect 7948 5272 7988 5312
rect 10060 5272 10100 5312
rect 1132 5188 1172 5228
rect 14476 5188 14516 5228
rect 940 5104 980 5144
rect 5452 5104 5492 5144
rect 5356 5020 5396 5060
rect 18808 5272 18848 5312
rect 18890 5272 18930 5312
rect 18972 5272 19012 5312
rect 19054 5272 19094 5312
rect 19136 5272 19176 5312
rect 20620 5020 20660 5060
rect 2380 4936 2420 4976
rect 14380 4936 14420 4976
rect 19084 4936 19124 4976
rect 19852 4936 19892 4976
rect 21484 4936 21524 4976
rect 1420 4852 1460 4892
rect 7948 4768 7988 4808
rect 10924 4768 10964 4808
rect 21292 4768 21332 4808
rect 8236 4684 8276 4724
rect 10540 4684 10580 4724
rect 18796 4684 18836 4724
rect 1324 4600 1364 4640
rect 19084 4600 19124 4640
rect 4928 4516 4968 4556
rect 5010 4516 5050 4556
rect 5092 4516 5132 4556
rect 5174 4516 5214 4556
rect 5256 4516 5296 4556
rect 16780 4516 16820 4556
rect 19852 4516 19892 4556
rect 18508 4432 18548 4472
rect 20048 4516 20088 4556
rect 20130 4516 20170 4556
rect 20212 4516 20252 4556
rect 20294 4516 20334 4556
rect 20376 4516 20416 4556
rect 14668 4348 14708 4388
rect 18220 4348 18260 4388
rect 19852 4348 19892 4388
rect 20140 4348 20180 4388
rect 4204 4264 4244 4304
rect 6508 4264 6548 4304
rect 7372 4264 7412 4304
rect 21292 4264 21332 4304
rect 10156 4180 10196 4220
rect 12940 4180 12980 4220
rect 20524 4180 20564 4220
rect 1420 4096 1460 4136
rect 2764 4096 2804 4136
rect 4108 4096 4148 4136
rect 7756 4096 7796 4136
rect 11980 4096 12020 4136
rect 12172 4096 12212 4136
rect 14284 4096 14324 4136
rect 16492 4096 16532 4136
rect 16684 4096 16724 4136
rect 18796 4096 18836 4136
rect 20428 4096 20468 4136
rect 5836 4012 5876 4052
rect 7564 4012 7604 4052
rect 13996 4012 14036 4052
rect 10348 3928 10388 3968
rect 13036 3928 13076 3968
rect 13228 3928 13268 3968
rect 13804 3928 13844 3968
rect 14188 3928 14228 3968
rect 8620 3844 8660 3884
rect 13612 3844 13652 3884
rect 15820 3928 15860 3968
rect 17356 3928 17396 3968
rect 18220 3928 18260 3968
rect 3688 3760 3728 3800
rect 3770 3760 3810 3800
rect 3852 3760 3892 3800
rect 3934 3760 3974 3800
rect 4016 3760 4056 3800
rect 8524 3760 8564 3800
rect 18808 3760 18848 3800
rect 18890 3760 18930 3800
rect 18972 3760 19012 3800
rect 19054 3760 19094 3800
rect 19136 3760 19176 3800
rect 14380 3676 14420 3716
rect 13708 3592 13748 3632
rect 20428 3592 20468 3632
rect 6316 3508 6356 3548
rect 7948 3508 7988 3548
rect 11980 3508 12020 3548
rect 2476 3424 2516 3464
rect 3052 3424 3092 3464
rect 17068 3424 17108 3464
rect 19276 3424 19316 3464
rect 20140 3424 20180 3464
rect 5644 3340 5684 3380
rect 6220 3340 6260 3380
rect 10060 3340 10100 3380
rect 18604 3340 18644 3380
rect 6988 3256 7028 3296
rect 21004 3256 21044 3296
rect 7180 3172 7220 3212
rect 8140 3172 8180 3212
rect 12172 3172 12212 3212
rect 14380 3172 14420 3212
rect 15916 3172 15956 3212
rect 17452 3172 17492 3212
rect 13900 3088 13940 3128
rect 4928 3004 4968 3044
rect 5010 3004 5050 3044
rect 5092 3004 5132 3044
rect 5174 3004 5214 3044
rect 5256 3004 5296 3044
rect 6028 3004 6068 3044
rect 8428 3004 8468 3044
rect 14284 3004 14324 3044
rect 20048 3004 20088 3044
rect 20130 3004 20170 3044
rect 20212 3004 20252 3044
rect 20294 3004 20334 3044
rect 20376 3004 20416 3044
rect 7180 2920 7220 2960
rect 16684 2920 16724 2960
rect 18604 2836 18644 2876
rect 1132 2752 1172 2792
rect 9100 2752 9140 2792
rect 2284 2668 2324 2708
rect 9484 2668 9524 2708
rect 17260 2752 17300 2792
rect 21004 2752 21044 2792
rect 14188 2668 14228 2708
rect 15916 2668 15956 2708
rect 19948 2668 19988 2708
rect 1804 2584 1844 2624
rect 8812 2584 8852 2624
rect 9196 2584 9236 2624
rect 9580 2584 9620 2624
rect 9964 2584 10004 2624
rect 10732 2584 10772 2624
rect 13228 2584 13268 2624
rect 13612 2584 13652 2624
rect 13996 2584 14036 2624
rect 14380 2584 14420 2624
rect 15436 2584 15476 2624
rect 16012 2584 16052 2624
rect 16780 2584 16820 2624
rect 18892 2584 18932 2624
rect 19372 2584 19412 2624
rect 1996 2500 2036 2540
rect 7660 2500 7700 2540
rect 11692 2500 11732 2540
rect 11884 2500 11924 2540
rect 15628 2500 15668 2540
rect 1324 2416 1364 2456
rect 8044 2416 8084 2456
rect 8908 2416 8948 2456
rect 9292 2416 9332 2456
rect 9676 2416 9716 2456
rect 10060 2416 10100 2456
rect 10444 2416 10484 2456
rect 10828 2416 10868 2456
rect 12556 2416 12596 2456
rect 13036 2416 13076 2456
rect 13324 2416 13364 2456
rect 13708 2416 13748 2456
rect 14092 2416 14132 2456
rect 14476 2416 14516 2456
rect 14860 2416 14900 2456
rect 15724 2416 15764 2456
rect 15916 2416 15956 2456
rect 1420 2332 1460 2372
rect 8332 2332 8372 2372
rect 11980 2332 12020 2372
rect 12172 2332 12212 2372
rect 14572 2332 14612 2372
rect 15340 2332 15380 2372
rect 3688 2248 3728 2288
rect 3770 2248 3810 2288
rect 3852 2248 3892 2288
rect 3934 2248 3974 2288
rect 4016 2248 4056 2288
rect 6796 2248 6836 2288
rect 15436 2248 15476 2288
rect 6604 2164 6644 2204
rect 9100 2164 9140 2204
rect 7660 2080 7700 2120
rect 8812 2080 8852 2120
rect 14380 2080 14420 2120
rect 15340 2080 15380 2120
rect 17260 2080 17300 2120
rect 7852 1996 7892 2036
rect 11500 1996 11540 2036
rect 13516 1996 13556 2036
rect 15724 1996 15764 2036
rect 17356 1996 17396 2036
rect 18220 1996 18260 2036
rect 8236 1912 8276 1952
rect 8428 1912 8468 1952
rect 9004 1912 9044 1952
rect 9772 1912 9812 1952
rect 10540 1912 10580 1952
rect 10924 1912 10964 1952
rect 11212 1912 11252 1952
rect 11404 1912 11444 1952
rect 12076 1912 12116 1952
rect 13132 1912 13172 1952
rect 13804 1912 13844 1952
rect 14668 1912 14708 1952
rect 15628 1912 15668 1952
rect 17452 1912 17492 1952
rect 18808 2248 18848 2288
rect 18890 2248 18930 2288
rect 18972 2248 19012 2288
rect 19054 2248 19094 2288
rect 19136 2248 19176 2288
rect 18604 1996 18644 2036
rect 6412 1828 6452 1868
rect 8620 1828 8660 1868
rect 12172 1828 12212 1868
rect 15820 1828 15860 1868
rect 20428 2416 20468 2456
rect 20428 1996 20468 2036
rect 20620 1912 20660 1952
rect 11404 1744 11444 1784
rect 11788 1744 11828 1784
rect 12748 1744 12788 1784
rect 14668 1744 14708 1784
rect 15628 1744 15668 1784
rect 19180 1744 19220 1784
rect 8716 1660 8756 1700
rect 9100 1660 9140 1700
rect 9484 1660 9524 1700
rect 9868 1660 9908 1700
rect 10252 1660 10292 1700
rect 10636 1660 10676 1700
rect 11020 1660 11060 1700
rect 11212 1660 11252 1700
rect 11596 1660 11636 1700
rect 11980 1660 12020 1700
rect 12172 1660 12212 1700
rect 20524 1660 20564 1700
rect 76 1576 116 1616
rect 11884 1576 11924 1616
rect 12364 1576 12404 1616
rect 13132 1576 13172 1616
rect 13516 1576 13556 1616
rect 15052 1576 15092 1616
rect 21484 1576 21524 1616
rect 4928 1492 4968 1532
rect 5010 1492 5050 1532
rect 5092 1492 5132 1532
rect 5174 1492 5214 1532
rect 5256 1492 5296 1532
rect 13900 1492 13940 1532
rect 15244 1492 15284 1532
rect 19372 1492 19412 1532
rect 20048 1492 20088 1532
rect 20130 1492 20170 1532
rect 20212 1492 20252 1532
rect 20294 1492 20334 1532
rect 20376 1492 20416 1532
rect 76 1408 116 1448
rect 21484 1408 21524 1448
rect 1420 1072 1460 1112
rect 19180 1072 19220 1112
rect 15916 736 15956 776
rect 20524 736 20564 776
rect 8812 148 8852 188
rect 17356 64 17396 104
<< metal3 >>
rect 1016 12100 1096 12180
rect 1976 12100 2056 12180
rect 2936 12100 3016 12180
rect 3896 12100 3976 12180
rect 4856 12100 4936 12180
rect 5816 12100 5896 12180
rect 6776 12100 6856 12180
rect 7736 12100 7816 12180
rect 8696 12100 8776 12180
rect 9656 12100 9736 12180
rect 10616 12100 10696 12180
rect 11576 12100 11656 12180
rect 12536 12100 12616 12180
rect 13496 12100 13576 12180
rect 14456 12100 14536 12180
rect 15416 12100 15496 12180
rect 16376 12100 16456 12180
rect 17336 12100 17416 12180
rect 18296 12100 18376 12180
rect 19256 12100 19336 12180
rect 20216 12100 20296 12180
rect 172 10520 212 10529
rect 76 6824 116 6835
rect 76 6740 116 6784
rect 76 6691 116 6700
rect 76 6572 116 6581
rect 76 6488 116 6532
rect 76 6437 116 6448
rect 76 5648 116 5657
rect 76 5480 116 5608
rect 172 5564 212 10480
rect 1036 10436 1076 12100
rect 1036 10387 1076 10396
rect 1324 11192 1364 11201
rect 1324 9764 1364 11152
rect 1996 10436 2036 12100
rect 1996 10387 2036 10396
rect 2668 10520 2708 10529
rect 1324 9715 1364 9724
rect 1420 10184 1460 10193
rect 1420 9680 1460 10144
rect 1420 9631 1460 9640
rect 1996 10184 2036 10193
rect 1228 9008 1268 9017
rect 172 5515 212 5524
rect 940 7328 980 7337
rect 76 5431 116 5440
rect 940 5144 980 7288
rect 1228 6152 1268 8968
rect 1708 8168 1748 8177
rect 1708 6488 1748 8128
rect 1996 8168 2036 10144
rect 2572 9512 2612 9521
rect 1996 8119 2036 8128
rect 2284 8672 2324 8681
rect 1708 6439 1748 6448
rect 2092 6488 2132 6497
rect 1228 6103 1268 6112
rect 940 5095 980 5104
rect 1132 5228 1172 5237
rect 1132 2792 1172 5188
rect 1420 4892 1460 4901
rect 1132 2743 1172 2752
rect 1324 4640 1364 4649
rect 1324 2456 1364 4600
rect 1420 4136 1460 4852
rect 1420 4087 1460 4096
rect 1324 2407 1364 2416
rect 1804 2624 1844 2633
rect 1420 2372 1460 2381
rect 76 1616 116 1625
rect 76 1448 116 1576
rect 76 1399 116 1408
rect 1420 1112 1460 2332
rect 1420 1063 1460 1072
rect 1804 80 1844 2584
rect 1996 2540 2036 2549
rect 1996 80 2036 2500
rect 2092 272 2132 6448
rect 2092 223 2132 232
rect 2188 5648 2228 5657
rect 2188 80 2228 5608
rect 2284 2708 2324 8632
rect 2284 2659 2324 2668
rect 2380 4976 2420 4985
rect 2380 80 2420 4936
rect 2476 3464 2516 3473
rect 2476 188 2516 3424
rect 2572 356 2612 9472
rect 2668 5648 2708 10480
rect 2956 10436 2996 12100
rect 2956 10387 2996 10396
rect 3916 10436 3956 12100
rect 4876 11108 4916 12100
rect 3916 10387 3956 10396
rect 4780 11068 4916 11108
rect 4780 10436 4820 11068
rect 4928 10604 5296 10613
rect 4968 10564 5010 10604
rect 5050 10564 5092 10604
rect 5132 10564 5174 10604
rect 5214 10564 5256 10604
rect 4928 10555 5296 10564
rect 4780 10387 4820 10396
rect 5836 10436 5876 12100
rect 5836 10387 5876 10396
rect 6796 10436 6836 12100
rect 6796 10387 6836 10396
rect 7756 10436 7796 12100
rect 7756 10387 7796 10396
rect 8620 10856 8660 10865
rect 3244 10184 3284 10193
rect 2668 5599 2708 5608
rect 2764 8000 2804 8009
rect 2764 4304 2804 7960
rect 3052 7832 3092 7841
rect 2668 4264 2804 4304
rect 2956 7160 2996 7169
rect 2668 524 2708 4264
rect 2668 475 2708 484
rect 2764 4136 2804 4145
rect 2572 316 2708 356
rect 2668 188 2708 316
rect 2476 148 2612 188
rect 2572 80 2612 148
rect 2668 139 2708 148
rect 2764 80 2804 4096
rect 2956 80 2996 7120
rect 3052 3464 3092 7792
rect 3244 6656 3284 10144
rect 4204 10184 4244 10193
rect 3532 9848 3572 9857
rect 3532 9344 3572 9808
rect 3688 9848 4056 9857
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 3688 9799 4056 9808
rect 3532 9295 3572 9304
rect 3244 6607 3284 6616
rect 3340 8756 3380 8765
rect 3052 3415 3092 3424
rect 3148 6488 3188 6497
rect 3340 6488 3380 8716
rect 4108 8504 4148 8513
rect 3688 8336 4056 8345
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 3688 8287 4056 8296
rect 3628 7160 3668 7169
rect 3148 80 3188 6448
rect 3244 6448 3380 6488
rect 3532 7120 3628 7160
rect 3244 3968 3284 6448
rect 3436 6404 3476 6413
rect 3244 3919 3284 3928
rect 3340 5648 3380 5657
rect 3244 3800 3284 3809
rect 3244 2120 3284 3760
rect 3244 2071 3284 2080
rect 3340 80 3380 5608
rect 3436 2036 3476 6364
rect 3532 2120 3572 7120
rect 3628 7111 3668 7120
rect 3688 6824 4056 6833
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 3688 6775 4056 6784
rect 3628 5984 3668 5993
rect 3628 5480 3668 5944
rect 3628 5431 3668 5440
rect 3688 5312 4056 5321
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 3688 5263 4056 5272
rect 4108 4136 4148 8464
rect 4204 4304 4244 10144
rect 5356 10184 5396 10193
rect 4928 9092 5296 9101
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 4928 9043 5296 9052
rect 4588 8840 4628 8849
rect 4204 4255 4244 4264
rect 4300 8000 4340 8009
rect 4108 4087 4148 4096
rect 4108 3968 4148 3977
rect 3688 3800 4056 3809
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 3688 3751 4056 3760
rect 3688 2288 4056 2297
rect 3728 2248 3770 2288
rect 3810 2248 3852 2288
rect 3892 2248 3934 2288
rect 3974 2248 4016 2288
rect 3688 2239 4056 2248
rect 3916 2120 3956 2129
rect 3532 2080 3764 2120
rect 3436 1996 3572 2036
rect 3532 80 3572 1996
rect 3724 80 3764 2080
rect 3916 80 3956 2080
rect 4108 80 4148 3928
rect 4300 80 4340 7960
rect 4492 7916 4532 7925
rect 4492 80 4532 7876
rect 4588 6824 4628 8800
rect 4588 6775 4628 6784
rect 4684 7832 4724 7841
rect 4684 80 4724 7792
rect 4928 7580 5296 7589
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 4928 7531 5296 7540
rect 4876 7160 4916 7169
rect 4876 7025 4916 7120
rect 5356 6740 5396 10144
rect 5548 10184 5588 10193
rect 5548 7160 5588 10144
rect 7084 10184 7124 10193
rect 6508 8840 6548 8849
rect 5548 7111 5588 7120
rect 6316 7580 6356 7589
rect 5452 7076 5492 7085
rect 5452 6992 5492 7036
rect 5740 6992 5780 7001
rect 5452 6952 5740 6992
rect 5740 6943 5780 6952
rect 5164 6700 5396 6740
rect 5164 6488 5204 6700
rect 5164 6439 5204 6448
rect 5452 6488 5492 6497
rect 4928 6068 5296 6077
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 4928 6019 5296 6028
rect 5452 5900 5492 6448
rect 5452 5851 5492 5860
rect 4780 5564 4820 5573
rect 4780 1364 4820 5524
rect 5452 5144 5492 5153
rect 5356 5060 5396 5069
rect 4928 4556 5296 4565
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 4928 4507 5296 4516
rect 4928 3044 5296 3053
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 4928 2995 5296 3004
rect 4928 1532 5296 1541
rect 4968 1492 5010 1532
rect 5050 1492 5092 1532
rect 5132 1492 5174 1532
rect 5214 1492 5256 1532
rect 4928 1483 5296 1492
rect 5356 1364 5396 5020
rect 4780 1324 5108 1364
rect 4876 1196 4916 1205
rect 4876 80 4916 1156
rect 5068 80 5108 1324
rect 5260 1324 5396 1364
rect 5260 80 5300 1324
rect 5452 80 5492 5104
rect 5836 4052 5876 4061
rect 5644 3380 5684 3389
rect 5644 80 5684 3340
rect 5836 80 5876 4012
rect 6316 3548 6356 7540
rect 6508 4304 6548 8800
rect 7084 8168 7124 10144
rect 7084 8119 7124 8128
rect 8044 10184 8084 10193
rect 8044 8168 8084 10144
rect 8044 8119 8084 8128
rect 8236 10184 8276 10193
rect 8236 8084 8276 10144
rect 8620 9596 8660 10816
rect 8716 10436 8756 12100
rect 8716 10387 8756 10396
rect 9676 10436 9716 12100
rect 9676 10387 9716 10396
rect 10636 10436 10676 12100
rect 10636 10387 10676 10396
rect 11596 10436 11636 12100
rect 11596 10387 11636 10396
rect 12556 10436 12596 12100
rect 12556 10387 12596 10396
rect 13516 10436 13556 12100
rect 13516 10387 13556 10396
rect 14476 10436 14516 12100
rect 14476 10387 14516 10396
rect 15436 10436 15476 12100
rect 15436 10387 15476 10396
rect 16396 10436 16436 12100
rect 16396 10387 16436 10396
rect 17356 10436 17396 12100
rect 17356 10387 17396 10396
rect 18316 10436 18356 12100
rect 18316 10387 18356 10396
rect 19276 10436 19316 12100
rect 19468 11192 19508 11201
rect 19276 10387 19316 10396
rect 19372 10856 19412 10865
rect 13420 10352 13460 10361
rect 8620 9547 8660 9556
rect 9964 10184 10004 10193
rect 9964 8924 10004 10144
rect 10924 10184 10964 10193
rect 10924 9680 10964 10144
rect 13036 10100 13076 10109
rect 10924 9631 10964 9640
rect 11116 9932 11156 9941
rect 11116 9512 11156 9892
rect 11116 9463 11156 9472
rect 10060 9428 10100 9437
rect 10060 9293 10100 9388
rect 9964 8875 10004 8884
rect 13036 8924 13076 10060
rect 13036 8875 13076 8884
rect 8236 8035 8276 8044
rect 8716 8672 8756 8681
rect 6508 4255 6548 4264
rect 6892 8000 6932 8009
rect 6316 3499 6356 3508
rect 6220 3380 6260 3389
rect 6028 3044 6068 3053
rect 6028 80 6068 3004
rect 6220 80 6260 3340
rect 6796 2288 6836 2297
rect 6604 2204 6644 2213
rect 6412 1868 6452 1877
rect 6412 80 6452 1828
rect 6604 80 6644 2164
rect 6796 80 6836 2248
rect 6892 356 6932 7960
rect 7660 8000 7700 8009
rect 7660 7244 7700 7960
rect 7660 7195 7700 7204
rect 7756 7160 7796 7169
rect 7756 5984 7796 7120
rect 7756 5935 7796 5944
rect 7852 6320 7892 6329
rect 7372 4304 7412 4313
rect 6892 307 6932 316
rect 6988 3296 7028 3305
rect 6988 80 7028 3256
rect 7180 3212 7220 3221
rect 7180 2960 7220 3172
rect 7180 2911 7220 2920
rect 7180 440 7220 449
rect 7180 80 7220 400
rect 7372 80 7412 4264
rect 7756 4136 7796 4145
rect 7564 4052 7604 4061
rect 7564 80 7604 4012
rect 7660 2540 7700 2549
rect 7660 2120 7700 2500
rect 7660 2071 7700 2080
rect 7756 80 7796 4096
rect 7852 2036 7892 6280
rect 7948 6236 7988 6245
rect 7948 5984 7988 6196
rect 7948 5935 7988 5944
rect 7948 5312 7988 5321
rect 7948 4808 7988 5272
rect 7948 4759 7988 4768
rect 8236 4724 8276 4733
rect 7852 1987 7892 1996
rect 7948 3548 7988 3557
rect 7948 80 7988 3508
rect 8140 3212 8180 3221
rect 8044 2456 8084 2465
rect 8044 1952 8084 2416
rect 8044 1903 8084 1912
rect 8140 80 8180 3172
rect 8236 1952 8276 4684
rect 8620 3884 8660 3893
rect 8524 3800 8564 3809
rect 8428 3044 8468 3053
rect 8332 2372 8372 2381
rect 8332 2237 8372 2332
rect 8428 2120 8468 3004
rect 8236 1903 8276 1912
rect 8332 2080 8468 2120
rect 8332 80 8372 2080
rect 8428 1952 8468 1961
rect 8428 1817 8468 1912
rect 8524 80 8564 3760
rect 8620 1868 8660 3844
rect 8716 1952 8756 8632
rect 13420 8672 13460 10312
rect 14380 10268 14420 10277
rect 19372 10268 19412 10816
rect 13516 10184 13556 10193
rect 13516 9596 13556 10144
rect 13804 10184 13844 10193
rect 13804 9764 13844 10144
rect 13804 9715 13844 9724
rect 13516 9547 13556 9556
rect 13804 9512 13844 9607
rect 13804 9463 13844 9472
rect 13420 8623 13460 8632
rect 13804 9344 13844 9353
rect 13804 8672 13844 9304
rect 13804 8623 13844 8632
rect 14380 8672 14420 10228
rect 19276 10228 19412 10268
rect 14764 10184 14804 10193
rect 14764 9680 14804 10144
rect 15724 10184 15764 10193
rect 14764 9631 14804 9640
rect 15532 10100 15572 10109
rect 15340 9176 15380 9185
rect 15244 8924 15284 8933
rect 15244 8789 15284 8884
rect 14380 8623 14420 8632
rect 15340 8000 15380 9136
rect 15340 7951 15380 7960
rect 12076 7832 12116 7841
rect 11500 7748 11540 7757
rect 9004 7160 9044 7169
rect 8908 6740 8948 6749
rect 8908 6488 8948 6700
rect 8908 6439 8948 6448
rect 8812 2624 8852 2633
rect 8812 2120 8852 2584
rect 8812 2071 8852 2080
rect 8908 2456 8948 2465
rect 8716 1912 8852 1952
rect 8620 1819 8660 1828
rect 8716 1700 8756 1709
rect 8716 80 8756 1660
rect 8812 188 8852 1912
rect 8812 139 8852 148
rect 8908 80 8948 2416
rect 9004 1952 9044 7120
rect 9484 7160 9524 7169
rect 9196 7076 9236 7085
rect 9100 6572 9140 6581
rect 9100 6437 9140 6532
rect 9196 6488 9236 7036
rect 9196 6439 9236 6448
rect 9388 6488 9428 6497
rect 9196 5396 9236 5405
rect 9100 2792 9140 2801
rect 9100 2624 9140 2752
rect 9100 2575 9140 2584
rect 9196 2624 9236 5356
rect 9196 2575 9236 2584
rect 9292 2456 9332 2465
rect 9100 2372 9140 2381
rect 9100 2204 9140 2332
rect 9100 2155 9140 2164
rect 9004 1903 9044 1912
rect 9100 1700 9140 1709
rect 9100 80 9140 1660
rect 9292 80 9332 2416
rect 9388 1196 9428 6448
rect 9484 6068 9524 7120
rect 9484 6019 9524 6028
rect 9964 6908 10004 6917
rect 9772 5984 9812 5993
rect 9484 5564 9524 5573
rect 9484 2708 9524 5524
rect 9484 2659 9524 2668
rect 9580 2624 9620 2633
rect 9580 2489 9620 2584
rect 9676 2456 9716 2465
rect 9388 1147 9428 1156
rect 9484 1700 9524 1709
rect 9484 80 9524 1660
rect 9676 80 9716 2416
rect 9772 1952 9812 5944
rect 9964 2624 10004 6868
rect 10732 6656 10772 6665
rect 10636 6572 10676 6581
rect 10636 6437 10676 6532
rect 10060 6320 10100 6329
rect 10060 5312 10100 6280
rect 10060 5263 10100 5272
rect 10540 4724 10580 4733
rect 10156 4220 10196 4229
rect 10060 3380 10100 3389
rect 10060 3245 10100 3340
rect 9964 2575 10004 2584
rect 9772 1903 9812 1912
rect 10060 2456 10100 2465
rect 9868 1700 9908 1709
rect 9868 80 9908 1660
rect 10060 80 10100 2416
rect 10156 1280 10196 4180
rect 10348 4220 10388 4229
rect 10348 3968 10388 4180
rect 10348 3919 10388 3928
rect 10444 2456 10484 2465
rect 10156 1231 10196 1240
rect 10252 1700 10292 1709
rect 10252 80 10292 1660
rect 10444 80 10484 2416
rect 10540 1952 10580 4684
rect 10732 2624 10772 6616
rect 11404 6236 11444 6245
rect 11212 5480 11252 5489
rect 10732 2575 10772 2584
rect 10924 4808 10964 4817
rect 10540 1903 10580 1912
rect 10828 2456 10868 2465
rect 10636 1700 10676 1709
rect 10636 80 10676 1660
rect 10828 80 10868 2416
rect 10924 1952 10964 4768
rect 10924 1903 10964 1912
rect 11212 1952 11252 5440
rect 11212 1903 11252 1912
rect 11404 1952 11444 6196
rect 11500 2036 11540 7708
rect 11596 6404 11636 6413
rect 11596 5732 11636 6364
rect 11596 5683 11636 5692
rect 11980 4136 12020 4145
rect 11980 3548 12020 4096
rect 11980 3499 12020 3508
rect 11692 2540 11732 2549
rect 11692 2405 11732 2500
rect 11884 2540 11924 2549
rect 11500 1987 11540 1996
rect 11404 1903 11444 1912
rect 11404 1784 11444 1793
rect 11020 1700 11060 1709
rect 11020 80 11060 1660
rect 11212 1700 11252 1709
rect 11212 80 11252 1660
rect 11404 80 11444 1744
rect 11788 1784 11828 1793
rect 11596 1700 11636 1709
rect 11596 80 11636 1660
rect 11788 80 11828 1744
rect 11884 1616 11924 2500
rect 11980 2456 12020 2465
rect 11980 2372 12020 2416
rect 11980 2321 12020 2332
rect 12076 1952 12116 7792
rect 13132 7664 13172 7673
rect 12844 7496 12884 7505
rect 12844 6488 12884 7456
rect 12844 6439 12884 6448
rect 12940 4220 12980 4229
rect 12172 4136 12212 4145
rect 12172 3212 12212 4096
rect 12940 4085 12980 4180
rect 12172 3163 12212 3172
rect 13036 3968 13076 3977
rect 13036 2624 13076 3928
rect 13036 2575 13076 2584
rect 12556 2456 12596 2465
rect 12076 1903 12116 1912
rect 12172 2372 12212 2381
rect 12172 1868 12212 2332
rect 12172 1819 12212 1828
rect 11884 1567 11924 1576
rect 11980 1700 12020 1709
rect 11980 80 12020 1660
rect 12172 1700 12212 1709
rect 12172 80 12212 1660
rect 12364 1616 12404 1625
rect 12364 80 12404 1576
rect 12556 80 12596 2416
rect 13036 2456 13076 2465
rect 12748 1784 12788 1793
rect 12748 80 12788 1744
rect 13036 440 13076 2416
rect 13132 1952 13172 7624
rect 15244 7160 15284 7169
rect 15244 6488 15284 7120
rect 15532 7160 15572 10060
rect 15628 9092 15668 9101
rect 15628 8924 15668 9052
rect 15628 8875 15668 8884
rect 15724 8924 15764 10144
rect 16876 10184 16916 10193
rect 15820 9932 15860 9941
rect 15820 9260 15860 9892
rect 15820 9211 15860 9220
rect 15724 8875 15764 8884
rect 16780 8336 16820 8345
rect 16780 8000 16820 8296
rect 16876 8168 16916 10144
rect 18604 10184 18644 10193
rect 18124 9848 18164 9857
rect 17932 9764 17972 9773
rect 17260 9512 17300 9521
rect 17260 8924 17300 9472
rect 17548 9512 17588 9521
rect 17452 9260 17492 9269
rect 17356 8924 17396 8933
rect 17260 8884 17356 8924
rect 17356 8875 17396 8884
rect 17452 8840 17492 9220
rect 17548 9008 17588 9472
rect 17548 8959 17588 8968
rect 17452 8800 17588 8840
rect 17068 8756 17108 8765
rect 17356 8756 17396 8765
rect 17108 8716 17356 8756
rect 17068 8707 17108 8716
rect 17356 8707 17396 8716
rect 16876 8119 16916 8128
rect 17260 8168 17300 8177
rect 17068 8000 17108 8009
rect 16780 7960 16916 8000
rect 15532 7111 15572 7120
rect 15244 6439 15284 6448
rect 16684 6488 16724 6497
rect 16588 6068 16628 6077
rect 16300 5900 16340 5909
rect 13900 5732 13940 5741
rect 13708 5648 13748 5657
rect 13228 3968 13268 3977
rect 13228 2624 13268 3928
rect 13612 3884 13652 3893
rect 13228 2575 13268 2584
rect 13516 2624 13556 2633
rect 13132 1903 13172 1912
rect 13324 2456 13364 2465
rect 12940 400 13076 440
rect 13132 1616 13172 1625
rect 12940 80 12980 400
rect 13132 80 13172 1576
rect 13324 80 13364 2416
rect 13516 2036 13556 2584
rect 13612 2624 13652 3844
rect 13708 3632 13748 5608
rect 13708 3583 13748 3592
rect 13804 3968 13844 3977
rect 13612 2575 13652 2584
rect 13516 1987 13556 1996
rect 13708 2456 13748 2465
rect 13516 1616 13556 1625
rect 13516 80 13556 1576
rect 13708 80 13748 2416
rect 13804 1952 13844 3928
rect 13900 3128 13940 5692
rect 14476 5648 14516 5657
rect 14476 5228 14516 5608
rect 14476 5179 14516 5188
rect 14380 4976 14420 4985
rect 14284 4136 14324 4145
rect 13900 3079 13940 3088
rect 13996 4052 14036 4061
rect 13996 2624 14036 4012
rect 14188 3968 14228 3977
rect 14188 2708 14228 3928
rect 14284 3044 14324 4096
rect 14380 3716 14420 4936
rect 14380 3667 14420 3676
rect 14668 4388 14708 4397
rect 14284 2995 14324 3004
rect 14380 3212 14420 3221
rect 14188 2659 14228 2668
rect 13996 2575 14036 2584
rect 14380 2624 14420 3172
rect 14380 2575 14420 2584
rect 13804 1903 13844 1912
rect 14092 2456 14132 2465
rect 13900 1532 13940 1541
rect 13900 80 13940 1492
rect 14092 80 14132 2416
rect 14476 2456 14516 2465
rect 14380 2120 14420 2129
rect 14380 860 14420 2080
rect 14284 820 14420 860
rect 14284 80 14324 820
rect 14476 80 14516 2416
rect 14572 2372 14612 2381
rect 14572 2237 14612 2332
rect 14668 1952 14708 4348
rect 15820 3968 15860 3977
rect 15436 2624 15476 2633
rect 14668 1903 14708 1912
rect 14860 2456 14900 2465
rect 14668 1784 14708 1793
rect 14668 80 14708 1744
rect 14860 80 14900 2416
rect 15340 2372 15380 2381
rect 15340 2120 15380 2332
rect 15436 2288 15476 2584
rect 15436 2239 15476 2248
rect 15628 2540 15668 2549
rect 15340 2071 15380 2080
rect 15628 1952 15668 2500
rect 15724 2456 15764 2465
rect 15724 2036 15764 2416
rect 15724 1987 15764 1996
rect 15628 1903 15668 1912
rect 15820 1868 15860 3928
rect 15916 3212 15956 3221
rect 15916 2708 15956 3172
rect 15916 2659 15956 2668
rect 16012 2624 16052 2633
rect 15820 1819 15860 1828
rect 15916 2456 15956 2465
rect 15628 1784 15668 1793
rect 15436 1744 15628 1784
rect 15052 1616 15092 1625
rect 15052 80 15092 1576
rect 15244 1532 15284 1541
rect 15244 80 15284 1492
rect 15436 80 15476 1744
rect 15628 1735 15668 1744
rect 15916 776 15956 2416
rect 16012 2372 16052 2584
rect 16012 2323 16052 2332
rect 15916 727 15956 736
rect 16204 1280 16244 1289
rect 15820 524 15860 533
rect 15628 188 15668 197
rect 15628 80 15668 148
rect 15820 80 15860 484
rect 16012 272 16052 281
rect 16012 80 16052 232
rect 16204 80 16244 1240
rect 16300 1028 16340 5860
rect 16492 4136 16532 4145
rect 16300 988 16436 1028
rect 16396 80 16436 988
rect 16492 440 16532 4096
rect 16492 391 16532 400
rect 16588 80 16628 6028
rect 16684 5816 16724 6448
rect 16684 5767 16724 5776
rect 16780 6236 16820 6245
rect 16780 4556 16820 6196
rect 16780 4507 16820 4516
rect 16684 4136 16724 4145
rect 16684 2960 16724 4096
rect 16684 2911 16724 2920
rect 16876 2900 16916 7960
rect 16972 7244 17012 7253
rect 16972 5984 17012 7204
rect 17068 6572 17108 7960
rect 17068 6523 17108 6532
rect 17068 6152 17108 6161
rect 17260 6152 17300 8128
rect 17356 8000 17396 8009
rect 17356 7328 17396 7960
rect 17356 7279 17396 7288
rect 17356 6488 17396 6497
rect 17356 6353 17396 6448
rect 17108 6112 17300 6152
rect 17068 6103 17108 6112
rect 16972 5944 17204 5984
rect 17068 3464 17108 3473
rect 17068 3380 17108 3424
rect 17068 3329 17108 3340
rect 16876 2860 17012 2900
rect 16780 2624 16820 2633
rect 16780 2456 16820 2584
rect 16780 2407 16820 2416
rect 16780 356 16820 365
rect 16780 80 16820 316
rect 16972 80 17012 2860
rect 17164 80 17204 5944
rect 17356 3968 17396 3977
rect 17260 2792 17300 2801
rect 17260 2120 17300 2752
rect 17260 2071 17300 2080
rect 17356 2036 17396 3928
rect 17356 1987 17396 1996
rect 17452 3212 17492 3221
rect 17452 1952 17492 3172
rect 17452 1903 17492 1912
rect 17356 104 17396 113
rect 1784 0 1864 80
rect 1976 0 2056 80
rect 2168 0 2248 80
rect 2360 0 2440 80
rect 2552 0 2632 80
rect 2744 0 2824 80
rect 2936 0 3016 80
rect 3128 0 3208 80
rect 3320 0 3400 80
rect 3512 0 3592 80
rect 3704 0 3784 80
rect 3896 0 3976 80
rect 4088 0 4168 80
rect 4280 0 4360 80
rect 4472 0 4552 80
rect 4664 0 4744 80
rect 4856 0 4936 80
rect 5048 0 5128 80
rect 5240 0 5320 80
rect 5432 0 5512 80
rect 5624 0 5704 80
rect 5816 0 5896 80
rect 6008 0 6088 80
rect 6200 0 6280 80
rect 6392 0 6472 80
rect 6584 0 6664 80
rect 6776 0 6856 80
rect 6968 0 7048 80
rect 7160 0 7240 80
rect 7352 0 7432 80
rect 7544 0 7624 80
rect 7736 0 7816 80
rect 7928 0 8008 80
rect 8120 0 8200 80
rect 8312 0 8392 80
rect 8504 0 8584 80
rect 8696 0 8776 80
rect 8888 0 8968 80
rect 9080 0 9160 80
rect 9272 0 9352 80
rect 9464 0 9544 80
rect 9656 0 9736 80
rect 9848 0 9928 80
rect 10040 0 10120 80
rect 10232 0 10312 80
rect 10424 0 10504 80
rect 10616 0 10696 80
rect 10808 0 10888 80
rect 11000 0 11080 80
rect 11192 0 11272 80
rect 11384 0 11464 80
rect 11576 0 11656 80
rect 11768 0 11848 80
rect 11960 0 12040 80
rect 12152 0 12232 80
rect 12344 0 12424 80
rect 12536 0 12616 80
rect 12728 0 12808 80
rect 12920 0 13000 80
rect 13112 0 13192 80
rect 13304 0 13384 80
rect 13496 0 13576 80
rect 13688 0 13768 80
rect 13880 0 13960 80
rect 14072 0 14152 80
rect 14264 0 14344 80
rect 14456 0 14536 80
rect 14648 0 14728 80
rect 14840 0 14920 80
rect 15032 0 15112 80
rect 15224 0 15304 80
rect 15416 0 15496 80
rect 15608 0 15688 80
rect 15800 0 15880 80
rect 15992 0 16072 80
rect 16184 0 16264 80
rect 16376 0 16456 80
rect 16568 0 16648 80
rect 16760 0 16840 80
rect 16952 0 17032 80
rect 17144 0 17224 80
rect 17336 64 17356 80
rect 17548 80 17588 8800
rect 17740 8756 17780 8765
rect 17740 80 17780 8716
rect 17932 80 17972 9724
rect 18028 9596 18068 9605
rect 18028 8756 18068 9556
rect 18028 8707 18068 8716
rect 18124 80 18164 9808
rect 18604 9680 18644 10144
rect 18604 9631 18644 9640
rect 18700 10100 18740 10109
rect 18508 9512 18548 9521
rect 18508 9377 18548 9472
rect 18700 9176 18740 10060
rect 18808 9848 19176 9857
rect 18848 9808 18890 9848
rect 18930 9808 18972 9848
rect 19012 9808 19054 9848
rect 19094 9808 19136 9848
rect 18808 9799 19176 9808
rect 19276 9764 19316 10228
rect 19276 9715 19316 9724
rect 19372 10100 19412 10109
rect 19372 9680 19412 10060
rect 19372 9631 19412 9640
rect 19180 9596 19220 9605
rect 18700 9127 18740 9136
rect 18892 9512 18932 9521
rect 18892 9092 18932 9472
rect 19180 9176 19220 9556
rect 19180 9127 19220 9136
rect 19372 9428 19412 9437
rect 18892 9043 18932 9052
rect 18988 9008 19028 9017
rect 19028 8968 19316 9008
rect 18988 8959 19028 8968
rect 18604 8840 18644 8849
rect 18316 8756 18356 8765
rect 18220 5480 18260 5489
rect 18220 4388 18260 5440
rect 18220 4339 18260 4348
rect 18220 3968 18260 3977
rect 18220 2036 18260 3928
rect 18220 1987 18260 1996
rect 18316 80 18356 8716
rect 18412 8504 18452 8513
rect 18412 2900 18452 8464
rect 18604 5900 18644 8800
rect 18988 8840 19028 8849
rect 19180 8840 19220 8849
rect 19028 8800 19180 8840
rect 18988 8791 19028 8800
rect 19180 8791 19220 8800
rect 18808 8336 19176 8345
rect 18848 8296 18890 8336
rect 18930 8296 18972 8336
rect 19012 8296 19054 8336
rect 19094 8296 19136 8336
rect 18808 8287 19176 8296
rect 18604 5851 18644 5860
rect 18700 7748 18740 7757
rect 18700 5732 18740 7708
rect 18808 6824 19176 6833
rect 18848 6784 18890 6824
rect 18930 6784 18972 6824
rect 19012 6784 19054 6824
rect 19094 6784 19136 6824
rect 18808 6775 19176 6784
rect 18700 5683 18740 5692
rect 18796 6572 18836 6581
rect 18508 5648 18548 5657
rect 18508 4472 18548 5608
rect 18796 5480 18836 6532
rect 19276 5816 19316 8968
rect 19372 8672 19412 9388
rect 19468 8924 19508 11152
rect 20236 10772 20276 12100
rect 20236 10732 20564 10772
rect 20048 10604 20416 10613
rect 20088 10564 20130 10604
rect 20170 10564 20212 10604
rect 20252 10564 20294 10604
rect 20334 10564 20376 10604
rect 20048 10555 20416 10564
rect 19756 10184 19796 10193
rect 19468 8875 19508 8884
rect 19660 9512 19700 9521
rect 19372 8623 19412 8632
rect 19564 8840 19604 8849
rect 19468 7664 19508 7673
rect 19276 5776 19412 5816
rect 18892 5648 18932 5657
rect 18892 5513 18932 5608
rect 18700 5440 18836 5480
rect 19276 5480 19316 5489
rect 18508 4423 18548 4432
rect 18604 5396 18644 5405
rect 18604 3380 18644 5356
rect 18604 3331 18644 3340
rect 18412 2860 18548 2900
rect 18508 80 18548 2860
rect 18604 2876 18644 2885
rect 18604 2036 18644 2836
rect 18604 1987 18644 1996
rect 18700 80 18740 5440
rect 18808 5312 19176 5321
rect 18848 5272 18890 5312
rect 18930 5272 18972 5312
rect 19012 5272 19054 5312
rect 19094 5272 19136 5312
rect 18808 5263 19176 5272
rect 19084 4976 19124 4985
rect 18796 4724 18836 4733
rect 18796 4136 18836 4684
rect 19084 4640 19124 4936
rect 19084 4591 19124 4600
rect 18796 4087 18836 4096
rect 18808 3800 19176 3809
rect 18848 3760 18890 3800
rect 18930 3760 18972 3800
rect 19012 3760 19054 3800
rect 19094 3760 19136 3800
rect 18808 3751 19176 3760
rect 19276 3464 19316 5440
rect 19276 3415 19316 3424
rect 19372 2900 19412 5776
rect 19276 2860 19412 2900
rect 18892 2624 18932 2633
rect 18892 2540 18932 2584
rect 18892 2489 18932 2500
rect 18808 2288 19176 2297
rect 18848 2248 18890 2288
rect 18930 2248 18972 2288
rect 19012 2248 19054 2288
rect 19094 2248 19136 2288
rect 18808 2239 19176 2248
rect 19180 1784 19220 1793
rect 18892 1532 18932 1541
rect 18892 80 18932 1492
rect 19084 1448 19124 1457
rect 19084 80 19124 1408
rect 19180 1112 19220 1744
rect 19180 1063 19220 1072
rect 19276 80 19316 2860
rect 19372 2624 19412 2633
rect 19372 1532 19412 2584
rect 19372 1483 19412 1492
rect 19468 1532 19508 7624
rect 19468 1483 19508 1492
rect 19564 1448 19604 8800
rect 19564 1399 19604 1408
rect 19660 188 19700 9472
rect 19756 8924 19796 10144
rect 20140 10016 20180 10025
rect 20140 9596 20180 9976
rect 20524 9764 20564 10732
rect 20140 9547 20180 9556
rect 20428 9724 20564 9764
rect 20716 10268 20756 10277
rect 20428 9344 20468 9724
rect 20428 9295 20468 9304
rect 20524 9512 20564 9521
rect 20048 9092 20416 9101
rect 20088 9052 20130 9092
rect 20170 9052 20212 9092
rect 20252 9052 20294 9092
rect 20334 9052 20376 9092
rect 20048 9043 20416 9052
rect 19756 8875 19796 8884
rect 19756 7832 19796 7841
rect 19756 6488 19796 7792
rect 20048 7580 20416 7589
rect 20088 7540 20130 7580
rect 20170 7540 20212 7580
rect 20252 7540 20294 7580
rect 20334 7540 20376 7580
rect 20048 7531 20416 7540
rect 19852 7160 19892 7169
rect 19852 6740 19892 7120
rect 20524 7160 20564 9472
rect 20524 7111 20564 7120
rect 20620 8672 20660 8681
rect 19852 6691 19892 6700
rect 19756 6439 19796 6448
rect 20620 6236 20660 8632
rect 20716 8252 20756 10228
rect 20908 10016 20948 10025
rect 20908 9176 20948 9976
rect 20908 9127 20948 9136
rect 21004 9260 21044 9269
rect 21004 8840 21044 9220
rect 21004 8791 21044 8800
rect 20716 8203 20756 8212
rect 20812 7160 20852 7169
rect 20812 6656 20852 7120
rect 20812 6607 20852 6616
rect 20620 6187 20660 6196
rect 20524 6152 20564 6161
rect 20048 6068 20416 6077
rect 20088 6028 20130 6068
rect 20170 6028 20212 6068
rect 20252 6028 20294 6068
rect 20334 6028 20376 6068
rect 20048 6019 20416 6028
rect 19852 4976 19892 4985
rect 19852 4556 19892 4936
rect 19852 4507 19892 4516
rect 20048 4556 20416 4565
rect 20088 4516 20130 4556
rect 20170 4516 20212 4556
rect 20252 4516 20294 4556
rect 20334 4516 20376 4556
rect 20048 4507 20416 4516
rect 19852 4388 19892 4397
rect 19852 2900 19892 4348
rect 20140 4388 20180 4397
rect 20140 3464 20180 4348
rect 20524 4220 20564 6112
rect 21484 5480 21524 5489
rect 20524 4171 20564 4180
rect 20620 5060 20660 5069
rect 20428 4136 20468 4145
rect 20428 3632 20468 4096
rect 20428 3583 20468 3592
rect 20140 3415 20180 3424
rect 20048 3044 20416 3053
rect 20088 3004 20130 3044
rect 20170 3004 20212 3044
rect 20252 3004 20294 3044
rect 20334 3004 20376 3044
rect 20048 2995 20416 3004
rect 19852 2860 19988 2900
rect 19948 2708 19988 2860
rect 19948 2659 19988 2668
rect 20428 2456 20468 2465
rect 20428 2036 20468 2416
rect 20428 1987 20468 1996
rect 20620 1952 20660 5020
rect 21484 4976 21524 5440
rect 21484 4927 21524 4936
rect 21292 4808 21332 4817
rect 21292 4304 21332 4768
rect 21292 4255 21332 4264
rect 21004 3296 21044 3305
rect 21004 2792 21044 3256
rect 21004 2743 21044 2752
rect 20620 1903 20660 1912
rect 20524 1700 20564 1709
rect 20048 1532 20416 1541
rect 20088 1492 20130 1532
rect 20170 1492 20212 1532
rect 20252 1492 20294 1532
rect 20334 1492 20376 1532
rect 20048 1483 20416 1492
rect 20524 776 20564 1660
rect 21484 1616 21524 1625
rect 21484 1448 21524 1576
rect 21484 1399 21524 1408
rect 20524 727 20564 736
rect 19468 148 19700 188
rect 19468 80 19508 148
rect 17396 64 17416 80
rect 17336 0 17416 64
rect 17528 0 17608 80
rect 17720 0 17800 80
rect 17912 0 17992 80
rect 18104 0 18184 80
rect 18296 0 18376 80
rect 18488 0 18568 80
rect 18680 0 18760 80
rect 18872 0 18952 80
rect 19064 0 19144 80
rect 19256 0 19336 80
rect 19448 0 19528 80
<< via3 >>
rect 76 6700 116 6740
rect 76 6532 116 6572
rect 1708 6448 1748 6488
rect 2092 232 2132 272
rect 4928 10564 4968 10604
rect 5010 10564 5050 10604
rect 5092 10564 5132 10604
rect 5174 10564 5214 10604
rect 5256 10564 5296 10604
rect 2668 484 2708 524
rect 2668 148 2708 188
rect 3688 9808 3728 9848
rect 3770 9808 3810 9848
rect 3852 9808 3892 9848
rect 3934 9808 3974 9848
rect 4016 9808 4056 9848
rect 3688 8296 3728 8336
rect 3770 8296 3810 8336
rect 3852 8296 3892 8336
rect 3934 8296 3974 8336
rect 4016 8296 4056 8336
rect 3244 3928 3284 3968
rect 3244 3760 3284 3800
rect 3244 2080 3284 2120
rect 3688 6784 3728 6824
rect 3770 6784 3810 6824
rect 3852 6784 3892 6824
rect 3934 6784 3974 6824
rect 4016 6784 4056 6824
rect 3628 5440 3668 5480
rect 3688 5272 3728 5312
rect 3770 5272 3810 5312
rect 3852 5272 3892 5312
rect 3934 5272 3974 5312
rect 4016 5272 4056 5312
rect 4928 9052 4968 9092
rect 5010 9052 5050 9092
rect 5092 9052 5132 9092
rect 5174 9052 5214 9092
rect 5256 9052 5296 9092
rect 4108 3928 4148 3968
rect 3688 3760 3728 3800
rect 3770 3760 3810 3800
rect 3852 3760 3892 3800
rect 3934 3760 3974 3800
rect 4016 3760 4056 3800
rect 3688 2248 3728 2288
rect 3770 2248 3810 2288
rect 3852 2248 3892 2288
rect 3934 2248 3974 2288
rect 4016 2248 4056 2288
rect 3916 2080 3956 2120
rect 4928 7540 4968 7580
rect 5010 7540 5050 7580
rect 5092 7540 5132 7580
rect 5174 7540 5214 7580
rect 5256 7540 5296 7580
rect 4876 7120 4916 7160
rect 4928 6028 4968 6068
rect 5010 6028 5050 6068
rect 5092 6028 5132 6068
rect 5174 6028 5214 6068
rect 5256 6028 5296 6068
rect 4928 4516 4968 4556
rect 5010 4516 5050 4556
rect 5092 4516 5132 4556
rect 5174 4516 5214 4556
rect 5256 4516 5296 4556
rect 4928 3004 4968 3044
rect 5010 3004 5050 3044
rect 5092 3004 5132 3044
rect 5174 3004 5214 3044
rect 5256 3004 5296 3044
rect 4928 1492 4968 1532
rect 5010 1492 5050 1532
rect 5092 1492 5132 1532
rect 5174 1492 5214 1532
rect 5256 1492 5296 1532
rect 4876 1156 4916 1196
rect 10060 9388 10100 9428
rect 6892 316 6932 356
rect 7180 400 7220 440
rect 8044 1912 8084 1952
rect 8332 2332 8372 2372
rect 8428 1912 8468 1952
rect 13804 9472 13844 9512
rect 15244 8884 15284 8924
rect 8908 6700 8948 6740
rect 9484 7120 9524 7160
rect 9100 6532 9140 6572
rect 9100 2584 9140 2624
rect 9100 2332 9140 2372
rect 9580 2584 9620 2624
rect 9388 1156 9428 1196
rect 10636 6532 10676 6572
rect 10060 3340 10100 3380
rect 10348 4180 10388 4220
rect 10156 1240 10196 1280
rect 11692 2500 11732 2540
rect 11980 2416 12020 2456
rect 12940 4180 12980 4220
rect 13036 2584 13076 2624
rect 15628 8884 15668 8924
rect 13516 2584 13556 2624
rect 14476 5608 14516 5648
rect 14572 2332 14612 2372
rect 16012 2332 16052 2372
rect 16204 1240 16244 1280
rect 15820 484 15860 524
rect 15628 148 15668 188
rect 16012 232 16052 272
rect 16492 400 16532 440
rect 17068 6532 17108 6572
rect 17356 6448 17396 6488
rect 17068 3340 17108 3380
rect 16780 2416 16820 2456
rect 16780 316 16820 356
rect 18508 9472 18548 9512
rect 18808 9808 18848 9848
rect 18890 9808 18930 9848
rect 18972 9808 19012 9848
rect 19054 9808 19094 9848
rect 19136 9808 19176 9848
rect 19372 9388 19412 9428
rect 18808 8296 18848 8336
rect 18890 8296 18930 8336
rect 18972 8296 19012 8336
rect 19054 8296 19094 8336
rect 19136 8296 19176 8336
rect 18808 6784 18848 6824
rect 18890 6784 18930 6824
rect 18972 6784 19012 6824
rect 19054 6784 19094 6824
rect 19136 6784 19176 6824
rect 20048 10564 20088 10604
rect 20130 10564 20170 10604
rect 20212 10564 20252 10604
rect 20294 10564 20334 10604
rect 20376 10564 20416 10604
rect 18892 5608 18932 5648
rect 18808 5272 18848 5312
rect 18890 5272 18930 5312
rect 18972 5272 19012 5312
rect 19054 5272 19094 5312
rect 19136 5272 19176 5312
rect 18808 3760 18848 3800
rect 18890 3760 18930 3800
rect 18972 3760 19012 3800
rect 19054 3760 19094 3800
rect 19136 3760 19176 3800
rect 18892 2500 18932 2540
rect 18808 2248 18848 2288
rect 18890 2248 18930 2288
rect 18972 2248 19012 2288
rect 19054 2248 19094 2288
rect 19136 2248 19176 2288
rect 18892 1492 18932 1532
rect 19084 1408 19124 1448
rect 19468 1492 19508 1532
rect 19564 1408 19604 1448
rect 20048 9052 20088 9092
rect 20130 9052 20170 9092
rect 20212 9052 20252 9092
rect 20294 9052 20334 9092
rect 20376 9052 20416 9092
rect 20048 7540 20088 7580
rect 20130 7540 20170 7580
rect 20212 7540 20252 7580
rect 20294 7540 20334 7580
rect 20376 7540 20416 7580
rect 20048 6028 20088 6068
rect 20130 6028 20170 6068
rect 20212 6028 20252 6068
rect 20294 6028 20334 6068
rect 20376 6028 20416 6068
rect 20048 4516 20088 4556
rect 20130 4516 20170 4556
rect 20212 4516 20252 4556
rect 20294 4516 20334 4556
rect 20376 4516 20416 4556
rect 20048 3004 20088 3044
rect 20130 3004 20170 3044
rect 20212 3004 20252 3044
rect 20294 3004 20334 3044
rect 20376 3004 20416 3044
rect 20048 1492 20088 1532
rect 20130 1492 20170 1532
rect 20212 1492 20252 1532
rect 20294 1492 20334 1532
rect 20376 1492 20416 1532
<< metal4 >>
rect 4919 10564 4928 10604
rect 4968 10564 5010 10604
rect 5050 10564 5092 10604
rect 5132 10564 5174 10604
rect 5214 10564 5256 10604
rect 5296 10564 5305 10604
rect 20039 10564 20048 10604
rect 20088 10564 20130 10604
rect 20170 10564 20212 10604
rect 20252 10564 20294 10604
rect 20334 10564 20376 10604
rect 20416 10564 20425 10604
rect 3679 9808 3688 9848
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 4056 9808 4065 9848
rect 18799 9808 18808 9848
rect 18848 9808 18890 9848
rect 18930 9808 18972 9848
rect 19012 9808 19054 9848
rect 19094 9808 19136 9848
rect 19176 9808 19185 9848
rect 13795 9472 13804 9512
rect 13844 9472 18508 9512
rect 18548 9472 18557 9512
rect 10051 9388 10060 9428
rect 10100 9388 19372 9428
rect 19412 9388 19421 9428
rect 4919 9052 4928 9092
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 5296 9052 5305 9092
rect 20039 9052 20048 9092
rect 20088 9052 20130 9092
rect 20170 9052 20212 9092
rect 20252 9052 20294 9092
rect 20334 9052 20376 9092
rect 20416 9052 20425 9092
rect 15235 8884 15244 8924
rect 15284 8884 15628 8924
rect 15668 8884 15677 8924
rect 3679 8296 3688 8336
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 4056 8296 4065 8336
rect 18799 8296 18808 8336
rect 18848 8296 18890 8336
rect 18930 8296 18972 8336
rect 19012 8296 19054 8336
rect 19094 8296 19136 8336
rect 19176 8296 19185 8336
rect 4919 7540 4928 7580
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 5296 7540 5305 7580
rect 20039 7540 20048 7580
rect 20088 7540 20130 7580
rect 20170 7540 20212 7580
rect 20252 7540 20294 7580
rect 20334 7540 20376 7580
rect 20416 7540 20425 7580
rect 4867 7120 4876 7160
rect 4916 7120 9484 7160
rect 9524 7120 9533 7160
rect 3679 6784 3688 6824
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 4056 6784 4065 6824
rect 18799 6784 18808 6824
rect 18848 6784 18890 6824
rect 18930 6784 18972 6824
rect 19012 6784 19054 6824
rect 19094 6784 19136 6824
rect 19176 6784 19185 6824
rect 67 6700 76 6740
rect 116 6700 8908 6740
rect 8948 6700 8957 6740
rect 67 6532 76 6572
rect 116 6532 9100 6572
rect 9140 6532 9149 6572
rect 10627 6532 10636 6572
rect 10676 6532 17068 6572
rect 17108 6532 17117 6572
rect 1699 6448 1708 6488
rect 1748 6448 17356 6488
rect 17396 6448 17405 6488
rect 4919 6028 4928 6068
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 5296 6028 5305 6068
rect 20039 6028 20048 6068
rect 20088 6028 20130 6068
rect 20170 6028 20212 6068
rect 20252 6028 20294 6068
rect 20334 6028 20376 6068
rect 20416 6028 20425 6068
rect 14467 5608 14476 5648
rect 14516 5608 18892 5648
rect 18932 5608 18941 5648
rect 3235 5440 3244 5480
rect 3284 5440 3628 5480
rect 3668 5440 3677 5480
rect 3679 5272 3688 5312
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 4056 5272 4065 5312
rect 18799 5272 18808 5312
rect 18848 5272 18890 5312
rect 18930 5272 18972 5312
rect 19012 5272 19054 5312
rect 19094 5272 19136 5312
rect 19176 5272 19185 5312
rect 4919 4516 4928 4556
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 5296 4516 5305 4556
rect 20039 4516 20048 4556
rect 20088 4516 20130 4556
rect 20170 4516 20212 4556
rect 20252 4516 20294 4556
rect 20334 4516 20376 4556
rect 20416 4516 20425 4556
rect 10339 4180 10348 4220
rect 10388 4180 12940 4220
rect 12980 4180 12989 4220
rect 3235 3928 3244 3968
rect 3284 3928 4108 3968
rect 4148 3928 4157 3968
rect 3149 3760 3244 3800
rect 3284 3760 3293 3800
rect 3679 3760 3688 3800
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 4056 3760 4065 3800
rect 18799 3760 18808 3800
rect 18848 3760 18890 3800
rect 18930 3760 18972 3800
rect 19012 3760 19054 3800
rect 19094 3760 19136 3800
rect 19176 3760 19185 3800
rect 10051 3340 10060 3380
rect 10100 3340 17068 3380
rect 17108 3340 17117 3380
rect 4919 3004 4928 3044
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 5296 3004 5305 3044
rect 20039 3004 20048 3044
rect 20088 3004 20130 3044
rect 20170 3004 20212 3044
rect 20252 3004 20294 3044
rect 20334 3004 20376 3044
rect 20416 3004 20425 3044
rect 9091 2584 9100 2624
rect 9140 2584 9580 2624
rect 9620 2584 9629 2624
rect 13027 2584 13036 2624
rect 13076 2584 13516 2624
rect 13556 2584 13565 2624
rect 11683 2500 11692 2540
rect 11732 2500 18892 2540
rect 18932 2500 18941 2540
rect 11971 2416 11980 2456
rect 12020 2416 16780 2456
rect 16820 2416 16829 2456
rect 8323 2332 8332 2372
rect 8372 2332 9100 2372
rect 9140 2332 9149 2372
rect 14563 2332 14572 2372
rect 14612 2332 16012 2372
rect 16052 2332 16061 2372
rect 3679 2248 3688 2288
rect 3728 2248 3770 2288
rect 3810 2248 3852 2288
rect 3892 2248 3934 2288
rect 3974 2248 4016 2288
rect 4056 2248 4065 2288
rect 18799 2248 18808 2288
rect 18848 2248 18890 2288
rect 18930 2248 18972 2288
rect 19012 2248 19054 2288
rect 19094 2248 19136 2288
rect 19176 2248 19185 2288
rect 3235 2080 3244 2120
rect 3284 2080 3916 2120
rect 3956 2080 3965 2120
rect 8035 1912 8044 1952
rect 8084 1912 8428 1952
rect 8468 1912 8477 1952
rect 4919 1492 4928 1532
rect 4968 1492 5010 1532
rect 5050 1492 5092 1532
rect 5132 1492 5174 1532
rect 5214 1492 5256 1532
rect 5296 1492 5305 1532
rect 18883 1492 18892 1532
rect 18932 1492 19468 1532
rect 19508 1492 19517 1532
rect 20039 1492 20048 1532
rect 20088 1492 20130 1532
rect 20170 1492 20212 1532
rect 20252 1492 20294 1532
rect 20334 1492 20376 1532
rect 20416 1492 20425 1532
rect 19075 1408 19084 1448
rect 19124 1408 19564 1448
rect 19604 1408 19613 1448
rect 10147 1240 10156 1280
rect 10196 1240 16204 1280
rect 16244 1240 16253 1280
rect 4867 1156 4876 1196
rect 4916 1156 9388 1196
rect 9428 1156 9437 1196
rect 2659 484 2668 524
rect 2708 484 15820 524
rect 15860 484 15869 524
rect 7171 400 7180 440
rect 7220 400 16492 440
rect 16532 400 16541 440
rect 6883 316 6892 356
rect 6932 316 16780 356
rect 16820 316 16829 356
rect 2083 232 2092 272
rect 2132 232 16012 272
rect 16052 232 16061 272
rect 2659 148 2668 188
rect 2708 148 15628 188
rect 15668 148 15677 188
<< via4 >>
rect 4928 10564 4968 10604
rect 5010 10564 5050 10604
rect 5092 10564 5132 10604
rect 5174 10564 5214 10604
rect 5256 10564 5296 10604
rect 20048 10564 20088 10604
rect 20130 10564 20170 10604
rect 20212 10564 20252 10604
rect 20294 10564 20334 10604
rect 20376 10564 20416 10604
rect 3688 9808 3728 9848
rect 3770 9808 3810 9848
rect 3852 9808 3892 9848
rect 3934 9808 3974 9848
rect 4016 9808 4056 9848
rect 18808 9808 18848 9848
rect 18890 9808 18930 9848
rect 18972 9808 19012 9848
rect 19054 9808 19094 9848
rect 19136 9808 19176 9848
rect 4928 9052 4968 9092
rect 5010 9052 5050 9092
rect 5092 9052 5132 9092
rect 5174 9052 5214 9092
rect 5256 9052 5296 9092
rect 20048 9052 20088 9092
rect 20130 9052 20170 9092
rect 20212 9052 20252 9092
rect 20294 9052 20334 9092
rect 20376 9052 20416 9092
rect 3688 8296 3728 8336
rect 3770 8296 3810 8336
rect 3852 8296 3892 8336
rect 3934 8296 3974 8336
rect 4016 8296 4056 8336
rect 18808 8296 18848 8336
rect 18890 8296 18930 8336
rect 18972 8296 19012 8336
rect 19054 8296 19094 8336
rect 19136 8296 19176 8336
rect 4928 7540 4968 7580
rect 5010 7540 5050 7580
rect 5092 7540 5132 7580
rect 5174 7540 5214 7580
rect 5256 7540 5296 7580
rect 20048 7540 20088 7580
rect 20130 7540 20170 7580
rect 20212 7540 20252 7580
rect 20294 7540 20334 7580
rect 20376 7540 20416 7580
rect 3688 6784 3728 6824
rect 3770 6784 3810 6824
rect 3852 6784 3892 6824
rect 3934 6784 3974 6824
rect 4016 6784 4056 6824
rect 18808 6784 18848 6824
rect 18890 6784 18930 6824
rect 18972 6784 19012 6824
rect 19054 6784 19094 6824
rect 19136 6784 19176 6824
rect 4928 6028 4968 6068
rect 5010 6028 5050 6068
rect 5092 6028 5132 6068
rect 5174 6028 5214 6068
rect 5256 6028 5296 6068
rect 20048 6028 20088 6068
rect 20130 6028 20170 6068
rect 20212 6028 20252 6068
rect 20294 6028 20334 6068
rect 20376 6028 20416 6068
rect 3244 5440 3284 5480
rect 3688 5272 3728 5312
rect 3770 5272 3810 5312
rect 3852 5272 3892 5312
rect 3934 5272 3974 5312
rect 4016 5272 4056 5312
rect 18808 5272 18848 5312
rect 18890 5272 18930 5312
rect 18972 5272 19012 5312
rect 19054 5272 19094 5312
rect 19136 5272 19176 5312
rect 4928 4516 4968 4556
rect 5010 4516 5050 4556
rect 5092 4516 5132 4556
rect 5174 4516 5214 4556
rect 5256 4516 5296 4556
rect 20048 4516 20088 4556
rect 20130 4516 20170 4556
rect 20212 4516 20252 4556
rect 20294 4516 20334 4556
rect 20376 4516 20416 4556
rect 3244 3760 3284 3800
rect 3688 3760 3728 3800
rect 3770 3760 3810 3800
rect 3852 3760 3892 3800
rect 3934 3760 3974 3800
rect 4016 3760 4056 3800
rect 18808 3760 18848 3800
rect 18890 3760 18930 3800
rect 18972 3760 19012 3800
rect 19054 3760 19094 3800
rect 19136 3760 19176 3800
rect 4928 3004 4968 3044
rect 5010 3004 5050 3044
rect 5092 3004 5132 3044
rect 5174 3004 5214 3044
rect 5256 3004 5296 3044
rect 20048 3004 20088 3044
rect 20130 3004 20170 3044
rect 20212 3004 20252 3044
rect 20294 3004 20334 3044
rect 20376 3004 20416 3044
rect 3688 2248 3728 2288
rect 3770 2248 3810 2288
rect 3852 2248 3892 2288
rect 3934 2248 3974 2288
rect 4016 2248 4056 2288
rect 18808 2248 18848 2288
rect 18890 2248 18930 2288
rect 18972 2248 19012 2288
rect 19054 2248 19094 2288
rect 19136 2248 19176 2288
rect 4928 1492 4968 1532
rect 5010 1492 5050 1532
rect 5092 1492 5132 1532
rect 5174 1492 5214 1532
rect 5256 1492 5296 1532
rect 20048 1492 20088 1532
rect 20130 1492 20170 1532
rect 20212 1492 20252 1532
rect 20294 1492 20334 1532
rect 20376 1492 20416 1532
<< metal5 >>
rect 3652 9848 4092 12180
rect 3652 9808 3688 9848
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 4056 9808 4092 9848
rect 3652 8336 4092 9808
rect 3652 8296 3688 8336
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 4056 8296 4092 8336
rect 3652 6824 4092 8296
rect 3652 6784 3688 6824
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 4056 6784 4092 6824
rect 3244 5480 3284 5489
rect 3244 3800 3284 5440
rect 3244 3751 3284 3760
rect 3652 5312 4092 6784
rect 3652 5272 3688 5312
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 4056 5272 4092 5312
rect 3652 3800 4092 5272
rect 3652 3760 3688 3800
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 4056 3760 4092 3800
rect 3652 2288 4092 3760
rect 3652 2248 3688 2288
rect 3728 2248 3770 2288
rect 3810 2248 3852 2288
rect 3892 2248 3934 2288
rect 3974 2248 4016 2288
rect 4056 2248 4092 2288
rect 3652 0 4092 2248
rect 4892 10604 5332 12180
rect 4892 10564 4928 10604
rect 4968 10564 5010 10604
rect 5050 10564 5092 10604
rect 5132 10564 5174 10604
rect 5214 10564 5256 10604
rect 5296 10564 5332 10604
rect 4892 9092 5332 10564
rect 4892 9052 4928 9092
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 5296 9052 5332 9092
rect 4892 7580 5332 9052
rect 4892 7540 4928 7580
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 5296 7540 5332 7580
rect 4892 6068 5332 7540
rect 4892 6028 4928 6068
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 5296 6028 5332 6068
rect 4892 4556 5332 6028
rect 4892 4516 4928 4556
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 5296 4516 5332 4556
rect 4892 3044 5332 4516
rect 4892 3004 4928 3044
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 5296 3004 5332 3044
rect 4892 1532 5332 3004
rect 4892 1492 4928 1532
rect 4968 1492 5010 1532
rect 5050 1492 5092 1532
rect 5132 1492 5174 1532
rect 5214 1492 5256 1532
rect 5296 1492 5332 1532
rect 4892 0 5332 1492
rect 18772 9848 19212 12180
rect 18772 9808 18808 9848
rect 18848 9808 18890 9848
rect 18930 9808 18972 9848
rect 19012 9808 19054 9848
rect 19094 9808 19136 9848
rect 19176 9808 19212 9848
rect 18772 8336 19212 9808
rect 18772 8296 18808 8336
rect 18848 8296 18890 8336
rect 18930 8296 18972 8336
rect 19012 8296 19054 8336
rect 19094 8296 19136 8336
rect 19176 8296 19212 8336
rect 18772 6824 19212 8296
rect 18772 6784 18808 6824
rect 18848 6784 18890 6824
rect 18930 6784 18972 6824
rect 19012 6784 19054 6824
rect 19094 6784 19136 6824
rect 19176 6784 19212 6824
rect 18772 5312 19212 6784
rect 18772 5272 18808 5312
rect 18848 5272 18890 5312
rect 18930 5272 18972 5312
rect 19012 5272 19054 5312
rect 19094 5272 19136 5312
rect 19176 5272 19212 5312
rect 18772 3800 19212 5272
rect 18772 3760 18808 3800
rect 18848 3760 18890 3800
rect 18930 3760 18972 3800
rect 19012 3760 19054 3800
rect 19094 3760 19136 3800
rect 19176 3760 19212 3800
rect 18772 2288 19212 3760
rect 18772 2248 18808 2288
rect 18848 2248 18890 2288
rect 18930 2248 18972 2288
rect 19012 2248 19054 2288
rect 19094 2248 19136 2288
rect 19176 2248 19212 2288
rect 18772 0 19212 2248
rect 20012 10604 20452 12180
rect 20012 10564 20048 10604
rect 20088 10564 20130 10604
rect 20170 10564 20212 10604
rect 20252 10564 20294 10604
rect 20334 10564 20376 10604
rect 20416 10564 20452 10604
rect 20012 9092 20452 10564
rect 20012 9052 20048 9092
rect 20088 9052 20130 9092
rect 20170 9052 20212 9092
rect 20252 9052 20294 9092
rect 20334 9052 20376 9092
rect 20416 9052 20452 9092
rect 20012 7580 20452 9052
rect 20012 7540 20048 7580
rect 20088 7540 20130 7580
rect 20170 7540 20212 7580
rect 20252 7540 20294 7580
rect 20334 7540 20376 7580
rect 20416 7540 20452 7580
rect 20012 6068 20452 7540
rect 20012 6028 20048 6068
rect 20088 6028 20130 6068
rect 20170 6028 20212 6068
rect 20252 6028 20294 6068
rect 20334 6028 20376 6068
rect 20416 6028 20452 6068
rect 20012 4556 20452 6028
rect 20012 4516 20048 4556
rect 20088 4516 20130 4556
rect 20170 4516 20212 4556
rect 20252 4516 20294 4556
rect 20334 4516 20376 4556
rect 20416 4516 20452 4556
rect 20012 3044 20452 4516
rect 20012 3004 20048 3044
rect 20088 3004 20130 3044
rect 20170 3004 20212 3044
rect 20252 3004 20294 3044
rect 20334 3004 20376 3044
rect 20416 3004 20452 3044
rect 20012 1532 20452 3004
rect 20012 1492 20048 1532
rect 20088 1492 20130 1532
rect 20170 1492 20212 1532
rect 20252 1492 20294 1532
rect 20334 1492 20376 1532
rect 20416 1492 20452 1532
rect 20012 0 20452 1492
use sg13g2_buf_1  _00_
timestamp 1676381911
transform 1 0 16896 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _01_
timestamp 1676381911
transform 1 0 17280 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _02_
timestamp 1676381911
transform -1 0 19584 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _03_
timestamp 1676381911
transform -1 0 19968 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _04_
timestamp 1676381911
transform 1 0 18816 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _05_
timestamp 1676381911
transform 1 0 19008 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _06_
timestamp 1676381911
transform 1 0 18816 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _07_
timestamp 1676381911
transform 1 0 16896 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _08_
timestamp 1676381911
transform 1 0 15648 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _09_
timestamp 1676381911
transform 1 0 16992 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _10_
timestamp 1676381911
transform 1 0 19392 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _11_
timestamp 1676381911
transform 1 0 18432 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _12_
timestamp 1676381911
transform 1 0 16992 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _13_
timestamp 1676381911
transform 1 0 17856 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _14_
timestamp 1676381911
transform 1 0 14400 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _15_
timestamp 1676381911
transform 1 0 16608 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _16_
timestamp 1676381911
transform 1 0 17184 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _17_
timestamp 1676381911
transform 1 0 16992 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _18_
timestamp 1676381911
transform 1 0 8832 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _19_
timestamp 1676381911
transform 1 0 19392 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _20_
timestamp 1676381911
transform 1 0 12768 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _21_
timestamp 1676381911
transform 1 0 5952 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _22_
timestamp 1676381911
transform 1 0 19200 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _23_
timestamp 1676381911
transform 1 0 6144 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _24_
timestamp 1676381911
transform 1 0 19776 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _25_
timestamp 1676381911
transform 1 0 15264 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _26_
timestamp 1676381911
transform 1 0 19296 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _27_
timestamp 1676381911
transform 1 0 13728 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _28_
timestamp 1676381911
transform 1 0 13344 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _29_
timestamp 1676381911
transform 1 0 2400 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _30_
timestamp 1676381911
transform 1 0 11232 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  _31_
timestamp 1676381911
transform -1 0 19584 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  _32_
timestamp 1676381911
transform -1 0 2304 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _33_
timestamp 1676381911
transform 1 0 2016 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _34_
timestamp 1676381911
transform 1 0 3552 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _35_
timestamp 1676381911
transform -1 0 5568 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _36_
timestamp 1676381911
transform 1 0 4800 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _37_
timestamp 1676381911
transform -1 0 7104 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _38_
timestamp 1676381911
transform -1 0 8736 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _39_
timestamp 1676381911
transform 1 0 7584 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _40_
timestamp 1676381911
transform 1 0 8736 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _41_
timestamp 1676381911
transform -1 0 11232 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  _42_
timestamp 1676381911
transform -1 0 13344 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _43_
timestamp 1676381911
transform -1 0 14496 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  _44_
timestamp 1676381911
transform -1 0 14112 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  _45_
timestamp 1676381911
transform -1 0 15168 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  _46_
timestamp 1676381911
transform -1 0 15744 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _47_
timestamp 1676381911
transform 1 0 15168 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _48_
timestamp 1676381911
transform 1 0 15648 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _49_
timestamp 1676381911
transform 1 0 16320 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  _50_
timestamp 1676381911
transform 1 0 17472 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  _51_
timestamp 1676381911
transform -1 0 19968 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  _52_
timestamp 1676381911
transform 1 0 4896 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _53_
timestamp 1676381911
transform 1 0 1920 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _54_
timestamp 1676381911
transform 1 0 2400 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _55_
timestamp 1676381911
transform 1 0 2016 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _56_
timestamp 1676381911
transform 1 0 7680 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _57_
timestamp 1676381911
transform 1 0 7296 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _58_
timestamp 1676381911
transform 1 0 6144 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _59_
timestamp 1676381911
transform 1 0 4608 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _60_
timestamp 1676381911
transform 1 0 3456 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _61_
timestamp 1676381911
transform 1 0 2016 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _62_
timestamp 1676381911
transform 1 0 2208 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _63_
timestamp 1676381911
transform 1 0 2400 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _64_
timestamp 1676381911
transform 1 0 9024 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _65_
timestamp 1676381911
transform 1 0 8640 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _66_
timestamp 1676381911
transform 1 0 8928 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _67_
timestamp 1676381911
transform 1 0 9312 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _68_
timestamp 1676381911
transform 1 0 9888 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _69_
timestamp 1676381911
transform 1 0 8928 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _70_
timestamp 1676381911
transform 1 0 4416 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _71_
timestamp 1676381911
transform 1 0 1824 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _72_
timestamp 1676381911
transform -1 0 14784 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _73_
timestamp 1676381911
transform -1 0 14400 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _74_
timestamp 1676381911
transform -1 0 13728 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _75_
timestamp 1676381911
transform 1 0 11904 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _76_
timestamp 1676381911
transform 1 0 10176 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _77_
timestamp 1676381911
transform 1 0 10560 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _78_
timestamp 1676381911
transform 1 0 11520 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _79_
timestamp 1676381911
transform -1 0 16512 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _80_
timestamp 1676381911
transform -1 0 15840 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _81_
timestamp 1676381911
transform -1 0 16896 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _82_
timestamp 1676381911
transform -1 0 15744 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _83_
timestamp 1676381911
transform -1 0 16128 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _84_
timestamp 1676381911
transform -1 0 17184 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _85_
timestamp 1676381911
transform -1 0 18048 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _86_
timestamp 1676381911
transform -1 0 19776 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _87_
timestamp 1676381911
transform -1 0 19680 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _88_
timestamp 1676381911
transform -1 0 2688 0 1 9072
box -48 -56 432 834
use sg13g2_decap_8  FILLER_0_0
timestamp 1679581782
transform 1 0 1152 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_7
timestamp 1679581782
transform 1 0 1824 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_14
timestamp 1679581782
transform 1 0 2496 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_21
timestamp 1679581782
transform 1 0 3168 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_28
timestamp 1679581782
transform 1 0 3840 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_35
timestamp 1679581782
transform 1 0 4512 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_42
timestamp 1679581782
transform 1 0 5184 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_49
timestamp 1679581782
transform 1 0 5856 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_56
timestamp 1679581782
transform 1 0 6528 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_63
timestamp 1679581782
transform 1 0 7200 0 1 1512
box -48 -56 720 834
use sg13g2_fill_2  FILLER_0_70
timestamp 1677580104
transform 1 0 7872 0 1 1512
box -48 -56 240 834
use sg13g2_fill_1  FILLER_0_72
timestamp 1677579658
transform 1 0 8064 0 1 1512
box -48 -56 144 834
use sg13g2_decap_8  FILLER_0_165
timestamp 1679581782
transform 1 0 16992 0 1 1512
box -48 -56 720 834
use sg13g2_decap_4  FILLER_0_172
timestamp 1679577901
transform 1 0 17664 0 1 1512
box -48 -56 432 834
use sg13g2_fill_1  FILLER_0_176
timestamp 1677579658
transform 1 0 18048 0 1 1512
box -48 -56 144 834
use sg13g2_decap_8  FILLER_1_0
timestamp 1679581782
transform 1 0 1152 0 -1 3024
box -48 -56 720 834
use sg13g2_fill_2  FILLER_1_7
timestamp 1677580104
transform 1 0 1824 0 -1 3024
box -48 -56 240 834
use sg13g2_decap_8  FILLER_1_17
timestamp 1679581782
transform 1 0 2784 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_24
timestamp 1679581782
transform 1 0 3456 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_31
timestamp 1679581782
transform 1 0 4128 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_38
timestamp 1679581782
transform 1 0 4800 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_45
timestamp 1679581782
transform 1 0 5472 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_52
timestamp 1679581782
transform 1 0 6144 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_59
timestamp 1679581782
transform 1 0 6816 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_66
timestamp 1679581782
transform 1 0 7488 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_73
timestamp 1679581782
transform 1 0 8160 0 -1 3024
box -48 -56 720 834
use sg13g2_fill_1  FILLER_1_80
timestamp 1677579658
transform 1 0 8832 0 -1 3024
box -48 -56 144 834
use sg13g2_decap_8  FILLER_1_105
timestamp 1679581782
transform 1 0 11232 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_112
timestamp 1679581782
transform 1 0 11904 0 -1 3024
box -48 -56 720 834
use sg13g2_fill_1  FILLER_1_147
timestamp 1677579658
transform 1 0 15264 0 -1 3024
box -48 -56 144 834
use sg13g2_decap_4  FILLER_1_156
timestamp 1679577901
transform 1 0 16128 0 -1 3024
box -48 -56 432 834
use sg13g2_decap_8  FILLER_1_172
timestamp 1679581782
transform 1 0 17664 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_4  FILLER_1_179
timestamp 1679577901
transform 1 0 18336 0 -1 3024
box -48 -56 432 834
use sg13g2_fill_1  FILLER_1_183
timestamp 1677579658
transform 1 0 18720 0 -1 3024
box -48 -56 144 834
use sg13g2_fill_1  FILLER_1_196
timestamp 1677579658
transform 1 0 19968 0 -1 3024
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_0
timestamp 1679581782
transform 1 0 1152 0 1 3024
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_7
timestamp 1679577901
transform 1 0 1824 0 1 3024
box -48 -56 432 834
use sg13g2_fill_2  FILLER_2_11
timestamp 1677580104
transform 1 0 2208 0 1 3024
box -48 -56 240 834
use sg13g2_decap_8  FILLER_2_17
timestamp 1679581782
transform 1 0 2784 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_24
timestamp 1679581782
transform 1 0 3456 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_31
timestamp 1679581782
transform 1 0 4128 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_38
timestamp 1679581782
transform 1 0 4800 0 1 3024
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_45
timestamp 1679577901
transform 1 0 5472 0 1 3024
box -48 -56 432 834
use sg13g2_fill_1  FILLER_2_49
timestamp 1677579658
transform 1 0 5856 0 1 3024
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_54
timestamp 1679581782
transform 1 0 6336 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_61
timestamp 1679581782
transform 1 0 7008 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_68
timestamp 1679581782
transform 1 0 7680 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_75
timestamp 1679581782
transform 1 0 8352 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_82
timestamp 1679581782
transform 1 0 9024 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_89
timestamp 1679581782
transform 1 0 9696 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_96
timestamp 1679581782
transform 1 0 10368 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_103
timestamp 1679581782
transform 1 0 11040 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_110
timestamp 1679581782
transform 1 0 11712 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_117
timestamp 1679581782
transform 1 0 12384 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_124
timestamp 1679581782
transform 1 0 13056 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_131
timestamp 1679581782
transform 1 0 13728 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_138
timestamp 1679581782
transform 1 0 14400 0 1 3024
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_145
timestamp 1679577901
transform 1 0 15072 0 1 3024
box -48 -56 432 834
use sg13g2_decap_8  FILLER_2_153
timestamp 1679581782
transform 1 0 15840 0 1 3024
box -48 -56 720 834
use sg13g2_fill_2  FILLER_2_160
timestamp 1677580104
transform 1 0 16512 0 1 3024
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_162
timestamp 1677579658
transform 1 0 16704 0 1 3024
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_167
timestamp 1679581782
transform 1 0 17184 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_174
timestamp 1679581782
transform 1 0 17856 0 1 3024
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_181
timestamp 1679577901
transform 1 0 18528 0 1 3024
box -48 -56 432 834
use sg13g2_decap_8  FILLER_3_0
timestamp 1679581782
transform 1 0 1152 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_7
timestamp 1679577901
transform 1 0 1824 0 -1 4536
box -48 -56 432 834
use sg13g2_decap_8  FILLER_3_15
timestamp 1679581782
transform 1 0 2592 0 -1 4536
box -48 -56 720 834
use sg13g2_fill_2  FILLER_3_22
timestamp 1677580104
transform 1 0 3264 0 -1 4536
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_24
timestamp 1677579658
transform 1 0 3456 0 -1 4536
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_29
timestamp 1679581782
transform 1 0 3936 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_36
timestamp 1679581782
transform 1 0 4608 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_43
timestamp 1679581782
transform 1 0 5280 0 -1 4536
box -48 -56 720 834
use sg13g2_fill_2  FILLER_3_50
timestamp 1677580104
transform 1 0 5952 0 -1 4536
box -48 -56 240 834
use sg13g2_decap_8  FILLER_3_56
timestamp 1679581782
transform 1 0 6528 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_63
timestamp 1679581782
transform 1 0 7200 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_70
timestamp 1679581782
transform 1 0 7872 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_77
timestamp 1679581782
transform 1 0 8544 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_84
timestamp 1679581782
transform 1 0 9216 0 -1 4536
box -48 -56 720 834
use sg13g2_fill_2  FILLER_3_91
timestamp 1677580104
transform 1 0 9888 0 -1 4536
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_93
timestamp 1677579658
transform 1 0 10080 0 -1 4536
box -48 -56 144 834
use sg13g2_decap_4  FILLER_3_102
timestamp 1679577901
transform 1 0 10944 0 -1 4536
box -48 -56 432 834
use sg13g2_fill_2  FILLER_3_106
timestamp 1677580104
transform 1 0 11328 0 -1 4536
box -48 -56 240 834
use sg13g2_decap_8  FILLER_3_116
timestamp 1679581782
transform 1 0 12288 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_123
timestamp 1679577901
transform 1 0 12960 0 -1 4536
box -48 -56 432 834
use sg13g2_fill_2  FILLER_3_131
timestamp 1677580104
transform 1 0 13728 0 -1 4536
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_133
timestamp 1677579658
transform 1 0 13920 0 -1 4536
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_142
timestamp 1679581782
transform 1 0 14784 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_149
timestamp 1679581782
transform 1 0 15456 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_160
timestamp 1679581782
transform 1 0 16512 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_167
timestamp 1679577901
transform 1 0 17184 0 -1 4536
box -48 -56 432 834
use sg13g2_fill_1  FILLER_3_171
timestamp 1677579658
transform 1 0 17568 0 -1 4536
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_176
timestamp 1679581782
transform 1 0 18048 0 -1 4536
box -48 -56 720 834
use sg13g2_fill_2  FILLER_3_183
timestamp 1677580104
transform 1 0 18720 0 -1 4536
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_185
timestamp 1677579658
transform 1 0 18912 0 -1 4536
box -48 -56 144 834
use sg13g2_fill_2  FILLER_3_194
timestamp 1677580104
transform 1 0 19776 0 -1 4536
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_196
timestamp 1677579658
transform 1 0 19968 0 -1 4536
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_0
timestamp 1679581782
transform 1 0 1152 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_7
timestamp 1679581782
transform 1 0 1824 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_14
timestamp 1679581782
transform 1 0 2496 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_21
timestamp 1679581782
transform 1 0 3168 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_28
timestamp 1679581782
transform 1 0 3840 0 1 4536
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_35
timestamp 1679577901
transform 1 0 4512 0 1 4536
box -48 -56 432 834
use sg13g2_decap_8  FILLER_4_43
timestamp 1679581782
transform 1 0 5280 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_50
timestamp 1679581782
transform 1 0 5952 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_57
timestamp 1679581782
transform 1 0 6624 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_64
timestamp 1679581782
transform 1 0 7296 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_71
timestamp 1679581782
transform 1 0 7968 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_86
timestamp 1679581782
transform 1 0 9408 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_93
timestamp 1679581782
transform 1 0 10080 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_100
timestamp 1679581782
transform 1 0 10752 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_107
timestamp 1679581782
transform 1 0 11424 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_114
timestamp 1679581782
transform 1 0 12096 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_121
timestamp 1679581782
transform 1 0 12768 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_128
timestamp 1679581782
transform 1 0 13440 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_135
timestamp 1679581782
transform 1 0 14112 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_142
timestamp 1679581782
transform 1 0 14784 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_149
timestamp 1679581782
transform 1 0 15456 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_156
timestamp 1679581782
transform 1 0 16128 0 1 4536
box -48 -56 720 834
use sg13g2_fill_2  FILLER_4_163
timestamp 1677580104
transform 1 0 16800 0 1 4536
box -48 -56 240 834
use sg13g2_decap_8  FILLER_4_169
timestamp 1679581782
transform 1 0 17376 0 1 4536
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_176
timestamp 1679577901
transform 1 0 18048 0 1 4536
box -48 -56 432 834
use sg13g2_fill_2  FILLER_4_180
timestamp 1677580104
transform 1 0 18432 0 1 4536
box -48 -56 240 834
use sg13g2_fill_2  FILLER_4_194
timestamp 1677580104
transform 1 0 19776 0 1 4536
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_196
timestamp 1677579658
transform 1 0 19968 0 1 4536
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_0
timestamp 1679581782
transform 1 0 1152 0 -1 6048
box -48 -56 720 834
use sg13g2_fill_1  FILLER_5_7
timestamp 1677579658
transform 1 0 1824 0 -1 6048
box -48 -56 144 834
use sg13g2_fill_1  FILLER_5_12
timestamp 1677579658
transform 1 0 2304 0 -1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_17
timestamp 1679581782
transform 1 0 2784 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_24
timestamp 1679581782
transform 1 0 3456 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_31
timestamp 1679577901
transform 1 0 4128 0 -1 6048
box -48 -56 432 834
use sg13g2_fill_1  FILLER_5_35
timestamp 1677579658
transform 1 0 4512 0 -1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_40
timestamp 1679581782
transform 1 0 4992 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_47
timestamp 1679581782
transform 1 0 5664 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_54
timestamp 1679581782
transform 1 0 6336 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_61
timestamp 1679581782
transform 1 0 7008 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_68
timestamp 1679581782
transform 1 0 7680 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_75
timestamp 1679577901
transform 1 0 8352 0 -1 6048
box -48 -56 432 834
use sg13g2_fill_2  FILLER_5_79
timestamp 1677580104
transform 1 0 8736 0 -1 6048
box -48 -56 240 834
use sg13g2_decap_8  FILLER_5_85
timestamp 1679581782
transform 1 0 9312 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_92
timestamp 1679581782
transform 1 0 9984 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_99
timestamp 1679581782
transform 1 0 10656 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_106
timestamp 1679581782
transform 1 0 11328 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_113
timestamp 1679581782
transform 1 0 12000 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_120
timestamp 1679581782
transform 1 0 12672 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_127
timestamp 1679581782
transform 1 0 13344 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_134
timestamp 1679581782
transform 1 0 14016 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_141
timestamp 1679581782
transform 1 0 14688 0 -1 6048
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_148
timestamp 1677580104
transform 1 0 15360 0 -1 6048
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_150
timestamp 1677579658
transform 1 0 15552 0 -1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_155
timestamp 1679581782
transform 1 0 16032 0 -1 6048
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_162
timestamp 1677580104
transform 1 0 16704 0 -1 6048
box -48 -56 240 834
use sg13g2_decap_8  FILLER_5_168
timestamp 1679581782
transform 1 0 17280 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_175
timestamp 1679577901
transform 1 0 17952 0 -1 6048
box -48 -56 432 834
use sg13g2_fill_1  FILLER_5_179
timestamp 1677579658
transform 1 0 18336 0 -1 6048
box -48 -56 144 834
use sg13g2_fill_1  FILLER_5_188
timestamp 1677579658
transform 1 0 19200 0 -1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_0
timestamp 1679581782
transform 1 0 1152 0 1 6048
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_7
timestamp 1677580104
transform 1 0 1824 0 1 6048
box -48 -56 240 834
use sg13g2_decap_8  FILLER_6_13
timestamp 1679581782
transform 1 0 2400 0 1 6048
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_20
timestamp 1679577901
transform 1 0 3072 0 1 6048
box -48 -56 432 834
use sg13g2_decap_8  FILLER_6_28
timestamp 1679581782
transform 1 0 3840 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_35
timestamp 1679581782
transform 1 0 4512 0 1 6048
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_46
timestamp 1679577901
transform 1 0 5568 0 1 6048
box -48 -56 432 834
use sg13g2_fill_2  FILLER_6_50
timestamp 1677580104
transform 1 0 5952 0 1 6048
box -48 -56 240 834
use sg13g2_decap_8  FILLER_6_56
timestamp 1679581782
transform 1 0 6528 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_63
timestamp 1679581782
transform 1 0 7200 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_70
timestamp 1679581782
transform 1 0 7872 0 1 6048
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_77
timestamp 1677580104
transform 1 0 8544 0 1 6048
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_79
timestamp 1677579658
transform 1 0 8736 0 1 6048
box -48 -56 144 834
use sg13g2_fill_1  FILLER_6_84
timestamp 1677579658
transform 1 0 9216 0 1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_89
timestamp 1679581782
transform 1 0 9696 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_96
timestamp 1679581782
transform 1 0 10368 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_103
timestamp 1679581782
transform 1 0 11040 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_110
timestamp 1679581782
transform 1 0 11712 0 1 6048
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_117
timestamp 1679577901
transform 1 0 12384 0 1 6048
box -48 -56 432 834
use sg13g2_decap_8  FILLER_6_125
timestamp 1679581782
transform 1 0 13152 0 1 6048
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_132
timestamp 1679577901
transform 1 0 13824 0 1 6048
box -48 -56 432 834
use sg13g2_fill_2  FILLER_6_136
timestamp 1677580104
transform 1 0 14208 0 1 6048
box -48 -56 240 834
use sg13g2_decap_8  FILLER_6_142
timestamp 1679581782
transform 1 0 14784 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_149
timestamp 1679581782
transform 1 0 15456 0 1 6048
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_156
timestamp 1679577901
transform 1 0 16128 0 1 6048
box -48 -56 432 834
use sg13g2_fill_1  FILLER_6_160
timestamp 1677579658
transform 1 0 16512 0 1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_169
timestamp 1679581782
transform 1 0 17376 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_176
timestamp 1679581782
transform 1 0 18048 0 1 6048
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_183
timestamp 1679577901
transform 1 0 18720 0 1 6048
box -48 -56 432 834
use sg13g2_fill_1  FILLER_6_187
timestamp 1677579658
transform 1 0 19104 0 1 6048
box -48 -56 144 834
use sg13g2_fill_1  FILLER_6_192
timestamp 1677579658
transform 1 0 19584 0 1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_0
timestamp 1679581782
transform 1 0 1152 0 -1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_7_7
timestamp 1677580104
transform 1 0 1824 0 -1 7560
box -48 -56 240 834
use sg13g2_decap_8  FILLER_7_13
timestamp 1679581782
transform 1 0 2400 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_20
timestamp 1679581782
transform 1 0 3072 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_27
timestamp 1679581782
transform 1 0 3744 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_4  FILLER_7_34
timestamp 1679577901
transform 1 0 4416 0 -1 7560
box -48 -56 432 834
use sg13g2_decap_8  FILLER_7_42
timestamp 1679581782
transform 1 0 5184 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_49
timestamp 1679581782
transform 1 0 5856 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_56
timestamp 1679581782
transform 1 0 6528 0 -1 7560
box -48 -56 720 834
use sg13g2_fill_1  FILLER_7_63
timestamp 1677579658
transform 1 0 7200 0 -1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_72
timestamp 1679581782
transform 1 0 8064 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_79
timestamp 1679581782
transform 1 0 8736 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_86
timestamp 1679581782
transform 1 0 9408 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_93
timestamp 1679581782
transform 1 0 10080 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_100
timestamp 1679581782
transform 1 0 10752 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_107
timestamp 1679581782
transform 1 0 11424 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_114
timestamp 1679581782
transform 1 0 12096 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_121
timestamp 1679581782
transform 1 0 12768 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_128
timestamp 1679581782
transform 1 0 13440 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_135
timestamp 1679581782
transform 1 0 14112 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_4  FILLER_7_142
timestamp 1679577901
transform 1 0 14784 0 -1 7560
box -48 -56 432 834
use sg13g2_decap_8  FILLER_7_150
timestamp 1679581782
transform 1 0 15552 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_157
timestamp 1679581782
transform 1 0 16224 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_164
timestamp 1679581782
transform 1 0 16896 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_171
timestamp 1679581782
transform 1 0 17568 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_178
timestamp 1679581782
transform 1 0 18240 0 -1 7560
box -48 -56 720 834
use sg13g2_fill_1  FILLER_7_185
timestamp 1677579658
transform 1 0 18912 0 -1 7560
box -48 -56 144 834
use sg13g2_fill_2  FILLER_7_198
timestamp 1677580104
transform 1 0 20160 0 -1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_200
timestamp 1677579658
transform 1 0 20352 0 -1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_0
timestamp 1679581782
transform 1 0 1152 0 1 7560
box -48 -56 720 834
use sg13g2_fill_1  FILLER_8_7
timestamp 1677579658
transform 1 0 1824 0 1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_12
timestamp 1679581782
transform 1 0 2304 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_19
timestamp 1679581782
transform 1 0 2976 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_26
timestamp 1679581782
transform 1 0 3648 0 1 7560
box -48 -56 720 834
use sg13g2_fill_1  FILLER_8_33
timestamp 1677579658
transform 1 0 4320 0 1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_38
timestamp 1679581782
transform 1 0 4800 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_45
timestamp 1679581782
transform 1 0 5472 0 1 7560
box -48 -56 720 834
use sg13g2_decap_4  FILLER_8_52
timestamp 1679577901
transform 1 0 6144 0 1 7560
box -48 -56 432 834
use sg13g2_fill_2  FILLER_8_56
timestamp 1677580104
transform 1 0 6528 0 1 7560
box -48 -56 240 834
use sg13g2_decap_4  FILLER_8_62
timestamp 1679577901
transform 1 0 7104 0 1 7560
box -48 -56 432 834
use sg13g2_fill_1  FILLER_8_66
timestamp 1677579658
transform 1 0 7488 0 1 7560
box -48 -56 144 834
use sg13g2_decap_4  FILLER_8_71
timestamp 1679577901
transform 1 0 7968 0 1 7560
box -48 -56 432 834
use sg13g2_fill_2  FILLER_8_79
timestamp 1677580104
transform 1 0 8736 0 1 7560
box -48 -56 240 834
use sg13g2_decap_4  FILLER_8_85
timestamp 1679577901
transform 1 0 9312 0 1 7560
box -48 -56 432 834
use sg13g2_fill_2  FILLER_8_89
timestamp 1677580104
transform 1 0 9696 0 1 7560
box -48 -56 240 834
use sg13g2_decap_8  FILLER_8_95
timestamp 1679581782
transform 1 0 10272 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_102
timestamp 1679581782
transform 1 0 10944 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_109
timestamp 1679581782
transform 1 0 11616 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_116
timestamp 1679581782
transform 1 0 12288 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_123
timestamp 1679581782
transform 1 0 12960 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_130
timestamp 1679581782
transform 1 0 13632 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_137
timestamp 1679581782
transform 1 0 14304 0 1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_8_144
timestamp 1677580104
transform 1 0 14976 0 1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_146
timestamp 1677579658
transform 1 0 15168 0 1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_155
timestamp 1679581782
transform 1 0 16032 0 1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_8_162
timestamp 1677580104
transform 1 0 16704 0 1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_164
timestamp 1677579658
transform 1 0 16896 0 1 7560
box -48 -56 144 834
use sg13g2_decap_4  FILLER_8_169
timestamp 1679577901
transform 1 0 17376 0 1 7560
box -48 -56 432 834
use sg13g2_fill_1  FILLER_8_173
timestamp 1677579658
transform 1 0 17760 0 1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_178
timestamp 1679581782
transform 1 0 18240 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_185
timestamp 1679581782
transform 1 0 18912 0 1 7560
box -48 -56 720 834
use sg13g2_fill_1  FILLER_8_192
timestamp 1677579658
transform 1 0 19584 0 1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_0
timestamp 1679581782
transform 1 0 1152 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_11
timestamp 1679581782
transform 1 0 2208 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_18
timestamp 1679581782
transform 1 0 2880 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_25
timestamp 1679581782
transform 1 0 3552 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_32
timestamp 1679581782
transform 1 0 4224 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_39
timestamp 1679581782
transform 1 0 4896 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_46
timestamp 1679581782
transform 1 0 5568 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_53
timestamp 1679581782
transform 1 0 6240 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_60
timestamp 1679581782
transform 1 0 6912 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_67
timestamp 1679581782
transform 1 0 7584 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_4  FILLER_9_74
timestamp 1679577901
transform 1 0 8256 0 -1 9072
box -48 -56 432 834
use sg13g2_fill_1  FILLER_9_78
timestamp 1677579658
transform 1 0 8640 0 -1 9072
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_83
timestamp 1679581782
transform 1 0 9120 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_90
timestamp 1679581782
transform 1 0 9792 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_97
timestamp 1679581782
transform 1 0 10464 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_104
timestamp 1679581782
transform 1 0 11136 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_111
timestamp 1679581782
transform 1 0 11808 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_4  FILLER_9_118
timestamp 1679577901
transform 1 0 12480 0 -1 9072
box -48 -56 432 834
use sg13g2_fill_1  FILLER_9_122
timestamp 1677579658
transform 1 0 12864 0 -1 9072
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_135
timestamp 1679581782
transform 1 0 14112 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_4  FILLER_9_142
timestamp 1679577901
transform 1 0 14784 0 -1 9072
box -48 -56 432 834
use sg13g2_fill_2  FILLER_9_146
timestamp 1677580104
transform 1 0 15168 0 -1 9072
box -48 -56 240 834
use sg13g2_decap_8  FILLER_9_152
timestamp 1679581782
transform 1 0 15744 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_159
timestamp 1679581782
transform 1 0 16416 0 -1 9072
box -48 -56 720 834
use sg13g2_fill_1  FILLER_9_166
timestamp 1677579658
transform 1 0 17088 0 -1 9072
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_171
timestamp 1679581782
transform 1 0 17568 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_178
timestamp 1679581782
transform 1 0 18240 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_0
timestamp 1679581782
transform 1 0 1152 0 1 9072
box -48 -56 720 834
use sg13g2_decap_4  FILLER_10_7
timestamp 1679577901
transform 1 0 1824 0 1 9072
box -48 -56 432 834
use sg13g2_fill_1  FILLER_10_11
timestamp 1677579658
transform 1 0 2208 0 1 9072
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_16
timestamp 1679581782
transform 1 0 2688 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_23
timestamp 1679581782
transform 1 0 3360 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_30
timestamp 1679581782
transform 1 0 4032 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_37
timestamp 1679581782
transform 1 0 4704 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_44
timestamp 1679581782
transform 1 0 5376 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_51
timestamp 1679581782
transform 1 0 6048 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_58
timestamp 1679581782
transform 1 0 6720 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_65
timestamp 1679581782
transform 1 0 7392 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_72
timestamp 1679581782
transform 1 0 8064 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_79
timestamp 1679581782
transform 1 0 8736 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_86
timestamp 1679581782
transform 1 0 9408 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_93
timestamp 1679581782
transform 1 0 10080 0 1 9072
box -48 -56 720 834
use sg13g2_fill_1  FILLER_10_100
timestamp 1677579658
transform 1 0 10752 0 1 9072
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_109
timestamp 1679581782
transform 1 0 11616 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_116
timestamp 1679581782
transform 1 0 12288 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_123
timestamp 1679581782
transform 1 0 12960 0 1 9072
box -48 -56 720 834
use sg13g2_fill_1  FILLER_10_130
timestamp 1677579658
transform 1 0 13632 0 1 9072
box -48 -56 144 834
use sg13g2_fill_2  FILLER_10_139
timestamp 1677580104
transform 1 0 14496 0 1 9072
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_141
timestamp 1677579658
transform 1 0 14688 0 1 9072
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_146
timestamp 1679581782
transform 1 0 15168 0 1 9072
box -48 -56 720 834
use sg13g2_decap_4  FILLER_10_153
timestamp 1679577901
transform 1 0 15840 0 1 9072
box -48 -56 432 834
use sg13g2_fill_1  FILLER_10_157
timestamp 1677579658
transform 1 0 16224 0 1 9072
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_162
timestamp 1679581782
transform 1 0 16704 0 1 9072
box -48 -56 720 834
use sg13g2_fill_1  FILLER_10_169
timestamp 1677579658
transform 1 0 17376 0 1 9072
box -48 -56 144 834
use sg13g2_fill_2  FILLER_10_174
timestamp 1677580104
transform 1 0 17856 0 1 9072
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_196
timestamp 1677579658
transform 1 0 19968 0 1 9072
box -48 -56 144 834
use sg13g2_decap_4  FILLER_11_4
timestamp 1679577901
transform 1 0 1536 0 -1 10584
box -48 -56 432 834
use sg13g2_fill_1  FILLER_11_8
timestamp 1677579658
transform 1 0 1920 0 -1 10584
box -48 -56 144 834
use sg13g2_decap_4  FILLER_11_13
timestamp 1679577901
transform 1 0 2400 0 -1 10584
box -48 -56 432 834
use sg13g2_fill_2  FILLER_11_17
timestamp 1677580104
transform 1 0 2784 0 -1 10584
box -48 -56 240 834
use sg13g2_decap_4  FILLER_11_23
timestamp 1679577901
transform 1 0 3360 0 -1 10584
box -48 -56 432 834
use sg13g2_fill_2  FILLER_11_27
timestamp 1677580104
transform 1 0 3744 0 -1 10584
box -48 -56 240 834
use sg13g2_decap_4  FILLER_11_33
timestamp 1679577901
transform 1 0 4320 0 -1 10584
box -48 -56 432 834
use sg13g2_fill_2  FILLER_11_37
timestamp 1677580104
transform 1 0 4704 0 -1 10584
box -48 -56 240 834
use sg13g2_decap_4  FILLER_11_43
timestamp 1679577901
transform 1 0 5280 0 -1 10584
box -48 -56 432 834
use sg13g2_fill_2  FILLER_11_47
timestamp 1677580104
transform 1 0 5664 0 -1 10584
box -48 -56 240 834
use sg13g2_decap_4  FILLER_11_53
timestamp 1679577901
transform 1 0 6240 0 -1 10584
box -48 -56 432 834
use sg13g2_fill_2  FILLER_11_57
timestamp 1677580104
transform 1 0 6624 0 -1 10584
box -48 -56 240 834
use sg13g2_decap_4  FILLER_11_63
timestamp 1679577901
transform 1 0 7200 0 -1 10584
box -48 -56 432 834
use sg13g2_fill_2  FILLER_11_67
timestamp 1677580104
transform 1 0 7584 0 -1 10584
box -48 -56 240 834
use sg13g2_decap_4  FILLER_11_73
timestamp 1679577901
transform 1 0 8160 0 -1 10584
box -48 -56 432 834
use sg13g2_fill_2  FILLER_11_77
timestamp 1677580104
transform 1 0 8544 0 -1 10584
box -48 -56 240 834
use sg13g2_decap_4  FILLER_11_83
timestamp 1679577901
transform 1 0 9120 0 -1 10584
box -48 -56 432 834
use sg13g2_fill_2  FILLER_11_87
timestamp 1677580104
transform 1 0 9504 0 -1 10584
box -48 -56 240 834
use sg13g2_decap_4  FILLER_11_93
timestamp 1679577901
transform 1 0 10080 0 -1 10584
box -48 -56 432 834
use sg13g2_fill_2  FILLER_11_97
timestamp 1677580104
transform 1 0 10464 0 -1 10584
box -48 -56 240 834
use sg13g2_decap_4  FILLER_11_103
timestamp 1679577901
transform 1 0 11040 0 -1 10584
box -48 -56 432 834
use sg13g2_fill_2  FILLER_11_107
timestamp 1677580104
transform 1 0 11424 0 -1 10584
box -48 -56 240 834
use sg13g2_decap_4  FILLER_11_113
timestamp 1679577901
transform 1 0 12000 0 -1 10584
box -48 -56 432 834
use sg13g2_fill_2  FILLER_11_117
timestamp 1677580104
transform 1 0 12384 0 -1 10584
box -48 -56 240 834
use sg13g2_decap_4  FILLER_11_123
timestamp 1679577901
transform 1 0 12960 0 -1 10584
box -48 -56 432 834
use sg13g2_fill_2  FILLER_11_127
timestamp 1677580104
transform 1 0 13344 0 -1 10584
box -48 -56 240 834
use sg13g2_decap_4  FILLER_11_133
timestamp 1679577901
transform 1 0 13920 0 -1 10584
box -48 -56 432 834
use sg13g2_fill_2  FILLER_11_137
timestamp 1677580104
transform 1 0 14304 0 -1 10584
box -48 -56 240 834
use sg13g2_decap_4  FILLER_11_143
timestamp 1679577901
transform 1 0 14880 0 -1 10584
box -48 -56 432 834
use sg13g2_fill_2  FILLER_11_147
timestamp 1677580104
transform 1 0 15264 0 -1 10584
box -48 -56 240 834
use sg13g2_decap_4  FILLER_11_153
timestamp 1679577901
transform 1 0 15840 0 -1 10584
box -48 -56 432 834
use sg13g2_fill_2  FILLER_11_157
timestamp 1677580104
transform 1 0 16224 0 -1 10584
box -48 -56 240 834
use sg13g2_decap_4  FILLER_11_163
timestamp 1679577901
transform 1 0 16800 0 -1 10584
box -48 -56 432 834
use sg13g2_fill_2  FILLER_11_167
timestamp 1677580104
transform 1 0 17184 0 -1 10584
box -48 -56 240 834
use sg13g2_fill_2  FILLER_11_173
timestamp 1677580104
transform 1 0 17760 0 -1 10584
box -48 -56 240 834
use sg13g2_fill_2  FILLER_11_183
timestamp 1677580104
transform 1 0 18720 0 -1 10584
box -48 -56 240 834
use sg13g2_buf_1  output1
timestamp 1676381911
transform 1 0 18912 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output2
timestamp 1676381911
transform 1 0 20064 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output3
timestamp 1676381911
transform 1 0 18624 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output4
timestamp 1676381911
transform 1 0 20064 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output5
timestamp 1676381911
transform 1 0 19296 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output6
timestamp 1676381911
transform 1 0 20064 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output7
timestamp 1676381911
transform 1 0 19680 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output8
timestamp 1676381911
transform 1 0 20064 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output9
timestamp 1676381911
transform 1 0 19680 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  output10
timestamp 1676381911
transform 1 0 19008 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  output11
timestamp 1676381911
transform 1 0 20064 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  output12
timestamp 1676381911
transform 1 0 18528 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output13
timestamp 1676381911
transform 1 0 20064 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  output14
timestamp 1676381911
transform 1 0 19680 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  output15
timestamp 1676381911
transform 1 0 20064 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output16
timestamp 1676381911
transform 1 0 19680 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output17
timestamp 1676381911
transform 1 0 20064 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output18
timestamp 1676381911
transform 1 0 20064 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output19
timestamp 1676381911
transform 1 0 19680 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output20
timestamp 1676381911
transform 1 0 18912 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output21
timestamp 1676381911
transform 1 0 18816 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output22
timestamp 1676381911
transform 1 0 17952 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output23
timestamp 1676381911
transform 1 0 18144 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output24
timestamp 1676381911
transform 1 0 18432 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output25
timestamp 1676381911
transform 1 0 18912 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output26
timestamp 1676381911
transform 1 0 19296 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output27
timestamp 1676381911
transform 1 0 19680 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output28
timestamp 1676381911
transform 1 0 20064 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output29
timestamp 1676381911
transform 1 0 18912 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output30
timestamp 1676381911
transform 1 0 20064 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output31
timestamp 1676381911
transform 1 0 19680 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output32
timestamp 1676381911
transform 1 0 19008 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output33
timestamp 1676381911
transform -1 0 2400 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output34
timestamp 1676381911
transform -1 0 12000 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output35
timestamp 1676381911
transform -1 0 12960 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output36
timestamp 1676381911
transform -1 0 13920 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output37
timestamp 1676381911
transform -1 0 14880 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output38
timestamp 1676381911
transform -1 0 15840 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output39
timestamp 1676381911
transform -1 0 16800 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output40
timestamp 1676381911
transform -1 0 17760 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output41
timestamp 1676381911
transform -1 0 18720 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output42
timestamp 1676381911
transform -1 0 19680 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output43
timestamp 1676381911
transform 1 0 18048 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output44
timestamp 1676381911
transform -1 0 3360 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output45
timestamp 1676381911
transform -1 0 4320 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output46
timestamp 1676381911
transform -1 0 5280 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output47
timestamp 1676381911
transform -1 0 6240 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output48
timestamp 1676381911
transform -1 0 7200 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output49
timestamp 1676381911
transform -1 0 8160 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output50
timestamp 1676381911
transform -1 0 9120 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output51
timestamp 1676381911
transform -1 0 10080 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output52
timestamp 1676381911
transform -1 0 11040 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output53
timestamp 1676381911
transform 1 0 8160 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output54
timestamp 1676381911
transform -1 0 9312 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output55
timestamp 1676381911
transform 1 0 8544 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output56
timestamp 1676381911
transform -1 0 9696 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output57
timestamp 1676381911
transform 1 0 8928 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output58
timestamp 1676381911
transform -1 0 10080 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output59
timestamp 1676381911
transform 1 0 9312 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output60
timestamp 1676381911
transform -1 0 10464 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output61
timestamp 1676381911
transform 1 0 9696 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output62
timestamp 1676381911
transform -1 0 10848 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output63
timestamp 1676381911
transform 1 0 10080 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output64
timestamp 1676381911
transform -1 0 11232 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output65
timestamp 1676381911
transform 1 0 10464 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output66
timestamp 1676381911
transform 1 0 10848 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output67
timestamp 1676381911
transform 1 0 11232 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output68
timestamp 1676381911
transform -1 0 12000 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output69
timestamp 1676381911
transform -1 0 12768 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output70
timestamp 1676381911
transform -1 0 12384 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output71
timestamp 1676381911
transform -1 0 13152 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output72
timestamp 1676381911
transform -1 0 13536 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output73
timestamp 1676381911
transform -1 0 12960 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output74
timestamp 1676381911
transform -1 0 14880 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output75
timestamp 1676381911
transform -1 0 15840 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output76
timestamp 1676381911
transform -1 0 15264 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output77
timestamp 1676381911
transform -1 0 16224 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output78
timestamp 1676381911
transform -1 0 16608 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output79
timestamp 1676381911
transform -1 0 16992 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output80
timestamp 1676381911
transform -1 0 13920 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output81
timestamp 1676381911
transform -1 0 13344 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output82
timestamp 1676381911
transform -1 0 14304 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output83
timestamp 1676381911
transform -1 0 13728 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output84
timestamp 1676381911
transform -1 0 14688 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output85
timestamp 1676381911
transform -1 0 14112 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output86
timestamp 1676381911
transform -1 0 15072 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output87
timestamp 1676381911
transform -1 0 14496 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output88
timestamp 1676381911
transform -1 0 15456 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output89
timestamp 1676381911
transform -1 0 1536 0 -1 10584
box -48 -56 432 834
<< labels >>
flabel metal2 s 0 716 90 796 0 FreeSans 320 0 0 0 FrameData[0]
port 0 nsew signal input
flabel metal2 s 0 4076 90 4156 0 FreeSans 320 0 0 0 FrameData[10]
port 1 nsew signal input
flabel metal2 s 0 4412 90 4492 0 FreeSans 320 0 0 0 FrameData[11]
port 2 nsew signal input
flabel metal2 s 0 4748 90 4828 0 FreeSans 320 0 0 0 FrameData[12]
port 3 nsew signal input
flabel metal2 s 0 5084 90 5164 0 FreeSans 320 0 0 0 FrameData[13]
port 4 nsew signal input
flabel metal2 s 0 5420 90 5500 0 FreeSans 320 0 0 0 FrameData[14]
port 5 nsew signal input
flabel metal2 s 0 5756 90 5836 0 FreeSans 320 0 0 0 FrameData[15]
port 6 nsew signal input
flabel metal2 s 0 6092 90 6172 0 FreeSans 320 0 0 0 FrameData[16]
port 7 nsew signal input
flabel metal2 s 0 6428 90 6508 0 FreeSans 320 0 0 0 FrameData[17]
port 8 nsew signal input
flabel metal2 s 0 6764 90 6844 0 FreeSans 320 0 0 0 FrameData[18]
port 9 nsew signal input
flabel metal2 s 0 7100 90 7180 0 FreeSans 320 0 0 0 FrameData[19]
port 10 nsew signal input
flabel metal2 s 0 1052 90 1132 0 FreeSans 320 0 0 0 FrameData[1]
port 11 nsew signal input
flabel metal2 s 0 7436 90 7516 0 FreeSans 320 0 0 0 FrameData[20]
port 12 nsew signal input
flabel metal2 s 0 7772 90 7852 0 FreeSans 320 0 0 0 FrameData[21]
port 13 nsew signal input
flabel metal2 s 0 8108 90 8188 0 FreeSans 320 0 0 0 FrameData[22]
port 14 nsew signal input
flabel metal2 s 0 8444 90 8524 0 FreeSans 320 0 0 0 FrameData[23]
port 15 nsew signal input
flabel metal2 s 0 8780 90 8860 0 FreeSans 320 0 0 0 FrameData[24]
port 16 nsew signal input
flabel metal2 s 0 9116 90 9196 0 FreeSans 320 0 0 0 FrameData[25]
port 17 nsew signal input
flabel metal2 s 0 9452 90 9532 0 FreeSans 320 0 0 0 FrameData[26]
port 18 nsew signal input
flabel metal2 s 0 9788 90 9868 0 FreeSans 320 0 0 0 FrameData[27]
port 19 nsew signal input
flabel metal2 s 0 10124 90 10204 0 FreeSans 320 0 0 0 FrameData[28]
port 20 nsew signal input
flabel metal2 s 0 10460 90 10540 0 FreeSans 320 0 0 0 FrameData[29]
port 21 nsew signal input
flabel metal2 s 0 1388 90 1468 0 FreeSans 320 0 0 0 FrameData[2]
port 22 nsew signal input
flabel metal2 s 0 10796 90 10876 0 FreeSans 320 0 0 0 FrameData[30]
port 23 nsew signal input
flabel metal2 s 0 11132 90 11212 0 FreeSans 320 0 0 0 FrameData[31]
port 24 nsew signal input
flabel metal2 s 0 1724 90 1804 0 FreeSans 320 0 0 0 FrameData[3]
port 25 nsew signal input
flabel metal2 s 0 2060 90 2140 0 FreeSans 320 0 0 0 FrameData[4]
port 26 nsew signal input
flabel metal2 s 0 2396 90 2476 0 FreeSans 320 0 0 0 FrameData[5]
port 27 nsew signal input
flabel metal2 s 0 2732 90 2812 0 FreeSans 320 0 0 0 FrameData[6]
port 28 nsew signal input
flabel metal2 s 0 3068 90 3148 0 FreeSans 320 0 0 0 FrameData[7]
port 29 nsew signal input
flabel metal2 s 0 3404 90 3484 0 FreeSans 320 0 0 0 FrameData[8]
port 30 nsew signal input
flabel metal2 s 0 3740 90 3820 0 FreeSans 320 0 0 0 FrameData[9]
port 31 nsew signal input
flabel metal2 s 21510 716 21600 796 0 FreeSans 320 0 0 0 FrameData_O[0]
port 32 nsew signal output
flabel metal2 s 21510 4076 21600 4156 0 FreeSans 320 0 0 0 FrameData_O[10]
port 33 nsew signal output
flabel metal2 s 21510 4412 21600 4492 0 FreeSans 320 0 0 0 FrameData_O[11]
port 34 nsew signal output
flabel metal2 s 21510 4748 21600 4828 0 FreeSans 320 0 0 0 FrameData_O[12]
port 35 nsew signal output
flabel metal2 s 21510 5084 21600 5164 0 FreeSans 320 0 0 0 FrameData_O[13]
port 36 nsew signal output
flabel metal2 s 21510 5420 21600 5500 0 FreeSans 320 0 0 0 FrameData_O[14]
port 37 nsew signal output
flabel metal2 s 21510 5756 21600 5836 0 FreeSans 320 0 0 0 FrameData_O[15]
port 38 nsew signal output
flabel metal2 s 21510 6092 21600 6172 0 FreeSans 320 0 0 0 FrameData_O[16]
port 39 nsew signal output
flabel metal2 s 21510 6428 21600 6508 0 FreeSans 320 0 0 0 FrameData_O[17]
port 40 nsew signal output
flabel metal2 s 21510 6764 21600 6844 0 FreeSans 320 0 0 0 FrameData_O[18]
port 41 nsew signal output
flabel metal2 s 21510 7100 21600 7180 0 FreeSans 320 0 0 0 FrameData_O[19]
port 42 nsew signal output
flabel metal2 s 21510 1052 21600 1132 0 FreeSans 320 0 0 0 FrameData_O[1]
port 43 nsew signal output
flabel metal2 s 21510 7436 21600 7516 0 FreeSans 320 0 0 0 FrameData_O[20]
port 44 nsew signal output
flabel metal2 s 21510 7772 21600 7852 0 FreeSans 320 0 0 0 FrameData_O[21]
port 45 nsew signal output
flabel metal2 s 21510 8108 21600 8188 0 FreeSans 320 0 0 0 FrameData_O[22]
port 46 nsew signal output
flabel metal2 s 21510 8444 21600 8524 0 FreeSans 320 0 0 0 FrameData_O[23]
port 47 nsew signal output
flabel metal2 s 21510 8780 21600 8860 0 FreeSans 320 0 0 0 FrameData_O[24]
port 48 nsew signal output
flabel metal2 s 21510 9116 21600 9196 0 FreeSans 320 0 0 0 FrameData_O[25]
port 49 nsew signal output
flabel metal2 s 21510 9452 21600 9532 0 FreeSans 320 0 0 0 FrameData_O[26]
port 50 nsew signal output
flabel metal2 s 21510 9788 21600 9868 0 FreeSans 320 0 0 0 FrameData_O[27]
port 51 nsew signal output
flabel metal2 s 21510 10124 21600 10204 0 FreeSans 320 0 0 0 FrameData_O[28]
port 52 nsew signal output
flabel metal2 s 21510 10460 21600 10540 0 FreeSans 320 0 0 0 FrameData_O[29]
port 53 nsew signal output
flabel metal2 s 21510 1388 21600 1468 0 FreeSans 320 0 0 0 FrameData_O[2]
port 54 nsew signal output
flabel metal2 s 21510 10796 21600 10876 0 FreeSans 320 0 0 0 FrameData_O[30]
port 55 nsew signal output
flabel metal2 s 21510 11132 21600 11212 0 FreeSans 320 0 0 0 FrameData_O[31]
port 56 nsew signal output
flabel metal2 s 21510 1724 21600 1804 0 FreeSans 320 0 0 0 FrameData_O[3]
port 57 nsew signal output
flabel metal2 s 21510 2060 21600 2140 0 FreeSans 320 0 0 0 FrameData_O[4]
port 58 nsew signal output
flabel metal2 s 21510 2396 21600 2476 0 FreeSans 320 0 0 0 FrameData_O[5]
port 59 nsew signal output
flabel metal2 s 21510 2732 21600 2812 0 FreeSans 320 0 0 0 FrameData_O[6]
port 60 nsew signal output
flabel metal2 s 21510 3068 21600 3148 0 FreeSans 320 0 0 0 FrameData_O[7]
port 61 nsew signal output
flabel metal2 s 21510 3404 21600 3484 0 FreeSans 320 0 0 0 FrameData_O[8]
port 62 nsew signal output
flabel metal2 s 21510 3740 21600 3820 0 FreeSans 320 0 0 0 FrameData_O[9]
port 63 nsew signal output
flabel metal3 s 15800 0 15880 80 0 FreeSans 320 0 0 0 FrameStrobe[0]
port 64 nsew signal input
flabel metal3 s 17720 0 17800 80 0 FreeSans 320 0 0 0 FrameStrobe[10]
port 65 nsew signal input
flabel metal3 s 17912 0 17992 80 0 FreeSans 320 0 0 0 FrameStrobe[11]
port 66 nsew signal input
flabel metal3 s 18104 0 18184 80 0 FreeSans 320 0 0 0 FrameStrobe[12]
port 67 nsew signal input
flabel metal3 s 18296 0 18376 80 0 FreeSans 320 0 0 0 FrameStrobe[13]
port 68 nsew signal input
flabel metal3 s 18488 0 18568 80 0 FreeSans 320 0 0 0 FrameStrobe[14]
port 69 nsew signal input
flabel metal3 s 18680 0 18760 80 0 FreeSans 320 0 0 0 FrameStrobe[15]
port 70 nsew signal input
flabel metal3 s 18872 0 18952 80 0 FreeSans 320 0 0 0 FrameStrobe[16]
port 71 nsew signal input
flabel metal3 s 19064 0 19144 80 0 FreeSans 320 0 0 0 FrameStrobe[17]
port 72 nsew signal input
flabel metal3 s 19256 0 19336 80 0 FreeSans 320 0 0 0 FrameStrobe[18]
port 73 nsew signal input
flabel metal3 s 19448 0 19528 80 0 FreeSans 320 0 0 0 FrameStrobe[19]
port 74 nsew signal input
flabel metal3 s 15992 0 16072 80 0 FreeSans 320 0 0 0 FrameStrobe[1]
port 75 nsew signal input
flabel metal3 s 16184 0 16264 80 0 FreeSans 320 0 0 0 FrameStrobe[2]
port 76 nsew signal input
flabel metal3 s 16376 0 16456 80 0 FreeSans 320 0 0 0 FrameStrobe[3]
port 77 nsew signal input
flabel metal3 s 16568 0 16648 80 0 FreeSans 320 0 0 0 FrameStrobe[4]
port 78 nsew signal input
flabel metal3 s 16760 0 16840 80 0 FreeSans 320 0 0 0 FrameStrobe[5]
port 79 nsew signal input
flabel metal3 s 16952 0 17032 80 0 FreeSans 320 0 0 0 FrameStrobe[6]
port 80 nsew signal input
flabel metal3 s 17144 0 17224 80 0 FreeSans 320 0 0 0 FrameStrobe[7]
port 81 nsew signal input
flabel metal3 s 17336 0 17416 80 0 FreeSans 320 0 0 0 FrameStrobe[8]
port 82 nsew signal input
flabel metal3 s 17528 0 17608 80 0 FreeSans 320 0 0 0 FrameStrobe[9]
port 83 nsew signal input
flabel metal3 s 1976 12100 2056 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[0]
port 84 nsew signal output
flabel metal3 s 11576 12100 11656 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[10]
port 85 nsew signal output
flabel metal3 s 12536 12100 12616 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[11]
port 86 nsew signal output
flabel metal3 s 13496 12100 13576 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[12]
port 87 nsew signal output
flabel metal3 s 14456 12100 14536 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[13]
port 88 nsew signal output
flabel metal3 s 15416 12100 15496 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[14]
port 89 nsew signal output
flabel metal3 s 16376 12100 16456 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[15]
port 90 nsew signal output
flabel metal3 s 17336 12100 17416 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[16]
port 91 nsew signal output
flabel metal3 s 18296 12100 18376 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[17]
port 92 nsew signal output
flabel metal3 s 19256 12100 19336 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[18]
port 93 nsew signal output
flabel metal3 s 20216 12100 20296 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[19]
port 94 nsew signal output
flabel metal3 s 2936 12100 3016 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[1]
port 95 nsew signal output
flabel metal3 s 3896 12100 3976 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[2]
port 96 nsew signal output
flabel metal3 s 4856 12100 4936 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[3]
port 97 nsew signal output
flabel metal3 s 5816 12100 5896 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[4]
port 98 nsew signal output
flabel metal3 s 6776 12100 6856 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[5]
port 99 nsew signal output
flabel metal3 s 7736 12100 7816 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[6]
port 100 nsew signal output
flabel metal3 s 8696 12100 8776 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[7]
port 101 nsew signal output
flabel metal3 s 9656 12100 9736 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[8]
port 102 nsew signal output
flabel metal3 s 10616 12100 10696 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[9]
port 103 nsew signal output
flabel metal3 s 1784 0 1864 80 0 FreeSans 320 0 0 0 N1END[0]
port 104 nsew signal input
flabel metal3 s 1976 0 2056 80 0 FreeSans 320 0 0 0 N1END[1]
port 105 nsew signal input
flabel metal3 s 2168 0 2248 80 0 FreeSans 320 0 0 0 N1END[2]
port 106 nsew signal input
flabel metal3 s 2360 0 2440 80 0 FreeSans 320 0 0 0 N1END[3]
port 107 nsew signal input
flabel metal3 s 4088 0 4168 80 0 FreeSans 320 0 0 0 N2END[0]
port 108 nsew signal input
flabel metal3 s 4280 0 4360 80 0 FreeSans 320 0 0 0 N2END[1]
port 109 nsew signal input
flabel metal3 s 4472 0 4552 80 0 FreeSans 320 0 0 0 N2END[2]
port 110 nsew signal input
flabel metal3 s 4664 0 4744 80 0 FreeSans 320 0 0 0 N2END[3]
port 111 nsew signal input
flabel metal3 s 4856 0 4936 80 0 FreeSans 320 0 0 0 N2END[4]
port 112 nsew signal input
flabel metal3 s 5048 0 5128 80 0 FreeSans 320 0 0 0 N2END[5]
port 113 nsew signal input
flabel metal3 s 5240 0 5320 80 0 FreeSans 320 0 0 0 N2END[6]
port 114 nsew signal input
flabel metal3 s 5432 0 5512 80 0 FreeSans 320 0 0 0 N2END[7]
port 115 nsew signal input
flabel metal3 s 2552 0 2632 80 0 FreeSans 320 0 0 0 N2MID[0]
port 116 nsew signal input
flabel metal3 s 2744 0 2824 80 0 FreeSans 320 0 0 0 N2MID[1]
port 117 nsew signal input
flabel metal3 s 2936 0 3016 80 0 FreeSans 320 0 0 0 N2MID[2]
port 118 nsew signal input
flabel metal3 s 3128 0 3208 80 0 FreeSans 320 0 0 0 N2MID[3]
port 119 nsew signal input
flabel metal3 s 3320 0 3400 80 0 FreeSans 320 0 0 0 N2MID[4]
port 120 nsew signal input
flabel metal3 s 3512 0 3592 80 0 FreeSans 320 0 0 0 N2MID[5]
port 121 nsew signal input
flabel metal3 s 3704 0 3784 80 0 FreeSans 320 0 0 0 N2MID[6]
port 122 nsew signal input
flabel metal3 s 3896 0 3976 80 0 FreeSans 320 0 0 0 N2MID[7]
port 123 nsew signal input
flabel metal3 s 5624 0 5704 80 0 FreeSans 320 0 0 0 N4END[0]
port 124 nsew signal input
flabel metal3 s 7544 0 7624 80 0 FreeSans 320 0 0 0 N4END[10]
port 125 nsew signal input
flabel metal3 s 7736 0 7816 80 0 FreeSans 320 0 0 0 N4END[11]
port 126 nsew signal input
flabel metal3 s 7928 0 8008 80 0 FreeSans 320 0 0 0 N4END[12]
port 127 nsew signal input
flabel metal3 s 8120 0 8200 80 0 FreeSans 320 0 0 0 N4END[13]
port 128 nsew signal input
flabel metal3 s 8312 0 8392 80 0 FreeSans 320 0 0 0 N4END[14]
port 129 nsew signal input
flabel metal3 s 8504 0 8584 80 0 FreeSans 320 0 0 0 N4END[15]
port 130 nsew signal input
flabel metal3 s 5816 0 5896 80 0 FreeSans 320 0 0 0 N4END[1]
port 131 nsew signal input
flabel metal3 s 6008 0 6088 80 0 FreeSans 320 0 0 0 N4END[2]
port 132 nsew signal input
flabel metal3 s 6200 0 6280 80 0 FreeSans 320 0 0 0 N4END[3]
port 133 nsew signal input
flabel metal3 s 6392 0 6472 80 0 FreeSans 320 0 0 0 N4END[4]
port 134 nsew signal input
flabel metal3 s 6584 0 6664 80 0 FreeSans 320 0 0 0 N4END[5]
port 135 nsew signal input
flabel metal3 s 6776 0 6856 80 0 FreeSans 320 0 0 0 N4END[6]
port 136 nsew signal input
flabel metal3 s 6968 0 7048 80 0 FreeSans 320 0 0 0 N4END[7]
port 137 nsew signal input
flabel metal3 s 7160 0 7240 80 0 FreeSans 320 0 0 0 N4END[8]
port 138 nsew signal input
flabel metal3 s 7352 0 7432 80 0 FreeSans 320 0 0 0 N4END[9]
port 139 nsew signal input
flabel metal3 s 8696 0 8776 80 0 FreeSans 320 0 0 0 S1BEG[0]
port 140 nsew signal output
flabel metal3 s 8888 0 8968 80 0 FreeSans 320 0 0 0 S1BEG[1]
port 141 nsew signal output
flabel metal3 s 9080 0 9160 80 0 FreeSans 320 0 0 0 S1BEG[2]
port 142 nsew signal output
flabel metal3 s 9272 0 9352 80 0 FreeSans 320 0 0 0 S1BEG[3]
port 143 nsew signal output
flabel metal3 s 9464 0 9544 80 0 FreeSans 320 0 0 0 S2BEG[0]
port 144 nsew signal output
flabel metal3 s 9656 0 9736 80 0 FreeSans 320 0 0 0 S2BEG[1]
port 145 nsew signal output
flabel metal3 s 9848 0 9928 80 0 FreeSans 320 0 0 0 S2BEG[2]
port 146 nsew signal output
flabel metal3 s 10040 0 10120 80 0 FreeSans 320 0 0 0 S2BEG[3]
port 147 nsew signal output
flabel metal3 s 10232 0 10312 80 0 FreeSans 320 0 0 0 S2BEG[4]
port 148 nsew signal output
flabel metal3 s 10424 0 10504 80 0 FreeSans 320 0 0 0 S2BEG[5]
port 149 nsew signal output
flabel metal3 s 10616 0 10696 80 0 FreeSans 320 0 0 0 S2BEG[6]
port 150 nsew signal output
flabel metal3 s 10808 0 10888 80 0 FreeSans 320 0 0 0 S2BEG[7]
port 151 nsew signal output
flabel metal3 s 11000 0 11080 80 0 FreeSans 320 0 0 0 S2BEGb[0]
port 152 nsew signal output
flabel metal3 s 11192 0 11272 80 0 FreeSans 320 0 0 0 S2BEGb[1]
port 153 nsew signal output
flabel metal3 s 11384 0 11464 80 0 FreeSans 320 0 0 0 S2BEGb[2]
port 154 nsew signal output
flabel metal3 s 11576 0 11656 80 0 FreeSans 320 0 0 0 S2BEGb[3]
port 155 nsew signal output
flabel metal3 s 11768 0 11848 80 0 FreeSans 320 0 0 0 S2BEGb[4]
port 156 nsew signal output
flabel metal3 s 11960 0 12040 80 0 FreeSans 320 0 0 0 S2BEGb[5]
port 157 nsew signal output
flabel metal3 s 12152 0 12232 80 0 FreeSans 320 0 0 0 S2BEGb[6]
port 158 nsew signal output
flabel metal3 s 12344 0 12424 80 0 FreeSans 320 0 0 0 S2BEGb[7]
port 159 nsew signal output
flabel metal3 s 12536 0 12616 80 0 FreeSans 320 0 0 0 S4BEG[0]
port 160 nsew signal output
flabel metal3 s 14456 0 14536 80 0 FreeSans 320 0 0 0 S4BEG[10]
port 161 nsew signal output
flabel metal3 s 14648 0 14728 80 0 FreeSans 320 0 0 0 S4BEG[11]
port 162 nsew signal output
flabel metal3 s 14840 0 14920 80 0 FreeSans 320 0 0 0 S4BEG[12]
port 163 nsew signal output
flabel metal3 s 15032 0 15112 80 0 FreeSans 320 0 0 0 S4BEG[13]
port 164 nsew signal output
flabel metal3 s 15224 0 15304 80 0 FreeSans 320 0 0 0 S4BEG[14]
port 165 nsew signal output
flabel metal3 s 15416 0 15496 80 0 FreeSans 320 0 0 0 S4BEG[15]
port 166 nsew signal output
flabel metal3 s 12728 0 12808 80 0 FreeSans 320 0 0 0 S4BEG[1]
port 167 nsew signal output
flabel metal3 s 12920 0 13000 80 0 FreeSans 320 0 0 0 S4BEG[2]
port 168 nsew signal output
flabel metal3 s 13112 0 13192 80 0 FreeSans 320 0 0 0 S4BEG[3]
port 169 nsew signal output
flabel metal3 s 13304 0 13384 80 0 FreeSans 320 0 0 0 S4BEG[4]
port 170 nsew signal output
flabel metal3 s 13496 0 13576 80 0 FreeSans 320 0 0 0 S4BEG[5]
port 171 nsew signal output
flabel metal3 s 13688 0 13768 80 0 FreeSans 320 0 0 0 S4BEG[6]
port 172 nsew signal output
flabel metal3 s 13880 0 13960 80 0 FreeSans 320 0 0 0 S4BEG[7]
port 173 nsew signal output
flabel metal3 s 14072 0 14152 80 0 FreeSans 320 0 0 0 S4BEG[8]
port 174 nsew signal output
flabel metal3 s 14264 0 14344 80 0 FreeSans 320 0 0 0 S4BEG[9]
port 175 nsew signal output
flabel metal3 s 15608 0 15688 80 0 FreeSans 320 0 0 0 UserCLK
port 176 nsew signal input
flabel metal3 s 1016 12100 1096 12180 0 FreeSans 320 0 0 0 UserCLKo
port 177 nsew signal output
flabel metal5 s 4892 0 5332 12180 0 FreeSans 2560 90 0 0 VGND
port 178 nsew ground bidirectional
flabel metal5 s 4892 0 5332 40 0 FreeSans 320 0 0 0 VGND
port 178 nsew ground bidirectional
flabel metal5 s 4892 12140 5332 12180 0 FreeSans 320 0 0 0 VGND
port 178 nsew ground bidirectional
flabel metal5 s 20012 0 20452 12180 0 FreeSans 2560 90 0 0 VGND
port 178 nsew ground bidirectional
flabel metal5 s 20012 0 20452 40 0 FreeSans 320 0 0 0 VGND
port 178 nsew ground bidirectional
flabel metal5 s 20012 12140 20452 12180 0 FreeSans 320 0 0 0 VGND
port 178 nsew ground bidirectional
flabel metal5 s 3652 0 4092 12180 0 FreeSans 2560 90 0 0 VPWR
port 179 nsew power bidirectional
flabel metal5 s 3652 0 4092 40 0 FreeSans 320 0 0 0 VPWR
port 179 nsew power bidirectional
flabel metal5 s 3652 12140 4092 12180 0 FreeSans 320 0 0 0 VPWR
port 179 nsew power bidirectional
flabel metal5 s 18772 0 19212 12180 0 FreeSans 2560 90 0 0 VPWR
port 179 nsew power bidirectional
flabel metal5 s 18772 0 19212 40 0 FreeSans 320 0 0 0 VPWR
port 179 nsew power bidirectional
flabel metal5 s 18772 12140 19212 12180 0 FreeSans 320 0 0 0 VPWR
port 179 nsew power bidirectional
rlabel metal1 10802 10584 10802 10584 0 VGND
rlabel metal1 10800 9828 10800 9828 0 VPWR
rlabel metal3 15936 1596 15936 1596 0 FrameData[0]
rlabel metal2 752 4116 752 4116 0 FrameData[10]
rlabel metal3 18528 5040 18528 5040 0 FrameData[11]
rlabel metal2 17088 6384 17088 6384 0 FrameData[12]
rlabel metal2 512 5124 512 5124 0 FrameData[13]
rlabel via2 80 5460 80 5460 0 FrameData[14]
rlabel metal3 16704 6132 16704 6132 0 FrameData[15]
rlabel metal2 656 6132 656 6132 0 FrameData[16]
rlabel via2 80 6468 80 6468 0 FrameData[17]
rlabel via2 80 6804 80 6804 0 FrameData[18]
rlabel metal2 1040 7140 1040 7140 0 FrameData[19]
rlabel metal2 752 1092 752 1092 0 FrameData[1]
rlabel metal3 12864 6972 12864 6972 0 FrameData[20]
rlabel metal3 3072 5628 3072 5628 0 FrameData[21]
rlabel metal2 896 8148 896 8148 0 FrameData[22]
rlabel metal3 4128 6300 4128 6300 0 FrameData[23]
rlabel metal3 19872 6930 19872 6930 0 FrameData[24]
rlabel metal3 15360 8568 15360 8568 0 FrameData[25]
rlabel metal2 1208 9492 1208 9492 0 FrameData[26]
rlabel metal3 13824 8988 13824 8988 0 FrameData[27]
rlabel metal2 128 10164 128 10164 0 FrameData[28]
rlabel metal2 1344 5544 1344 5544 0 FrameData[29]
rlabel via2 80 1428 80 1428 0 FrameData[2]
rlabel metal3 8640 10206 8640 10206 0 FrameData[30]
rlabel metal2 704 11172 704 11172 0 FrameData[31]
rlabel metal2 8352 1680 8352 1680 0 FrameData[3]
rlabel metal3 7680 2310 7680 2310 0 FrameData[4]
rlabel metal2 704 2436 704 2436 0 FrameData[5]
rlabel metal2 608 2772 608 2772 0 FrameData[6]
rlabel metal3 13920 4410 13920 4410 0 FrameData[7]
rlabel metal2 1136 3444 1136 3444 0 FrameData[8]
rlabel metal3 14400 4326 14400 4326 0 FrameData[9]
rlabel metal2 21039 756 21039 756 0 FrameData_O[0]
rlabel metal2 20424 3612 20424 3612 0 FrameData_O[10]
rlabel metal2 21039 4452 21039 4452 0 FrameData_O[11]
rlabel metal2 20856 4284 20856 4284 0 FrameData_O[12]
rlabel metal2 21039 5124 21039 5124 0 FrameData_O[13]
rlabel metal2 20952 4956 20952 4956 0 FrameData_O[14]
rlabel metal2 20775 5796 20775 5796 0 FrameData_O[15]
rlabel metal2 20712 5880 20712 5880 0 FrameData_O[16]
rlabel metal2 21423 6468 21423 6468 0 FrameData_O[17]
rlabel metal2 20967 6804 20967 6804 0 FrameData_O[18]
rlabel metal2 20616 6636 20616 6636 0 FrameData_O[19]
rlabel metal2 20367 1092 20367 1092 0 FrameData_O[1]
rlabel metal2 21279 7476 21279 7476 0 FrameData_O[20]
rlabel metal2 20775 7812 20775 7812 0 FrameData_O[21]
rlabel metal2 21279 8148 21279 8148 0 FrameData_O[22]
rlabel metal2 21183 8484 21183 8484 0 FrameData_O[23]
rlabel metal2 21279 8820 21279 8820 0 FrameData_O[24]
rlabel metal2 21231 9156 21231 9156 0 FrameData_O[25]
rlabel metal2 21183 9492 21183 9492 0 FrameData_O[26]
rlabel metal2 20703 9828 20703 9828 0 FrameData_O[27]
rlabel metal2 19272 9660 19272 9660 0 FrameData_O[28]
rlabel metal2 19128 10332 19128 10332 0 FrameData_O[29]
rlabel via2 21519 1428 21519 1428 0 FrameData_O[2]
rlabel metal2 18888 9660 18888 9660 0 FrameData_O[30]
rlabel metal2 19368 8904 19368 8904 0 FrameData_O[31]
rlabel metal2 20583 1764 20583 1764 0 FrameData_O[3]
rlabel metal2 20775 2100 20775 2100 0 FrameData_O[4]
rlabel metal2 20424 2016 20424 2016 0 FrameData_O[5]
rlabel metal2 21279 2772 21279 2772 0 FrameData_O[6]
rlabel metal2 20712 2856 20712 2856 0 FrameData_O[7]
rlabel metal2 21183 3444 21183 3444 0 FrameData_O[8]
rlabel metal2 20991 3780 20991 3780 0 FrameData_O[9]
rlabel metal3 2736 4284 2736 4284 0 FrameStrobe[0]
rlabel metal2 17568 8736 17568 8736 0 FrameStrobe[10]
rlabel metal2 16176 9744 16176 9744 0 FrameStrobe[11]
rlabel metal2 16224 9828 16224 9828 0 FrameStrobe[12]
rlabel metal2 18192 8736 18192 8736 0 FrameStrobe[13]
rlabel metal3 18528 1470 18528 1470 0 FrameStrobe[14]
rlabel metal3 18768 5460 18768 5460 0 FrameStrobe[15]
rlabel metal3 18912 786 18912 786 0 FrameStrobe[16]
rlabel metal3 19104 744 19104 744 0 FrameStrobe[17]
rlabel metal3 19296 1470 19296 1470 0 FrameStrobe[18]
rlabel metal3 19488 114 19488 114 0 FrameStrobe[19]
rlabel metal3 2112 3360 2112 3360 0 FrameStrobe[1]
rlabel metal2 3648 4158 3648 4158 0 FrameStrobe[2]
rlabel metal3 16416 534 16416 534 0 FrameStrobe[3]
rlabel metal3 16608 3054 16608 3054 0 FrameStrobe[4]
rlabel metal3 16800 198 16800 198 0 FrameStrobe[5]
rlabel metal3 16992 1470 16992 1470 0 FrameStrobe[6]
rlabel metal3 16992 6594 16992 6594 0 FrameStrobe[7]
rlabel metal3 8784 1932 8784 1932 0 FrameStrobe[8]
rlabel metal3 15840 9576 15840 9576 0 FrameStrobe[9]
rlabel metal2 2040 10416 2040 10416 0 FrameStrobe_O[0]
rlabel metal2 11640 10416 11640 10416 0 FrameStrobe_O[10]
rlabel metal2 12600 10416 12600 10416 0 FrameStrobe_O[11]
rlabel metal2 13560 10416 13560 10416 0 FrameStrobe_O[12]
rlabel metal2 14520 10416 14520 10416 0 FrameStrobe_O[13]
rlabel metal2 15480 10416 15480 10416 0 FrameStrobe_O[14]
rlabel metal2 16440 10416 16440 10416 0 FrameStrobe_O[15]
rlabel metal2 17400 10416 17400 10416 0 FrameStrobe_O[16]
rlabel metal2 18360 10416 18360 10416 0 FrameStrobe_O[17]
rlabel metal2 19320 10416 19320 10416 0 FrameStrobe_O[18]
rlabel metal2 18696 9240 18696 9240 0 FrameStrobe_O[19]
rlabel metal2 3000 10416 3000 10416 0 FrameStrobe_O[1]
rlabel metal2 3960 10416 3960 10416 0 FrameStrobe_O[2]
rlabel metal2 4872 10416 4872 10416 0 FrameStrobe_O[3]
rlabel metal2 5880 10416 5880 10416 0 FrameStrobe_O[4]
rlabel metal2 6840 10416 6840 10416 0 FrameStrobe_O[5]
rlabel metal2 7800 10416 7800 10416 0 FrameStrobe_O[6]
rlabel metal2 8760 10416 8760 10416 0 FrameStrobe_O[7]
rlabel metal2 9720 10416 9720 10416 0 FrameStrobe_O[8]
rlabel metal2 10680 10416 10680 10416 0 FrameStrobe_O[9]
rlabel metal3 1824 1332 1824 1332 0 N1END[0]
rlabel metal3 2016 1290 2016 1290 0 N1END[1]
rlabel metal3 2208 2844 2208 2844 0 N1END[2]
rlabel metal3 2400 2508 2400 2508 0 N1END[3]
rlabel metal2 1920 8694 1920 8694 0 N2END[0]
rlabel metal2 4416 7980 4416 7980 0 N2END[1]
rlabel metal2 6768 7896 6768 7896 0 N2END[2]
rlabel metal2 6912 7812 6912 7812 0 N2END[3]
rlabel metal3 4896 618 4896 618 0 N2END[4]
rlabel metal3 5088 702 5088 702 0 N2END[5]
rlabel metal3 5280 702 5280 702 0 N2END[6]
rlabel metal2 7152 5124 7152 5124 0 N2END[7]
rlabel metal3 2592 114 2592 114 0 N2MID[0]
rlabel metal3 2784 2088 2784 2088 0 N2MID[1]
rlabel metal2 2544 7140 2544 7140 0 N2MID[2]
rlabel metal2 3360 6468 3360 6468 0 N2MID[3]
rlabel metal2 4032 5628 4032 5628 0 N2MID[4]
rlabel metal3 3552 1038 3552 1038 0 N2MID[5]
rlabel metal3 3744 1080 3744 1080 0 N2MID[6]
rlabel metal3 3936 1080 3936 1080 0 N2MID[7]
rlabel metal2 19584 3486 19584 3486 0 N4END[0]
rlabel metal2 9024 4032 9024 4032 0 N4END[10]
rlabel metal2 9024 4116 9024 4116 0 N4END[11]
rlabel metal2 9984 3528 9984 3528 0 N4END[12]
rlabel metal2 10176 3192 10176 3192 0 N4END[13]
rlabel metal3 8352 1080 8352 1080 0 N4END[14]
rlabel metal2 14688 3948 14688 3948 0 N4END[15]
rlabel metal2 19680 4158 19680 4158 0 N4END[1]
rlabel metal3 16704 3528 16704 3528 0 N4END[2]
rlabel metal3 6240 1710 6240 1710 0 N4END[3]
rlabel metal3 6432 954 6432 954 0 N4END[4]
rlabel metal3 6624 1122 6624 1122 0 N4END[5]
rlabel metal3 6816 1164 6816 1164 0 N4END[6]
rlabel metal3 7008 1668 7008 1668 0 N4END[7]
rlabel metal3 7200 240 7200 240 0 N4END[8]
rlabel metal3 7392 2172 7392 2172 0 N4END[9]
rlabel metal3 8736 870 8736 870 0 S1BEG[0]
rlabel metal3 8928 1248 8928 1248 0 S1BEG[1]
rlabel metal3 9120 870 9120 870 0 S1BEG[2]
rlabel metal3 9312 1248 9312 1248 0 S1BEG[3]
rlabel metal3 9504 870 9504 870 0 S2BEG[0]
rlabel metal3 9696 1248 9696 1248 0 S2BEG[1]
rlabel metal3 9888 870 9888 870 0 S2BEG[2]
rlabel metal3 10080 1248 10080 1248 0 S2BEG[3]
rlabel metal3 10272 870 10272 870 0 S2BEG[4]
rlabel metal3 10464 1248 10464 1248 0 S2BEG[5]
rlabel metal3 10656 870 10656 870 0 S2BEG[6]
rlabel metal3 10848 1248 10848 1248 0 S2BEG[7]
rlabel metal3 11040 870 11040 870 0 S2BEGb[0]
rlabel metal3 11232 870 11232 870 0 S2BEGb[1]
rlabel metal3 11424 912 11424 912 0 S2BEGb[2]
rlabel metal3 11616 870 11616 870 0 S2BEGb[3]
rlabel metal3 11808 912 11808 912 0 S2BEGb[4]
rlabel metal3 12000 870 12000 870 0 S2BEGb[5]
rlabel metal3 12192 870 12192 870 0 S2BEGb[6]
rlabel metal3 12384 828 12384 828 0 S2BEGb[7]
rlabel metal3 12576 1248 12576 1248 0 S4BEG[0]
rlabel metal3 14496 1248 14496 1248 0 S4BEG[10]
rlabel metal3 14688 912 14688 912 0 S4BEG[11]
rlabel metal3 14880 1248 14880 1248 0 S4BEG[12]
rlabel metal3 15072 828 15072 828 0 S4BEG[13]
rlabel metal3 15264 786 15264 786 0 S4BEG[14]
rlabel metal3 15456 912 15456 912 0 S4BEG[15]
rlabel metal3 12768 912 12768 912 0 S4BEG[1]
rlabel metal3 12960 240 12960 240 0 S4BEG[2]
rlabel metal3 13152 828 13152 828 0 S4BEG[3]
rlabel metal3 13344 1248 13344 1248 0 S4BEG[4]
rlabel metal3 13536 828 13536 828 0 S4BEG[5]
rlabel metal3 13728 1248 13728 1248 0 S4BEG[6]
rlabel metal3 13920 786 13920 786 0 S4BEG[7]
rlabel metal3 14112 1248 14112 1248 0 S4BEG[8]
rlabel metal3 14304 450 14304 450 0 S4BEG[9]
rlabel metal3 2640 336 2640 336 0 UserCLK
rlabel metal2 1128 10416 1128 10416 0 UserCLKo
rlabel metal2 19008 1974 19008 1974 0 net1
rlabel metal2 19104 7098 19104 7098 0 net10
rlabel metal2 20064 6468 20064 6468 0 net11
rlabel metal2 18576 1932 18576 1932 0 net12
rlabel metal2 13848 6216 13848 6216 0 net13
rlabel metal2 15072 7812 15072 7812 0 net14
rlabel metal2 20088 6216 20088 6216 0 net15
rlabel metal2 17184 8694 17184 8694 0 net16
rlabel metal2 20328 7140 20328 7140 0 net17
rlabel metal2 15720 8148 15720 8148 0 net18
rlabel metal2 19704 8904 19704 8904 0 net19
rlabel metal3 20160 3906 20160 3906 0 net2
rlabel metal2 14232 8652 14232 8652 0 net20
rlabel metal2 14472 8904 14472 8904 0 net21
rlabel metal2 2712 5628 2712 5628 0 net22
rlabel metal2 18240 1890 18240 1890 0 net23
rlabel metal4 16176 9492 16176 9492 0 net24
rlabel metal2 19056 8652 19056 8652 0 net25
rlabel metal2 19440 1932 19440 1932 0 net26
rlabel metal2 19776 2226 19776 2226 0 net27
rlabel metal2 20400 1932 20400 1932 0 net28
rlabel metal2 19152 3444 19152 3444 0 net29
rlabel via1 18744 4956 18744 4956 0 net3
rlabel metal2 19968 2646 19968 2646 0 net30
rlabel metal2 19776 3402 19776 3402 0 net31
rlabel metal2 18960 4116 18960 4116 0 net32
rlabel metal2 1992 8148 1992 8148 0 net33
rlabel metal2 13032 8904 13032 8904 0 net34
rlabel metal2 13848 9576 13848 9576 0 net35
rlabel metal2 13800 9660 13800 9660 0 net36
rlabel metal2 14808 9660 14808 9660 0 net37
rlabel metal2 15576 8904 15576 8904 0 net38
rlabel metal2 15528 7140 15528 7140 0 net39
rlabel metal2 20160 4158 20160 4158 0 net4
rlabel metal2 16440 8148 16440 8148 0 net40
rlabel metal2 17640 9660 17640 9660 0 net41
rlabel metal2 18024 9240 18024 9240 0 net42
rlabel metal2 18144 9534 18144 9534 0 net43
rlabel metal3 3264 8400 3264 8400 0 net44
rlabel metal2 4056 4284 4056 4284 0 net45
rlabel metal2 5208 6468 5208 6468 0 net46
rlabel metal2 5352 7140 5352 7140 0 net47
rlabel metal2 6936 8148 6936 8148 0 net48
rlabel metal2 8232 8148 8232 8148 0 net49
rlabel metal2 19392 5670 19392 5670 0 net5
rlabel metal2 8088 8064 8088 8064 0 net50
rlabel metal2 9528 8904 9528 8904 0 net51
rlabel metal2 10920 9660 10920 9660 0 net52
rlabel metal2 6744 4704 6744 4704 0 net53
rlabel metal2 2568 5460 2568 5460 0 net54
rlabel metal3 8064 2184 8064 2184 0 net55
rlabel metal4 9360 2604 9360 2604 0 net56
rlabel metal2 8520 7140 8520 7140 0 net57
rlabel metal2 9024 6888 9024 6888 0 net58
rlabel metal2 8640 2016 8640 2016 0 net59
rlabel metal2 20016 4956 20016 4956 0 net6
rlabel metal2 10368 2646 10368 2646 0 net60
rlabel metal2 8880 5964 8880 5964 0 net61
rlabel metal3 10752 4620 10752 4620 0 net62
rlabel metal2 9408 1848 9408 1848 0 net63
rlabel metal2 11136 2730 11136 2730 0 net64
rlabel metal2 9960 4704 9960 4704 0 net65
rlabel metal2 9960 4788 9960 4788 0 net66
rlabel metal2 11256 1932 11256 1932 0 net67
rlabel metal2 11664 1932 11664 1932 0 net68
rlabel metal2 12096 2016 12096 2016 0 net69
rlabel metal2 19632 5628 19632 5628 0 net7
rlabel metal2 12192 1932 12192 1932 0 net70
rlabel metal2 13104 1932 13104 1932 0 net71
rlabel metal2 2232 8652 2232 8652 0 net72
rlabel metal2 12864 2646 12864 2646 0 net73
rlabel metal2 14784 2562 14784 2562 0 net74
rlabel metal2 15768 1932 15768 1932 0 net75
rlabel metal2 15552 2688 15552 2688 0 net76
rlabel metal2 16752 2016 16752 2016 0 net77
rlabel metal2 18192 2016 18192 2016 0 net78
rlabel metal2 17184 1932 17184 1932 0 net79
rlabel metal2 20160 5670 20160 5670 0 net8
rlabel metal2 13944 3948 13944 3948 0 net80
rlabel metal2 13320 3948 13320 3948 0 net81
rlabel metal4 13296 2604 13296 2604 0 net82
rlabel metal3 13632 3234 13632 3234 0 net83
rlabel metal2 14640 1932 14640 1932 0 net84
rlabel metal3 14016 3318 14016 3318 0 net85
rlabel metal2 15408 1848 15408 1848 0 net86
rlabel metal2 14952 3192 14952 3192 0 net87
rlabel metal2 15504 1932 15504 1932 0 net88
rlabel metal2 1896 9660 1896 9660 0 net89
rlabel metal3 19776 7140 19776 7140 0 net9
<< properties >>
string FIXED_BBOX 0 0 21600 12180
<< end >>
