magic
tech sky130A
magscale 1 2
timestamp 1740383514
<< viali >>
rect 1593 8585 1627 8619
rect 3525 8585 3559 8619
rect 3893 8585 3927 8619
rect 4445 8585 4479 8619
rect 5457 8585 5491 8619
rect 5733 8585 5767 8619
rect 6101 8585 6135 8619
rect 6561 8585 6595 8619
rect 6929 8585 6963 8619
rect 7113 8585 7147 8619
rect 7481 8585 7515 8619
rect 8309 8585 8343 8619
rect 8585 8585 8619 8619
rect 9137 8585 9171 8619
rect 10517 8585 10551 8619
rect 11805 8585 11839 8619
rect 13093 8585 13127 8619
rect 15209 8585 15243 8619
rect 15577 8585 15611 8619
rect 16313 8585 16347 8619
rect 18061 8585 18095 8619
rect 18337 8585 18371 8619
rect 20637 8585 20671 8619
rect 23857 8585 23891 8619
rect 24777 8585 24811 8619
rect 25237 8585 25271 8619
rect 27813 8585 27847 8619
rect 32781 8585 32815 8619
rect 33517 8585 33551 8619
rect 34805 8585 34839 8619
rect 35173 8585 35207 8619
rect 36645 8585 36679 8619
rect 37749 8585 37783 8619
rect 38485 8585 38519 8619
rect 14749 8517 14783 8551
rect 16681 8517 16715 8551
rect 19717 8517 19751 8551
rect 24009 8517 24043 8551
rect 24225 8517 24259 8551
rect 24685 8517 24719 8551
rect 28641 8517 28675 8551
rect 29729 8517 29763 8551
rect 29929 8517 29963 8551
rect 30481 8517 30515 8551
rect 30665 8517 30699 8551
rect 28411 8483 28445 8517
rect 1409 8449 1443 8483
rect 1685 8449 1719 8483
rect 1869 8449 1903 8483
rect 1961 8449 1995 8483
rect 2145 8449 2179 8483
rect 2513 8449 2547 8483
rect 3249 8449 3283 8483
rect 3341 8449 3375 8483
rect 4997 8449 5031 8483
rect 5457 8449 5491 8483
rect 5549 8449 5583 8483
rect 5917 8449 5951 8483
rect 6745 8449 6779 8483
rect 6837 8449 6871 8483
rect 7297 8449 7331 8483
rect 7389 8449 7423 8483
rect 7665 8449 7699 8483
rect 7757 8449 7791 8483
rect 8125 8449 8159 8483
rect 8769 8449 8803 8483
rect 9321 8449 9355 8483
rect 10333 8449 10367 8483
rect 11621 8449 11655 8483
rect 11989 8449 12023 8483
rect 12173 8449 12207 8483
rect 12265 8449 12299 8483
rect 12357 8449 12391 8483
rect 12817 8449 12851 8483
rect 12909 8449 12943 8483
rect 13553 8449 13587 8483
rect 13645 8449 13679 8483
rect 15025 8449 15059 8483
rect 15393 8449 15427 8483
rect 15761 8449 15795 8483
rect 16129 8449 16163 8483
rect 16497 8449 16531 8483
rect 17601 8449 17635 8483
rect 17877 8449 17911 8483
rect 18245 8449 18279 8483
rect 18521 8449 18555 8483
rect 18981 8449 19015 8483
rect 19073 8449 19107 8483
rect 19441 8449 19475 8483
rect 21465 8449 21499 8483
rect 23029 8449 23063 8483
rect 25451 8449 25485 8483
rect 25605 8449 25639 8483
rect 26065 8449 26099 8483
rect 27077 8449 27111 8483
rect 27629 8449 27663 8483
rect 28181 8449 28215 8483
rect 28917 8449 28951 8483
rect 29101 8449 29135 8483
rect 29219 8449 29253 8483
rect 30205 8449 30239 8483
rect 30757 8449 30791 8483
rect 30849 8449 30883 8483
rect 31493 8449 31527 8483
rect 31585 8449 31619 8483
rect 31677 8449 31711 8483
rect 32137 8449 32171 8483
rect 32603 8449 32637 8483
rect 32965 8449 32999 8483
rect 33333 8449 33367 8483
rect 33977 8449 34011 8483
rect 34345 8449 34379 8483
rect 34989 8449 35023 8483
rect 35357 8449 35391 8483
rect 35725 8449 35759 8483
rect 36093 8449 36127 8483
rect 36461 8449 36495 8483
rect 36829 8449 36863 8483
rect 37289 8449 37323 8483
rect 37933 8449 37967 8483
rect 38025 8449 38059 8483
rect 38669 8449 38703 8483
rect 38853 8449 38887 8483
rect 39221 8449 39255 8483
rect 2237 8381 2271 8415
rect 4537 8381 4571 8415
rect 4721 8381 4755 8415
rect 9413 8381 9447 8415
rect 9965 8381 9999 8415
rect 11345 8381 11379 8415
rect 14105 8381 14139 8415
rect 17233 8381 17267 8415
rect 17417 8381 17451 8415
rect 18705 8381 18739 8415
rect 18797 8381 18831 8415
rect 20361 8381 20395 8415
rect 21281 8381 21315 8415
rect 22017 8381 22051 8415
rect 22661 8381 22695 8415
rect 22753 8381 22787 8415
rect 23765 8381 23799 8415
rect 24593 8381 24627 8415
rect 25789 8381 25823 8415
rect 31125 8381 31159 8415
rect 31309 8381 31343 8415
rect 2053 8313 2087 8347
rect 4077 8313 4111 8347
rect 5181 8313 5215 8347
rect 7941 8313 7975 8347
rect 13369 8313 13403 8347
rect 13829 8313 13863 8347
rect 15945 8313 15979 8347
rect 17785 8313 17819 8347
rect 18889 8313 18923 8347
rect 19625 8313 19659 8347
rect 22845 8313 22879 8347
rect 23305 8313 23339 8347
rect 23489 8313 23523 8347
rect 25145 8313 25179 8347
rect 27997 8313 28031 8347
rect 28273 8313 28307 8347
rect 29377 8313 29411 8347
rect 31033 8313 31067 8347
rect 33149 8313 33183 8347
rect 34161 8313 34195 8347
rect 35541 8313 35575 8347
rect 35909 8313 35943 8347
rect 38209 8313 38243 8347
rect 39037 8313 39071 8347
rect 39405 8313 39439 8347
rect 1777 8245 1811 8279
rect 10701 8245 10735 8279
rect 12633 8245 12667 8279
rect 14841 8245 14875 8279
rect 21649 8245 21683 8279
rect 23213 8245 23247 8279
rect 24041 8245 24075 8279
rect 26801 8245 26835 8279
rect 28457 8245 28491 8279
rect 28733 8245 28767 8279
rect 29561 8245 29595 8279
rect 29745 8245 29779 8279
rect 30021 8245 30055 8279
rect 31861 8245 31895 8279
rect 32321 8245 32355 8279
rect 33793 8245 33827 8279
rect 36277 8245 36311 8279
rect 37473 8245 37507 8279
rect 3525 8041 3559 8075
rect 4813 8041 4847 8075
rect 6929 8041 6963 8075
rect 7849 8041 7883 8075
rect 12173 8041 12207 8075
rect 16681 8041 16715 8075
rect 18245 8041 18279 8075
rect 29561 8041 29595 8075
rect 30205 8041 30239 8075
rect 33885 8041 33919 8075
rect 34805 8041 34839 8075
rect 35725 8041 35759 8075
rect 36277 8041 36311 8075
rect 36829 8041 36863 8075
rect 38025 8041 38059 8075
rect 38669 8041 38703 8075
rect 6745 7973 6779 8007
rect 14289 7973 14323 8007
rect 16497 7973 16531 8007
rect 28457 7973 28491 8007
rect 28733 7973 28767 8007
rect 29193 7973 29227 8007
rect 2329 7905 2363 7939
rect 5457 7905 5491 7939
rect 5733 7905 5767 7939
rect 7481 7905 7515 7939
rect 8769 7905 8803 7939
rect 8953 7905 8987 7939
rect 19901 7905 19935 7939
rect 28089 7905 28123 7939
rect 30481 7905 30515 7939
rect 32321 7905 32355 7939
rect 32965 7905 32999 7939
rect 33149 7905 33183 7939
rect 1409 7837 1443 7871
rect 1685 7837 1719 7871
rect 2605 7837 2639 7871
rect 3341 7837 3375 7871
rect 3801 7837 3835 7871
rect 4077 7837 4111 7871
rect 5273 7837 5307 7871
rect 6009 7837 6043 7871
rect 7297 7837 7331 7871
rect 8033 7837 8067 7871
rect 8125 7837 8159 7871
rect 8309 7837 8343 7871
rect 8401 7837 8435 7871
rect 8539 7837 8573 7871
rect 9220 7837 9254 7871
rect 10517 7837 10551 7871
rect 10701 7837 10735 7871
rect 10793 7837 10827 7871
rect 12357 7837 12391 7871
rect 12624 7837 12658 7871
rect 14105 7837 14139 7871
rect 14289 7837 14323 7871
rect 14381 7837 14415 7871
rect 14565 7837 14599 7871
rect 14657 7837 14691 7871
rect 14749 7837 14783 7871
rect 15117 7837 15151 7871
rect 17794 7837 17828 7871
rect 18061 7837 18095 7871
rect 18429 7837 18463 7871
rect 18613 7837 18647 7871
rect 18705 7837 18739 7871
rect 18889 7837 18923 7871
rect 20453 7837 20487 7871
rect 24041 7837 24075 7871
rect 27905 7837 27939 7871
rect 28365 7837 28399 7871
rect 28641 7837 28675 7871
rect 28917 7837 28951 7871
rect 29009 7837 29043 7871
rect 29745 7837 29779 7871
rect 30021 7837 30055 7871
rect 30297 7837 30331 7871
rect 30389 7837 30423 7871
rect 32229 7837 32263 7871
rect 33057 7837 33091 7871
rect 33333 7837 33367 7871
rect 33793 7837 33827 7871
rect 34069 7837 34103 7871
rect 34989 7837 35023 7871
rect 35909 7837 35943 7871
rect 36461 7837 36495 7871
rect 37013 7837 37047 7871
rect 37841 7837 37875 7871
rect 38485 7837 38519 7871
rect 38853 7837 38887 7871
rect 39221 7837 39255 7871
rect 11060 7769 11094 7803
rect 15025 7769 15059 7803
rect 15362 7769 15396 7803
rect 19073 7769 19107 7803
rect 20177 7769 20211 7803
rect 20361 7769 20395 7803
rect 23774 7769 23808 7803
rect 24501 7769 24535 7803
rect 26249 7769 26283 7803
rect 26341 7769 26375 7803
rect 30113 7769 30147 7803
rect 30748 7769 30782 7803
rect 4905 7701 4939 7735
rect 5365 7701 5399 7735
rect 7389 7701 7423 7735
rect 10333 7701 10367 7735
rect 10701 7701 10735 7735
rect 13737 7701 13771 7735
rect 19257 7701 19291 7735
rect 19993 7701 20027 7735
rect 22661 7701 22695 7735
rect 28181 7701 28215 7735
rect 29929 7701 29963 7735
rect 31861 7701 31895 7735
rect 32045 7701 32079 7735
rect 33517 7701 33551 7735
rect 33609 7701 33643 7735
rect 39037 7701 39071 7735
rect 39405 7701 39439 7735
rect 2513 7497 2547 7531
rect 2697 7497 2731 7531
rect 3157 7497 3191 7531
rect 4997 7497 5031 7531
rect 5181 7497 5215 7531
rect 6653 7497 6687 7531
rect 16891 7497 16925 7531
rect 18521 7497 18555 7531
rect 20177 7497 20211 7531
rect 21649 7497 21683 7531
rect 22477 7497 22511 7531
rect 24961 7497 24995 7531
rect 26801 7497 26835 7531
rect 27353 7497 27387 7531
rect 30021 7497 30055 7531
rect 31953 7497 31987 7531
rect 32965 7497 32999 7531
rect 34345 7497 34379 7531
rect 37473 7497 37507 7531
rect 38301 7497 38335 7531
rect 38669 7497 38703 7531
rect 39037 7497 39071 7531
rect 7021 7429 7055 7463
rect 8217 7429 8251 7463
rect 8554 7429 8588 7463
rect 13102 7429 13136 7463
rect 14942 7429 14976 7463
rect 16681 7429 16715 7463
rect 20536 7429 20570 7463
rect 23866 7429 23900 7463
rect 26249 7429 26283 7463
rect 27445 7429 27479 7463
rect 28264 7429 28298 7463
rect 30205 7429 30239 7463
rect 30840 7429 30874 7463
rect 1409 7361 1443 7395
rect 2329 7361 2363 7395
rect 2881 7361 2915 7395
rect 2973 7361 3007 7395
rect 3617 7361 3651 7395
rect 4721 7361 4755 7395
rect 4813 7361 4847 7395
rect 5917 7361 5951 7395
rect 6837 7361 6871 7395
rect 7113 7361 7147 7395
rect 7757 7361 7791 7395
rect 8033 7361 8067 7395
rect 8309 7361 8343 7395
rect 9965 7361 9999 7395
rect 10232 7361 10266 7395
rect 11713 7361 11747 7395
rect 13461 7361 13495 7395
rect 15209 7361 15243 7395
rect 15393 7361 15427 7395
rect 15669 7361 15703 7395
rect 15853 7361 15887 7395
rect 16129 7361 16163 7395
rect 16497 7361 16531 7395
rect 17141 7361 17175 7395
rect 17397 7361 17431 7395
rect 18804 7361 18838 7395
rect 19064 7361 19098 7395
rect 20269 7361 20303 7395
rect 21833 7361 21867 7395
rect 24133 7361 24167 7395
rect 24409 7361 24443 7395
rect 26525 7361 26559 7395
rect 26617 7361 26651 7395
rect 27997 7361 28031 7395
rect 29653 7361 29687 7395
rect 30113 7361 30147 7395
rect 30573 7361 30607 7395
rect 32597 7361 32631 7395
rect 32873 7361 32907 7395
rect 33149 7361 33183 7395
rect 33425 7361 33459 7395
rect 33701 7361 33735 7395
rect 33977 7361 34011 7395
rect 34253 7361 34287 7395
rect 34529 7361 34563 7395
rect 37657 7361 37691 7395
rect 37749 7361 37783 7395
rect 38117 7361 38151 7395
rect 38485 7361 38519 7395
rect 38853 7361 38887 7395
rect 39221 7361 39255 7395
rect 1685 7293 1719 7327
rect 3341 7293 3375 7327
rect 6193 7293 6227 7327
rect 7849 7293 7883 7327
rect 11529 7293 11563 7327
rect 13369 7293 13403 7327
rect 15485 7293 15519 7327
rect 27537 7293 27571 7327
rect 29745 7293 29779 7327
rect 32137 7293 32171 7327
rect 7297 7225 7331 7259
rect 7573 7225 7607 7259
rect 13645 7225 13679 7259
rect 15577 7225 15611 7259
rect 16313 7225 16347 7259
rect 17049 7225 17083 7259
rect 29377 7225 29411 7259
rect 32229 7225 32263 7259
rect 33241 7225 33275 7259
rect 33517 7225 33551 7259
rect 37933 7225 37967 7259
rect 4353 7157 4387 7191
rect 4721 7157 4755 7191
rect 9689 7157 9723 7191
rect 11345 7157 11379 7191
rect 11897 7157 11931 7191
rect 11989 7157 12023 7191
rect 13829 7157 13863 7191
rect 16037 7157 16071 7191
rect 16865 7157 16899 7191
rect 22753 7157 22787 7191
rect 24225 7157 24259 7191
rect 26341 7157 26375 7191
rect 26985 7157 27019 7191
rect 32689 7157 32723 7191
rect 33793 7157 33827 7191
rect 34069 7157 34103 7191
rect 39405 7157 39439 7191
rect 2789 6953 2823 6987
rect 7389 6953 7423 6987
rect 11069 6953 11103 6987
rect 11161 6953 11195 6987
rect 12357 6953 12391 6987
rect 18613 6953 18647 6987
rect 18889 6953 18923 6987
rect 23673 6953 23707 6987
rect 29101 6953 29135 6987
rect 34529 6953 34563 6987
rect 2421 6885 2455 6919
rect 6469 6885 6503 6919
rect 13737 6885 13771 6919
rect 18061 6885 18095 6919
rect 18153 6885 18187 6919
rect 24041 6885 24075 6919
rect 25789 6885 25823 6919
rect 26893 6885 26927 6919
rect 29377 6885 29411 6919
rect 31033 6885 31067 6919
rect 33701 6885 33735 6919
rect 38209 6885 38243 6919
rect 4445 6817 4479 6851
rect 7021 6817 7055 6851
rect 7113 6817 7147 6851
rect 11805 6817 11839 6851
rect 15577 6817 15611 6851
rect 15669 6817 15703 6851
rect 16589 6817 16623 6851
rect 17417 6817 17451 6851
rect 18245 6817 18279 6851
rect 18429 6817 18463 6851
rect 19349 6817 19383 6851
rect 20453 6817 20487 6851
rect 22385 6817 22419 6851
rect 27721 6817 27755 6851
rect 29929 6817 29963 6851
rect 30757 6817 30791 6851
rect 31401 6817 31435 6851
rect 33885 6817 33919 6851
rect 1961 6749 1995 6783
rect 2513 6749 2547 6783
rect 2605 6749 2639 6783
rect 3249 6749 3283 6783
rect 3617 6749 3651 6783
rect 4261 6749 4295 6783
rect 4353 6749 4387 6783
rect 4997 6749 5031 6783
rect 5365 6749 5399 6783
rect 5457 6749 5491 6783
rect 5733 6749 5767 6783
rect 6929 6749 6963 6783
rect 8769 6749 8803 6783
rect 8953 6749 8987 6783
rect 10425 6749 10459 6783
rect 10609 6749 10643 6783
rect 10701 6749 10735 6783
rect 10793 6749 10827 6783
rect 13737 6749 13771 6783
rect 13921 6749 13955 6783
rect 16681 6749 16715 6783
rect 17233 6749 17267 6783
rect 18142 6749 18176 6783
rect 18797 6765 18831 6799
rect 19064 6749 19098 6783
rect 19625 6749 19659 6783
rect 22201 6749 22235 6783
rect 23305 6749 23339 6783
rect 23489 6749 23523 6783
rect 23765 6749 23799 6783
rect 24225 6749 24259 6783
rect 24409 6749 24443 6783
rect 24685 6749 24719 6783
rect 25697 6749 25731 6783
rect 26525 6749 26559 6783
rect 26801 6749 26835 6783
rect 27077 6749 27111 6783
rect 27353 6749 27387 6783
rect 27629 6749 27663 6783
rect 27988 6749 28022 6783
rect 29193 6749 29227 6783
rect 29561 6749 29595 6783
rect 29837 6749 29871 6783
rect 30021 6749 30055 6783
rect 30297 6749 30331 6783
rect 30665 6749 30699 6783
rect 31493 6749 31527 6783
rect 31953 6749 31987 6783
rect 32229 6749 32263 6783
rect 32505 6749 32539 6783
rect 32689 6749 32723 6783
rect 32965 6749 32999 6783
rect 35357 6749 35391 6783
rect 36001 6749 36035 6783
rect 37933 6749 37967 6783
rect 38117 6749 38151 6783
rect 38393 6749 38427 6783
rect 38485 6749 38519 6783
rect 38853 6749 38887 6783
rect 39221 6749 39255 6783
rect 2145 6681 2179 6715
rect 8502 6681 8536 6715
rect 9198 6681 9232 6715
rect 13645 6681 13679 6715
rect 15332 6681 15366 6715
rect 1777 6613 1811 6647
rect 2237 6613 2271 6647
rect 3065 6613 3099 6647
rect 3433 6613 3467 6647
rect 3893 6613 3927 6647
rect 4813 6613 4847 6647
rect 5181 6613 5215 6647
rect 6561 6613 6595 6647
rect 7389 6613 7423 6647
rect 10333 6613 10367 6647
rect 11161 6613 11195 6647
rect 14197 6613 14231 6647
rect 16313 6613 16347 6647
rect 16865 6613 16899 6647
rect 17049 6613 17083 6647
rect 17601 6613 17635 6647
rect 17693 6613 17727 6647
rect 20361 6613 20395 6647
rect 22569 6613 22603 6647
rect 22661 6613 22695 6647
rect 23029 6613 23063 6647
rect 23121 6613 23155 6647
rect 23949 6613 23983 6647
rect 25421 6613 25455 6647
rect 25513 6613 25547 6647
rect 27169 6613 27203 6647
rect 27445 6613 27479 6647
rect 29101 6613 29135 6647
rect 29745 6613 29779 6647
rect 30113 6613 30147 6647
rect 31125 6613 31159 6647
rect 31769 6613 31803 6647
rect 32045 6613 32079 6647
rect 32321 6613 32355 6647
rect 34069 6613 34103 6647
rect 34161 6613 34195 6647
rect 35541 6613 35575 6647
rect 35817 6613 35851 6647
rect 37749 6613 37783 6647
rect 38025 6613 38059 6647
rect 38669 6613 38703 6647
rect 39037 6613 39071 6647
rect 39405 6613 39439 6647
rect 1593 6409 1627 6443
rect 2329 6409 2363 6443
rect 6009 6409 6043 6443
rect 6469 6409 6503 6443
rect 6837 6409 6871 6443
rect 7205 6409 7239 6443
rect 7573 6409 7607 6443
rect 9413 6409 9447 6443
rect 10793 6409 10827 6443
rect 26525 6409 26559 6443
rect 26801 6409 26835 6443
rect 27445 6409 27479 6443
rect 29837 6409 29871 6443
rect 31401 6409 31435 6443
rect 31677 6409 31711 6443
rect 33793 6409 33827 6443
rect 33885 6409 33919 6443
rect 36093 6409 36127 6443
rect 39405 6409 39439 6443
rect 1961 6341 1995 6375
rect 3709 6341 3743 6375
rect 8309 6341 8343 6375
rect 9505 6341 9539 6375
rect 10333 6341 10367 6375
rect 11345 6341 11379 6375
rect 16405 6341 16439 6375
rect 19533 6341 19567 6375
rect 21281 6341 21315 6375
rect 22201 6341 22235 6375
rect 36461 6341 36495 6375
rect 22431 6307 22465 6341
rect 1777 6273 1811 6307
rect 2513 6273 2547 6307
rect 3157 6273 3191 6307
rect 4261 6273 4295 6307
rect 4629 6273 4663 6307
rect 4997 6273 5031 6307
rect 6193 6273 6227 6307
rect 6653 6273 6687 6307
rect 7021 6273 7055 6307
rect 7389 6273 7423 6307
rect 7757 6273 7791 6307
rect 7849 6273 7883 6307
rect 8033 6273 8067 6307
rect 8217 6273 8251 6307
rect 8585 6273 8619 6307
rect 8677 6273 8711 6307
rect 8769 6273 8803 6307
rect 8953 6273 8987 6307
rect 9229 6273 9263 6307
rect 10149 6273 10183 6307
rect 10517 6273 10551 6307
rect 10609 6273 10643 6307
rect 11069 6273 11103 6307
rect 11161 6273 11195 6307
rect 11888 6273 11922 6307
rect 13645 6273 13679 6307
rect 15954 6273 15988 6307
rect 16313 6273 16347 6307
rect 16491 6273 16525 6307
rect 16865 6273 16899 6307
rect 17141 6273 17175 6307
rect 17693 6273 17727 6307
rect 18613 6273 18647 6307
rect 18797 6273 18831 6307
rect 19073 6273 19107 6307
rect 19441 6273 19475 6307
rect 21557 6273 21591 6307
rect 22017 6273 22051 6307
rect 22753 6273 22787 6307
rect 22937 6273 22971 6307
rect 24133 6273 24167 6307
rect 25237 6273 25271 6307
rect 25697 6273 25731 6307
rect 25973 6273 26007 6307
rect 26341 6273 26375 6307
rect 26617 6273 26651 6307
rect 26985 6273 27019 6307
rect 27629 6273 27663 6307
rect 27997 6273 28031 6307
rect 29101 6273 29135 6307
rect 30297 6273 30331 6307
rect 30665 6273 30699 6307
rect 31493 6273 31527 6307
rect 31953 6273 31987 6307
rect 32597 6273 32631 6307
rect 35265 6273 35299 6307
rect 38577 6273 38611 6307
rect 38669 6273 38703 6307
rect 39129 6273 39163 6307
rect 39221 6273 39255 6307
rect 2145 6205 2179 6239
rect 3249 6205 3283 6239
rect 3341 6205 3375 6239
rect 4721 6205 4755 6239
rect 9045 6205 9079 6239
rect 11621 6205 11655 6239
rect 14565 6205 14599 6239
rect 16221 6205 16255 6239
rect 16681 6205 16715 6239
rect 17049 6205 17083 6239
rect 17417 6205 17451 6239
rect 21925 6205 21959 6239
rect 23857 6205 23891 6239
rect 27721 6205 27755 6239
rect 28825 6205 28859 6239
rect 30389 6205 30423 6239
rect 32321 6205 32355 6239
rect 33885 6205 33919 6239
rect 33977 6205 34011 6239
rect 34989 6205 35023 6239
rect 36553 6205 36587 6239
rect 36645 6205 36679 6239
rect 3893 6137 3927 6171
rect 4445 6137 4479 6171
rect 22569 6137 22603 6171
rect 33333 6137 33367 6171
rect 36001 6137 36035 6171
rect 38393 6137 38427 6171
rect 39037 6137 39071 6171
rect 2789 6069 2823 6103
rect 4077 6069 4111 6103
rect 5733 6069 5767 6103
rect 10333 6069 10367 6103
rect 10885 6069 10919 6103
rect 11345 6069 11379 6103
rect 13001 6069 13035 6103
rect 13093 6069 13127 6103
rect 14013 6069 14047 6103
rect 14841 6069 14875 6103
rect 17325 6069 17359 6103
rect 18429 6069 18463 6103
rect 18613 6069 18647 6103
rect 18889 6069 18923 6103
rect 19257 6069 19291 6103
rect 20821 6069 20855 6103
rect 21373 6069 21407 6103
rect 22385 6069 22419 6103
rect 22937 6069 22971 6103
rect 24869 6069 24903 6103
rect 25053 6069 25087 6103
rect 25513 6069 25547 6103
rect 25789 6069 25823 6103
rect 27169 6069 27203 6103
rect 28733 6069 28767 6103
rect 30113 6069 30147 6103
rect 31769 6069 31803 6103
rect 33425 6069 33459 6103
rect 38853 6069 38887 6103
rect 2053 5865 2087 5899
rect 2605 5865 2639 5899
rect 4261 5865 4295 5899
rect 7021 5865 7055 5899
rect 7573 5865 7607 5899
rect 8125 5865 8159 5899
rect 10425 5865 10459 5899
rect 14105 5865 14139 5899
rect 15577 5865 15611 5899
rect 17325 5865 17359 5899
rect 17693 5865 17727 5899
rect 28181 5865 28215 5899
rect 30021 5865 30055 5899
rect 31217 5865 31251 5899
rect 32229 5865 32263 5899
rect 37473 5865 37507 5899
rect 37933 5865 37967 5899
rect 1777 5797 1811 5831
rect 3893 5797 3927 5831
rect 23121 5797 23155 5831
rect 24041 5797 24075 5831
rect 27077 5797 27111 5831
rect 28641 5797 28675 5831
rect 29377 5797 29411 5831
rect 38577 5797 38611 5831
rect 39405 5797 39439 5831
rect 5549 5729 5583 5763
rect 5733 5729 5767 5763
rect 8401 5729 8435 5763
rect 9045 5729 9079 5763
rect 11069 5729 11103 5763
rect 17969 5729 18003 5763
rect 19257 5729 19291 5763
rect 21281 5729 21315 5763
rect 21925 5729 21959 5763
rect 22318 5729 22352 5763
rect 24869 5729 24903 5763
rect 24961 5729 24995 5763
rect 27721 5729 27755 5763
rect 28917 5729 28951 5763
rect 34805 5729 34839 5763
rect 1961 5661 1995 5695
rect 2329 5661 2363 5695
rect 2513 5661 2547 5695
rect 3341 5661 3375 5695
rect 3617 5661 3651 5695
rect 4077 5661 4111 5695
rect 4445 5661 4479 5695
rect 4813 5661 4847 5695
rect 5273 5661 5307 5695
rect 6009 5661 6043 5695
rect 7205 5661 7239 5695
rect 7757 5661 7791 5695
rect 8309 5661 8343 5695
rect 8585 5661 8619 5695
rect 11437 5661 11471 5695
rect 11621 5661 11655 5695
rect 11713 5661 11747 5695
rect 11805 5661 11839 5695
rect 13921 5661 13955 5695
rect 15485 5661 15519 5695
rect 15853 5661 15887 5695
rect 15945 5661 15979 5695
rect 16037 5661 16071 5695
rect 16221 5661 16255 5695
rect 16313 5661 16347 5695
rect 16589 5661 16623 5695
rect 17509 5661 17543 5695
rect 18153 5661 18187 5695
rect 18797 5661 18831 5695
rect 19073 5661 19107 5695
rect 19513 5661 19547 5695
rect 21096 5661 21130 5695
rect 21189 5661 21223 5695
rect 21465 5661 21499 5695
rect 22201 5661 22235 5695
rect 22477 5661 22511 5695
rect 23397 5661 23431 5695
rect 24225 5661 24259 5695
rect 24777 5661 24811 5695
rect 26893 5637 26927 5671
rect 28365 5661 28399 5695
rect 28457 5661 28491 5695
rect 28733 5661 28767 5695
rect 29009 5661 29043 5695
rect 29745 5661 29779 5695
rect 29837 5661 29871 5695
rect 30205 5661 30239 5695
rect 30481 5661 30515 5695
rect 31777 5661 31811 5695
rect 32045 5661 32079 5695
rect 33425 5661 33459 5695
rect 35081 5661 35115 5695
rect 37657 5661 37691 5695
rect 37749 5661 37783 5695
rect 38485 5661 38519 5695
rect 38761 5661 38795 5695
rect 38853 5661 38887 5695
rect 39221 5661 39255 5695
rect 1593 5593 1627 5627
rect 8769 5593 8803 5627
rect 9290 5593 9324 5627
rect 12081 5593 12115 5627
rect 12173 5593 12207 5627
rect 15240 5593 15274 5627
rect 27537 5593 27571 5627
rect 4905 5525 4939 5559
rect 5365 5525 5399 5559
rect 6745 5525 6779 5559
rect 10517 5525 10551 5559
rect 18061 5525 18095 5559
rect 18521 5525 18555 5559
rect 18613 5525 18647 5559
rect 18889 5525 18923 5559
rect 20637 5525 20671 5559
rect 20821 5525 20855 5559
rect 23213 5525 23247 5559
rect 24409 5525 24443 5559
rect 27169 5525 27203 5559
rect 27629 5525 27663 5559
rect 29561 5525 29595 5559
rect 31953 5525 31987 5559
rect 33241 5525 33275 5559
rect 35817 5525 35851 5559
rect 38301 5525 38335 5559
rect 39037 5525 39071 5559
rect 2053 5321 2087 5355
rect 3065 5321 3099 5355
rect 6009 5321 6043 5355
rect 6929 5321 6963 5355
rect 16221 5321 16255 5355
rect 18751 5321 18785 5355
rect 21833 5321 21867 5355
rect 23489 5321 23523 5355
rect 25145 5321 25179 5355
rect 26985 5321 27019 5355
rect 29101 5321 29135 5355
rect 29193 5321 29227 5355
rect 29837 5321 29871 5355
rect 30205 5321 30239 5355
rect 31769 5321 31803 5355
rect 37289 5321 37323 5355
rect 38301 5321 38335 5355
rect 38577 5321 38611 5355
rect 39405 5321 39439 5355
rect 5181 5253 5215 5287
rect 6469 5253 6503 5287
rect 15678 5253 15712 5287
rect 18061 5253 18095 5287
rect 18153 5253 18187 5287
rect 1593 5185 1627 5219
rect 1869 5185 1903 5219
rect 2237 5185 2271 5219
rect 2605 5185 2639 5219
rect 3249 5185 3283 5219
rect 3341 5185 3375 5219
rect 3617 5185 3651 5219
rect 4537 5185 4571 5219
rect 5273 5185 5307 5219
rect 6193 5185 6227 5219
rect 6745 5185 6779 5219
rect 8134 5185 8168 5219
rect 8760 5185 8794 5219
rect 10241 5185 10275 5219
rect 10333 5185 10367 5219
rect 10425 5185 10459 5219
rect 10609 5185 10643 5219
rect 11529 5185 11563 5219
rect 11713 5185 11747 5219
rect 11805 5185 11839 5219
rect 11897 5185 11931 5219
rect 12449 5185 12483 5219
rect 15945 5185 15979 5219
rect 16037 5185 16071 5219
rect 16681 5185 16715 5219
rect 16957 5185 16991 5219
rect 18854 5185 18888 5219
rect 19165 5185 19199 5219
rect 19717 5185 19751 5219
rect 20821 5185 20855 5219
rect 22201 5185 22235 5219
rect 23029 5185 23063 5219
rect 23121 5185 23155 5219
rect 23581 5185 23615 5219
rect 23765 5185 23799 5219
rect 25789 5185 25823 5219
rect 26065 5185 26099 5219
rect 27169 5185 27203 5219
rect 28319 5185 28353 5219
rect 30941 5185 30975 5219
rect 31953 5185 31987 5219
rect 32137 5185 32171 5219
rect 32413 5185 32447 5219
rect 37473 5185 37507 5219
rect 38485 5185 38519 5219
rect 38761 5185 38795 5219
rect 38853 5185 38887 5219
rect 39221 5185 39255 5219
rect 4997 5117 5031 5151
rect 8401 5117 8435 5151
rect 8493 5117 8527 5151
rect 11345 5117 11379 5151
rect 17877 5117 17911 5151
rect 19441 5117 19475 5151
rect 20545 5117 20579 5151
rect 22293 5117 22327 5151
rect 22385 5117 22419 5151
rect 23213 5117 23247 5151
rect 23305 5117 23339 5151
rect 23673 5117 23707 5151
rect 24961 5117 24995 5151
rect 25053 5117 25087 5151
rect 27261 5117 27295 5151
rect 27445 5117 27479 5151
rect 28181 5117 28215 5151
rect 28457 5117 28491 5151
rect 29377 5117 29411 5151
rect 29469 5117 29503 5151
rect 31217 5117 31251 5151
rect 1777 5049 1811 5083
rect 2789 5049 2823 5083
rect 4353 5049 4387 5083
rect 6653 5049 6687 5083
rect 12173 5049 12207 5083
rect 17693 5049 17727 5083
rect 19349 5049 19383 5083
rect 27905 5049 27939 5083
rect 2329 4981 2363 5015
rect 4629 4981 4663 5015
rect 5641 4981 5675 5015
rect 7021 4981 7055 5015
rect 9873 4981 9907 5015
rect 9965 4981 9999 5015
rect 10701 4981 10735 5015
rect 14565 4981 14599 5015
rect 18521 4981 18555 5015
rect 20453 4981 20487 5015
rect 21557 4981 21591 5015
rect 25513 4981 25547 5015
rect 26801 4981 26835 5015
rect 33149 4981 33183 5015
rect 39037 4981 39071 5015
rect 1593 4777 1627 4811
rect 2421 4777 2455 4811
rect 3433 4777 3467 4811
rect 8125 4777 8159 4811
rect 14105 4777 14139 4811
rect 17141 4777 17175 4811
rect 18981 4777 19015 4811
rect 22753 4777 22787 4811
rect 23305 4777 23339 4811
rect 27261 4777 27295 4811
rect 29193 4777 29227 4811
rect 34713 4777 34747 4811
rect 36001 4777 36035 4811
rect 37381 4777 37415 4811
rect 38393 4777 38427 4811
rect 3801 4709 3835 4743
rect 4721 4709 4755 4743
rect 7757 4709 7791 4743
rect 11345 4709 11379 4743
rect 13001 4709 13035 4743
rect 16129 4709 16163 4743
rect 18429 4709 18463 4743
rect 20545 4709 20579 4743
rect 29745 4709 29779 4743
rect 31953 4709 31987 4743
rect 38209 4709 38243 4743
rect 39405 4709 39439 4743
rect 4353 4641 4387 4675
rect 5616 4641 5650 4675
rect 6009 4641 6043 4675
rect 6653 4641 6687 4675
rect 9045 4641 9079 4675
rect 9413 4641 9447 4675
rect 9505 4641 9539 4675
rect 13277 4641 13311 4675
rect 13921 4641 13955 4675
rect 14749 4641 14783 4675
rect 17325 4641 17359 4675
rect 19533 4641 19567 4675
rect 21097 4641 21131 4675
rect 21557 4641 21591 4675
rect 21833 4641 21867 4675
rect 21971 4641 22005 4675
rect 22109 4641 22143 4675
rect 23857 4641 23891 4675
rect 24961 4641 24995 4675
rect 27997 4641 28031 4675
rect 32597 4641 32631 4675
rect 32689 4641 32723 4675
rect 33517 4641 33551 4675
rect 38301 4641 38335 4675
rect 1501 4573 1535 4607
rect 2237 4573 2271 4607
rect 2513 4573 2547 4607
rect 2881 4573 2915 4607
rect 3249 4573 3283 4607
rect 4169 4573 4203 4607
rect 4629 4573 4663 4607
rect 5457 4573 5491 4607
rect 5733 4573 5767 4607
rect 6469 4573 6503 4607
rect 6745 4573 6779 4607
rect 7021 4573 7055 4607
rect 8401 4573 8435 4607
rect 8493 4573 8527 4607
rect 8585 4567 8619 4601
rect 8769 4573 8803 4607
rect 9229 4573 9263 4607
rect 10977 4573 11011 4607
rect 11161 4573 11195 4607
rect 11621 4573 11655 4607
rect 14289 4573 14323 4607
rect 14473 4573 14507 4607
rect 16313 4573 16347 4607
rect 16497 4573 16531 4607
rect 16589 4573 16623 4607
rect 16681 4573 16715 4607
rect 17049 4573 17083 4607
rect 17601 4573 17635 4607
rect 18613 4573 18647 4607
rect 18797 4573 18831 4607
rect 19257 4573 19291 4607
rect 19809 4573 19843 4607
rect 20821 4573 20855 4607
rect 20913 4573 20947 4607
rect 23673 4573 23707 4607
rect 24869 4573 24903 4607
rect 26249 4573 26283 4607
rect 26525 4573 26559 4607
rect 27353 4573 27387 4607
rect 27537 4573 27571 4607
rect 28273 4573 28307 4607
rect 28390 4573 28424 4607
rect 28549 4573 28583 4607
rect 30481 4573 30515 4607
rect 30757 4573 30791 4607
rect 30941 4573 30975 4607
rect 31217 4573 31251 4607
rect 32505 4573 32539 4607
rect 33425 4573 33459 4607
rect 35449 4573 35483 4607
rect 35725 4573 35759 4607
rect 35817 4573 35851 4607
rect 37565 4573 37599 4607
rect 38577 4573 38611 4607
rect 38669 4573 38703 4607
rect 39129 4573 39163 4607
rect 39221 4573 39255 4607
rect 1869 4505 1903 4539
rect 2053 4505 2087 4539
rect 4261 4505 4295 4539
rect 9772 4505 9806 4539
rect 11888 4505 11922 4539
rect 15016 4505 15050 4539
rect 16957 4505 16991 4539
rect 23765 4505 23799 4539
rect 33333 4505 33367 4539
rect 2697 4437 2731 4471
rect 3065 4437 3099 4471
rect 4813 4437 4847 4471
rect 10885 4437 10919 4471
rect 16129 4437 16163 4471
rect 18337 4437 18371 4471
rect 19441 4437 19475 4471
rect 20637 4437 20671 4471
rect 24409 4437 24443 4471
rect 24777 4437 24811 4471
rect 32137 4437 32171 4471
rect 32965 4437 32999 4471
rect 38853 4437 38887 4471
rect 39129 4437 39163 4471
rect 3801 4233 3835 4267
rect 5549 4233 5583 4267
rect 6653 4233 6687 4267
rect 6745 4233 6779 4267
rect 7113 4233 7147 4267
rect 8861 4233 8895 4267
rect 9413 4233 9447 4267
rect 10885 4233 10919 4267
rect 12909 4233 12943 4267
rect 13277 4233 13311 4267
rect 13461 4233 13495 4267
rect 14013 4233 14047 4267
rect 15577 4233 15611 4267
rect 15669 4233 15703 4267
rect 18889 4233 18923 4267
rect 22201 4233 22235 4267
rect 22293 4233 22327 4267
rect 23213 4233 23247 4267
rect 25329 4233 25363 4267
rect 25421 4233 25455 4267
rect 30849 4233 30883 4267
rect 10977 4165 11011 4199
rect 11774 4165 11808 4199
rect 13921 4165 13955 4199
rect 14473 4165 14507 4199
rect 18429 4165 18463 4199
rect 20821 4165 20855 4199
rect 27997 4165 28031 4199
rect 28917 4165 28951 4199
rect 36369 4165 36403 4199
rect 2513 4097 2547 4131
rect 3065 4097 3099 4131
rect 4169 4097 4203 4131
rect 5181 4097 5215 4131
rect 5273 4097 5307 4131
rect 5733 4097 5767 4131
rect 5825 4097 5859 4131
rect 6653 4097 6687 4131
rect 8217 4097 8251 4131
rect 8493 4097 8527 4131
rect 8677 4097 8711 4131
rect 8769 4097 8803 4131
rect 8944 4095 8978 4129
rect 9045 4097 9079 4131
rect 9229 4097 9263 4131
rect 9321 4097 9355 4131
rect 9505 4095 9539 4129
rect 10333 4097 10367 4131
rect 10517 4097 10551 4131
rect 11529 4097 11563 4131
rect 13093 4097 13127 4131
rect 13277 4097 13311 4131
rect 13553 4097 13587 4131
rect 14933 4097 14967 4131
rect 15393 4097 15427 4131
rect 15853 4097 15887 4131
rect 16037 4097 16071 4131
rect 16221 4097 16255 4131
rect 16313 4097 16347 4131
rect 23305 4097 23339 4131
rect 23949 4097 23983 4131
rect 24409 4097 24443 4131
rect 27537 4097 27571 4131
rect 28089 4097 28123 4131
rect 29929 4097 29963 4131
rect 30205 4097 30239 4131
rect 30389 4097 30423 4131
rect 30665 4097 30699 4131
rect 32413 4097 32447 4131
rect 32965 4097 32999 4131
rect 34897 4097 34931 4131
rect 35173 4097 35207 4131
rect 36461 4097 36495 4131
rect 37565 4097 37599 4131
rect 38853 4097 38887 4131
rect 39221 4097 39255 4131
rect 1409 4029 1443 4063
rect 1685 4029 1719 4063
rect 2789 4029 2823 4063
rect 3893 4029 3927 4063
rect 6561 4029 6595 4063
rect 10241 4029 10275 4063
rect 10793 4029 10827 4063
rect 13829 4029 13863 4063
rect 14749 4029 14783 4063
rect 15209 4029 15243 4063
rect 16129 4029 16163 4063
rect 18981 4029 19015 4063
rect 19073 4029 19107 4063
rect 20913 4029 20947 4063
rect 21005 4029 21039 4063
rect 22477 4029 22511 4063
rect 23121 4029 23155 4063
rect 25237 4029 25271 4063
rect 25329 4029 25363 4063
rect 28273 4029 28307 4063
rect 28457 4029 28491 4063
rect 36553 4029 36587 4063
rect 4905 3961 4939 3995
rect 4997 3961 5031 3995
rect 6009 3961 6043 3995
rect 8033 3961 8067 3995
rect 8585 3961 8619 3995
rect 9137 3961 9171 3995
rect 14381 3961 14415 3995
rect 17141 3961 17175 3995
rect 20453 3961 20487 3995
rect 21833 3961 21867 3995
rect 27629 3961 27663 3995
rect 28549 3961 28583 3995
rect 32229 3961 32263 3995
rect 35909 3961 35943 3995
rect 37381 3961 37415 3995
rect 39405 3961 39439 3995
rect 2697 3893 2731 3927
rect 5457 3893 5491 3927
rect 9597 3893 9631 3927
rect 10425 3893 10459 3927
rect 11345 3893 11379 3927
rect 14565 3893 14599 3927
rect 15117 3893 15151 3927
rect 16497 3893 16531 3927
rect 18521 3893 18555 3927
rect 23673 3893 23707 3927
rect 23765 3893 23799 3927
rect 24225 3893 24259 3927
rect 25789 3893 25823 3927
rect 27353 3893 27387 3927
rect 29745 3893 29779 3927
rect 30113 3893 30147 3927
rect 30573 3893 30607 3927
rect 32781 3893 32815 3927
rect 36001 3893 36035 3927
rect 39037 3893 39071 3927
rect 2789 3689 2823 3723
rect 5457 3689 5491 3723
rect 5733 3689 5767 3723
rect 8953 3689 8987 3723
rect 11437 3689 11471 3723
rect 11621 3689 11655 3723
rect 13369 3689 13403 3723
rect 14473 3689 14507 3723
rect 21005 3689 21039 3723
rect 23121 3689 23155 3723
rect 24225 3689 24259 3723
rect 26341 3689 26375 3723
rect 28917 3689 28951 3723
rect 29193 3689 29227 3723
rect 1961 3621 1995 3655
rect 2513 3621 2547 3655
rect 3433 3621 3467 3655
rect 8677 3621 8711 3655
rect 14197 3621 14231 3655
rect 18337 3621 18371 3655
rect 24501 3621 24535 3655
rect 24777 3621 24811 3655
rect 30941 3621 30975 3655
rect 39405 3621 39439 3655
rect 4445 3553 4479 3587
rect 7573 3553 7607 3587
rect 7665 3553 7699 3587
rect 9505 3553 9539 3587
rect 10425 3553 10459 3587
rect 11897 3553 11931 3587
rect 15025 3553 15059 3587
rect 25329 3553 25363 3587
rect 25789 3553 25823 3587
rect 25881 3553 25915 3587
rect 26801 3553 26835 3587
rect 27905 3553 27939 3587
rect 30573 3553 30607 3587
rect 1501 3485 1535 3519
rect 1777 3485 1811 3519
rect 2053 3485 2087 3519
rect 2329 3485 2363 3519
rect 2605 3485 2639 3519
rect 2881 3485 2915 3519
rect 3617 3485 3651 3519
rect 4721 3485 4755 3519
rect 5549 3485 5583 3519
rect 7389 3485 7423 3519
rect 7941 3485 7975 3519
rect 9321 3485 9355 3519
rect 10701 3485 10735 3519
rect 11529 3485 11563 3519
rect 11713 3485 11747 3519
rect 13553 3485 13587 3519
rect 13921 3485 13955 3519
rect 14381 3485 14415 3519
rect 14841 3485 14875 3519
rect 15301 3485 15335 3519
rect 15853 3485 15887 3519
rect 16957 3485 16991 3519
rect 17969 3485 18003 3519
rect 18245 3485 18279 3519
rect 18521 3485 18555 3519
rect 18797 3485 18831 3519
rect 19073 3485 19107 3519
rect 20821 3485 20855 3519
rect 21281 3485 21315 3519
rect 21465 3485 21499 3519
rect 22109 3485 22143 3519
rect 22385 3485 22419 3519
rect 23213 3485 23247 3519
rect 23489 3485 23523 3519
rect 24685 3485 24719 3519
rect 25145 3485 25179 3519
rect 25973 3485 26007 3519
rect 27077 3485 27111 3519
rect 28181 3485 28215 3519
rect 29009 3485 29043 3519
rect 30297 3485 30331 3519
rect 31677 3485 31711 3519
rect 31953 3485 31987 3519
rect 32689 3485 32723 3519
rect 35909 3485 35943 3519
rect 38853 3485 38887 3519
rect 39221 3485 39255 3519
rect 1685 3417 1719 3451
rect 3893 3417 3927 3451
rect 10149 3417 10183 3451
rect 12164 3417 12198 3451
rect 25237 3417 25271 3451
rect 2237 3349 2271 3383
rect 3065 3349 3099 3383
rect 3433 3349 3467 3383
rect 3985 3349 4019 3383
rect 9413 3349 9447 3383
rect 10241 3349 10275 3383
rect 13277 3349 13311 3383
rect 13737 3349 13771 3383
rect 14933 3349 14967 3383
rect 15485 3349 15519 3383
rect 15669 3349 15703 3383
rect 17141 3349 17175 3383
rect 17233 3349 17267 3383
rect 18613 3349 18647 3383
rect 18889 3349 18923 3383
rect 21097 3349 21131 3383
rect 21649 3349 21683 3383
rect 27813 3349 27847 3383
rect 29561 3349 29595 3383
rect 32505 3349 32539 3383
rect 35817 3349 35851 3383
rect 39037 3349 39071 3383
rect 1685 3145 1719 3179
rect 6745 3145 6779 3179
rect 9965 3145 9999 3179
rect 11529 3145 11563 3179
rect 13921 3145 13955 3179
rect 17049 3145 17083 3179
rect 17141 3145 17175 3179
rect 24133 3145 24167 3179
rect 25237 3145 25271 3179
rect 25329 3145 25363 3179
rect 29929 3145 29963 3179
rect 30297 3145 30331 3179
rect 30389 3145 30423 3179
rect 34897 3145 34931 3179
rect 34989 3145 35023 3179
rect 36829 3145 36863 3179
rect 39405 3145 39439 3179
rect 4721 3077 4755 3111
rect 29837 3077 29871 3111
rect 1501 3009 1535 3043
rect 1777 3009 1811 3043
rect 2053 3009 2087 3043
rect 2329 3009 2363 3043
rect 2605 3009 2639 3043
rect 2881 3009 2915 3043
rect 5273 3009 5307 3043
rect 6837 3009 6871 3043
rect 7573 3009 7607 3043
rect 7849 3009 7883 3043
rect 8953 3009 8987 3043
rect 9781 3009 9815 3043
rect 10333 3009 10367 3043
rect 10609 3009 10643 3043
rect 11713 3009 11747 3043
rect 11805 3009 11839 3043
rect 12081 3009 12115 3043
rect 12909 3009 12943 3043
rect 13185 3009 13219 3043
rect 14289 3009 14323 3043
rect 15393 3009 15427 3043
rect 17785 3009 17819 3043
rect 18797 3009 18831 3043
rect 19809 3009 19843 3043
rect 20453 3009 20487 3043
rect 20729 3009 20763 3043
rect 22293 3009 22327 3043
rect 23489 3009 23523 3043
rect 23949 3009 23983 3043
rect 24501 3009 24535 3043
rect 25513 3009 25547 3043
rect 25789 3009 25823 3043
rect 26801 3009 26835 3043
rect 27721 3009 27755 3043
rect 28089 3009 28123 3043
rect 30573 3009 30607 3043
rect 31585 3009 31619 3043
rect 32413 3009 32447 3043
rect 33425 3009 33459 3043
rect 33701 3009 33735 3043
rect 35357 3009 35391 3043
rect 36645 3009 36679 3043
rect 38761 3009 38795 3043
rect 38853 3009 38887 3043
rect 39221 3009 39255 3043
rect 4997 2941 5031 2975
rect 6929 2941 6963 2975
rect 8677 2941 8711 2975
rect 14013 2941 14047 2975
rect 15117 2941 15151 2975
rect 16957 2941 16991 2975
rect 17049 2941 17083 2975
rect 17601 2941 17635 2975
rect 18521 2941 18555 2975
rect 18659 2941 18693 2975
rect 19533 2941 19567 2975
rect 22017 2941 22051 2975
rect 23581 2941 23615 2975
rect 23673 2941 23707 2975
rect 24225 2941 24259 2975
rect 27997 2941 28031 2975
rect 29653 2941 29687 2975
rect 31861 2941 31895 2975
rect 32137 2941 32171 2975
rect 34989 2941 35023 2975
rect 35081 2941 35115 2975
rect 1961 2873 1995 2907
rect 2237 2873 2271 2907
rect 2513 2873 2547 2907
rect 4905 2873 4939 2907
rect 6009 2873 6043 2907
rect 16129 2873 16163 2907
rect 18245 2873 18279 2907
rect 23029 2873 23063 2907
rect 28273 2873 28307 2907
rect 30849 2873 30883 2907
rect 34529 2873 34563 2907
rect 35541 2873 35575 2907
rect 2789 2805 2823 2839
rect 3065 2805 3099 2839
rect 6377 2805 6411 2839
rect 8585 2805 8619 2839
rect 9689 2805 9723 2839
rect 11345 2805 11379 2839
rect 12817 2805 12851 2839
rect 15025 2805 15059 2839
rect 17509 2805 17543 2839
rect 19441 2805 19475 2839
rect 21465 2805 21499 2839
rect 23121 2805 23155 2839
rect 25973 2805 26007 2839
rect 26617 2805 26651 2839
rect 26985 2805 27019 2839
rect 33149 2805 33183 2839
rect 34437 2805 34471 2839
rect 38577 2805 38611 2839
rect 39037 2805 39071 2839
rect 1961 2601 1995 2635
rect 6009 2601 6043 2635
rect 10517 2601 10551 2635
rect 11529 2601 11563 2635
rect 13185 2601 13219 2635
rect 14565 2601 14599 2635
rect 15761 2601 15795 2635
rect 17969 2601 18003 2635
rect 21557 2601 21591 2635
rect 22937 2601 22971 2635
rect 26985 2601 27019 2635
rect 30849 2601 30883 2635
rect 32505 2601 32539 2635
rect 33701 2601 33735 2635
rect 10977 2533 11011 2567
rect 20177 2533 20211 2567
rect 39405 2533 39439 2567
rect 9045 2465 9079 2499
rect 12081 2465 12115 2499
rect 13737 2465 13771 2499
rect 15209 2465 15243 2499
rect 15301 2465 15335 2499
rect 18981 2465 19015 2499
rect 21005 2465 21039 2499
rect 27445 2465 27479 2499
rect 27537 2465 27571 2499
rect 33057 2465 33091 2499
rect 1869 2397 1903 2431
rect 2237 2397 2271 2431
rect 2605 2397 2639 2431
rect 2697 2397 2731 2431
rect 2973 2397 3007 2431
rect 4077 2397 4111 2431
rect 4813 2397 4847 2431
rect 5917 2397 5951 2431
rect 6193 2397 6227 2431
rect 7021 2397 7055 2431
rect 8033 2397 8067 2431
rect 8401 2397 8435 2431
rect 8585 2397 8619 2431
rect 10333 2397 10367 2431
rect 10701 2397 10735 2431
rect 10793 2397 10827 2431
rect 11075 2397 11109 2431
rect 11897 2397 11931 2431
rect 12633 2397 12667 2431
rect 12909 2397 12943 2431
rect 13553 2397 13587 2431
rect 14105 2397 14139 2431
rect 14749 2397 14783 2431
rect 16129 2397 16163 2431
rect 16957 2397 16991 2431
rect 17693 2397 17727 2431
rect 18705 2397 18739 2431
rect 19441 2397 19475 2431
rect 19993 2397 20027 2431
rect 21833 2397 21867 2431
rect 23121 2397 23155 2431
rect 27353 2397 27387 2431
rect 30665 2397 30699 2431
rect 31769 2397 31803 2431
rect 32873 2397 32907 2431
rect 33517 2397 33551 2431
rect 34345 2397 34379 2431
rect 37749 2397 37783 2431
rect 38117 2397 38151 2431
rect 38485 2397 38519 2431
rect 38853 2397 38887 2431
rect 39221 2397 39255 2431
rect 1501 2329 1535 2363
rect 8769 2329 8803 2363
rect 11989 2329 12023 2363
rect 13645 2329 13679 2363
rect 15393 2329 15427 2363
rect 1593 2261 1627 2295
rect 2421 2261 2455 2295
rect 2881 2261 2915 2295
rect 3157 2261 3191 2295
rect 3893 2261 3927 2295
rect 4629 2261 4663 2295
rect 5733 2261 5767 2295
rect 6837 2261 6871 2295
rect 7849 2261 7883 2295
rect 8217 2261 8251 2295
rect 9229 2261 9263 2295
rect 9321 2261 9355 2295
rect 9689 2261 9723 2295
rect 10149 2261 10183 2295
rect 11253 2261 11287 2295
rect 12449 2261 12483 2295
rect 13093 2261 13127 2295
rect 14289 2261 14323 2295
rect 15945 2261 15979 2295
rect 16773 2261 16807 2295
rect 17509 2261 17543 2295
rect 19257 2261 19291 2295
rect 21097 2261 21131 2295
rect 21189 2261 21223 2295
rect 22017 2261 22051 2295
rect 31953 2261 31987 2295
rect 32965 2261 32999 2295
rect 34253 2261 34287 2295
rect 37933 2261 37967 2295
rect 38301 2261 38335 2295
rect 38669 2261 38703 2295
rect 39037 2261 39071 2295
<< metal1 >>
rect 6638 11160 6644 11212
rect 6696 11200 6702 11212
rect 12894 11200 12900 11212
rect 6696 11172 12900 11200
rect 6696 11160 6702 11172
rect 12894 11160 12900 11172
rect 12952 11160 12958 11212
rect 17218 10820 17224 10872
rect 17276 10860 17282 10872
rect 18414 10860 18420 10872
rect 17276 10832 18420 10860
rect 17276 10820 17282 10832
rect 18414 10820 18420 10832
rect 18472 10820 18478 10872
rect 12986 10684 12992 10736
rect 13044 10724 13050 10736
rect 14550 10724 14556 10736
rect 13044 10696 14556 10724
rect 13044 10684 13050 10696
rect 14550 10684 14556 10696
rect 14608 10684 14614 10736
rect 12894 10480 12900 10532
rect 12952 10520 12958 10532
rect 20990 10520 20996 10532
rect 12952 10492 20996 10520
rect 12952 10480 12958 10492
rect 20990 10480 20996 10492
rect 21048 10480 21054 10532
rect 1486 10412 1492 10464
rect 1544 10452 1550 10464
rect 3510 10452 3516 10464
rect 1544 10424 3516 10452
rect 1544 10412 1550 10424
rect 3510 10412 3516 10424
rect 3568 10412 3574 10464
rect 23014 10452 23020 10464
rect 4632 10424 23020 10452
rect 2038 10208 2044 10260
rect 2096 10248 2102 10260
rect 4632 10248 4660 10424
rect 23014 10412 23020 10424
rect 23072 10412 23078 10464
rect 7282 10344 7288 10396
rect 7340 10384 7346 10396
rect 22370 10384 22376 10396
rect 7340 10356 22376 10384
rect 7340 10344 7346 10356
rect 22370 10344 22376 10356
rect 22428 10344 22434 10396
rect 8938 10276 8944 10328
rect 8996 10316 9002 10328
rect 17126 10316 17132 10328
rect 8996 10288 17132 10316
rect 8996 10276 9002 10288
rect 17126 10276 17132 10288
rect 17184 10276 17190 10328
rect 28902 10276 28908 10328
rect 28960 10316 28966 10328
rect 32398 10316 32404 10328
rect 28960 10288 32404 10316
rect 28960 10276 28966 10288
rect 32398 10276 32404 10288
rect 32456 10276 32462 10328
rect 2096 10220 4660 10248
rect 2096 10208 2102 10220
rect 9490 10208 9496 10260
rect 9548 10248 9554 10260
rect 17494 10248 17500 10260
rect 9548 10220 17500 10248
rect 9548 10208 9554 10220
rect 17494 10208 17500 10220
rect 17552 10208 17558 10260
rect 6454 10140 6460 10192
rect 6512 10180 6518 10192
rect 8754 10180 8760 10192
rect 6512 10152 8760 10180
rect 6512 10140 6518 10152
rect 8754 10140 8760 10152
rect 8812 10140 8818 10192
rect 12802 10140 12808 10192
rect 12860 10180 12866 10192
rect 19058 10180 19064 10192
rect 12860 10152 19064 10180
rect 12860 10140 12866 10152
rect 19058 10140 19064 10152
rect 19116 10140 19122 10192
rect 23566 10140 23572 10192
rect 23624 10180 23630 10192
rect 30466 10180 30472 10192
rect 23624 10152 30472 10180
rect 23624 10140 23630 10152
rect 30466 10140 30472 10152
rect 30524 10140 30530 10192
rect 7006 10072 7012 10124
rect 7064 10112 7070 10124
rect 7064 10084 9720 10112
rect 7064 10072 7070 10084
rect 7834 10004 7840 10056
rect 7892 10044 7898 10056
rect 9582 10044 9588 10056
rect 7892 10016 9588 10044
rect 7892 10004 7898 10016
rect 9582 10004 9588 10016
rect 9640 10004 9646 10056
rect 9692 10044 9720 10084
rect 10226 10072 10232 10124
rect 10284 10112 10290 10124
rect 10284 10084 17172 10112
rect 10284 10072 10290 10084
rect 9692 10016 17080 10044
rect 3694 9936 3700 9988
rect 3752 9976 3758 9988
rect 6546 9976 6552 9988
rect 3752 9948 6552 9976
rect 3752 9936 3758 9948
rect 6546 9936 6552 9948
rect 6604 9936 6610 9988
rect 8386 9936 8392 9988
rect 8444 9976 8450 9988
rect 13722 9976 13728 9988
rect 8444 9948 13728 9976
rect 8444 9936 8450 9948
rect 13722 9936 13728 9948
rect 13780 9936 13786 9988
rect 6086 9868 6092 9920
rect 6144 9908 6150 9920
rect 11790 9908 11796 9920
rect 6144 9880 11796 9908
rect 6144 9868 6150 9880
rect 11790 9868 11796 9880
rect 11848 9868 11854 9920
rect 11882 9868 11888 9920
rect 11940 9908 11946 9920
rect 12618 9908 12624 9920
rect 11940 9880 12624 9908
rect 11940 9868 11946 9880
rect 12618 9868 12624 9880
rect 12676 9868 12682 9920
rect 17052 9908 17080 10016
rect 17144 9976 17172 10084
rect 19150 10072 19156 10124
rect 19208 10112 19214 10124
rect 20898 10112 20904 10124
rect 19208 10084 20904 10112
rect 19208 10072 19214 10084
rect 20898 10072 20904 10084
rect 20956 10072 20962 10124
rect 20990 10072 20996 10124
rect 21048 10112 21054 10124
rect 30742 10112 30748 10124
rect 21048 10084 30748 10112
rect 21048 10072 21054 10084
rect 30742 10072 30748 10084
rect 30800 10072 30806 10124
rect 17494 10004 17500 10056
rect 17552 10044 17558 10056
rect 26602 10044 26608 10056
rect 17552 10016 26608 10044
rect 17552 10004 17558 10016
rect 26602 10004 26608 10016
rect 26660 10004 26666 10056
rect 27982 9976 27988 9988
rect 17144 9948 27988 9976
rect 27982 9936 27988 9948
rect 28040 9936 28046 9988
rect 26786 9908 26792 9920
rect 17052 9880 26792 9908
rect 26786 9868 26792 9880
rect 26844 9868 26850 9920
rect 35618 9908 35624 9920
rect 31726 9880 35624 9908
rect 6178 9800 6184 9852
rect 6236 9840 6242 9852
rect 7926 9840 7932 9852
rect 6236 9812 7932 9840
rect 6236 9800 6242 9812
rect 7926 9800 7932 9812
rect 7984 9800 7990 9852
rect 9582 9800 9588 9852
rect 9640 9840 9646 9852
rect 13998 9840 14004 9852
rect 9640 9812 14004 9840
rect 9640 9800 9646 9812
rect 13998 9800 14004 9812
rect 14056 9800 14062 9852
rect 16942 9800 16948 9852
rect 17000 9840 17006 9852
rect 18966 9840 18972 9852
rect 17000 9812 18972 9840
rect 17000 9800 17006 9812
rect 18966 9800 18972 9812
rect 19024 9800 19030 9852
rect 19058 9800 19064 9852
rect 19116 9840 19122 9852
rect 23566 9840 23572 9852
rect 19116 9812 23572 9840
rect 19116 9800 19122 9812
rect 23566 9800 23572 9812
rect 23624 9800 23630 9852
rect 24118 9800 24124 9852
rect 24176 9840 24182 9852
rect 31726 9840 31754 9880
rect 35618 9868 35624 9880
rect 35676 9868 35682 9920
rect 24176 9812 31754 9840
rect 24176 9800 24182 9812
rect 1762 9732 1768 9784
rect 1820 9772 1826 9784
rect 4338 9772 4344 9784
rect 1820 9744 4344 9772
rect 1820 9732 1826 9744
rect 4338 9732 4344 9744
rect 4396 9732 4402 9784
rect 8570 9732 8576 9784
rect 8628 9772 8634 9784
rect 12342 9772 12348 9784
rect 8628 9744 12348 9772
rect 8628 9732 8634 9744
rect 12342 9732 12348 9744
rect 12400 9732 12406 9784
rect 33778 9772 33784 9784
rect 12452 9744 24256 9772
rect 3418 9664 3424 9716
rect 3476 9704 3482 9716
rect 4614 9704 4620 9716
rect 3476 9676 4620 9704
rect 3476 9664 3482 9676
rect 4614 9664 4620 9676
rect 4672 9664 4678 9716
rect 7190 9664 7196 9716
rect 7248 9704 7254 9716
rect 12066 9704 12072 9716
rect 7248 9676 12072 9704
rect 7248 9664 7254 9676
rect 12066 9664 12072 9676
rect 12124 9664 12130 9716
rect 6362 9596 6368 9648
rect 6420 9636 6426 9648
rect 8938 9636 8944 9648
rect 6420 9608 8944 9636
rect 6420 9596 6426 9608
rect 8938 9596 8944 9608
rect 8996 9596 9002 9648
rect 9030 9596 9036 9648
rect 9088 9636 9094 9648
rect 12452 9636 12480 9744
rect 17126 9664 17132 9716
rect 17184 9704 17190 9716
rect 24118 9704 24124 9716
rect 17184 9676 24124 9704
rect 17184 9664 17190 9676
rect 24118 9664 24124 9676
rect 24176 9664 24182 9716
rect 24228 9704 24256 9744
rect 26896 9744 33784 9772
rect 26896 9704 26924 9744
rect 33778 9732 33784 9744
rect 33836 9732 33842 9784
rect 24228 9676 26924 9704
rect 27798 9664 27804 9716
rect 27856 9704 27862 9716
rect 32306 9704 32312 9716
rect 27856 9676 32312 9704
rect 27856 9664 27862 9676
rect 32306 9664 32312 9676
rect 32364 9664 32370 9716
rect 9088 9608 12480 9636
rect 9088 9596 9094 9608
rect 5902 9528 5908 9580
rect 5960 9568 5966 9580
rect 11790 9568 11796 9580
rect 5960 9540 11796 9568
rect 5960 9528 5966 9540
rect 11790 9528 11796 9540
rect 11848 9528 11854 9580
rect 1670 9460 1676 9512
rect 1728 9500 1734 9512
rect 9766 9500 9772 9512
rect 1728 9472 9772 9500
rect 1728 9460 1734 9472
rect 9766 9460 9772 9472
rect 9824 9460 9830 9512
rect 9858 9460 9864 9512
rect 9916 9500 9922 9512
rect 17126 9500 17132 9512
rect 9916 9472 17132 9500
rect 9916 9460 9922 9472
rect 17126 9460 17132 9472
rect 17184 9460 17190 9512
rect 17494 9460 17500 9512
rect 17552 9500 17558 9512
rect 24394 9500 24400 9512
rect 17552 9472 24400 9500
rect 17552 9460 17558 9472
rect 24394 9460 24400 9472
rect 24452 9460 24458 9512
rect 29546 9500 29552 9512
rect 27586 9472 29552 9500
rect 10778 9432 10784 9444
rect 3804 9404 10784 9432
rect 3804 9296 3832 9404
rect 10778 9392 10784 9404
rect 10836 9392 10842 9444
rect 17954 9432 17960 9444
rect 17144 9404 17960 9432
rect 4246 9324 4252 9376
rect 4304 9364 4310 9376
rect 10318 9364 10324 9376
rect 4304 9336 10324 9364
rect 4304 9324 4310 9336
rect 10318 9324 10324 9336
rect 10376 9324 10382 9376
rect 10502 9324 10508 9376
rect 10560 9364 10566 9376
rect 17144 9364 17172 9404
rect 17954 9392 17960 9404
rect 18012 9392 18018 9444
rect 23658 9392 23664 9444
rect 23716 9432 23722 9444
rect 26418 9432 26424 9444
rect 23716 9404 26424 9432
rect 23716 9392 23722 9404
rect 26418 9392 26424 9404
rect 26476 9392 26482 9444
rect 27338 9392 27344 9444
rect 27396 9432 27402 9444
rect 27586 9432 27614 9472
rect 29546 9460 29552 9472
rect 29604 9460 29610 9512
rect 27396 9404 27614 9432
rect 27396 9392 27402 9404
rect 28994 9392 29000 9444
rect 29052 9432 29058 9444
rect 34238 9432 34244 9444
rect 29052 9404 34244 9432
rect 29052 9392 29058 9404
rect 34238 9392 34244 9404
rect 34296 9392 34302 9444
rect 22738 9364 22744 9376
rect 10560 9336 17172 9364
rect 17236 9336 22744 9364
rect 10560 9324 10566 9336
rect 2746 9268 3832 9296
rect 2130 9188 2136 9240
rect 2188 9228 2194 9240
rect 2746 9228 2774 9268
rect 5626 9256 5632 9308
rect 5684 9296 5690 9308
rect 16298 9296 16304 9308
rect 5684 9268 16304 9296
rect 5684 9256 5690 9268
rect 16298 9256 16304 9268
rect 16356 9256 16362 9308
rect 16850 9256 16856 9308
rect 16908 9296 16914 9308
rect 17236 9296 17264 9336
rect 22738 9324 22744 9336
rect 22796 9324 22802 9376
rect 29822 9364 29828 9376
rect 23676 9336 29828 9364
rect 23676 9308 23704 9336
rect 29822 9324 29828 9336
rect 29880 9324 29886 9376
rect 30006 9324 30012 9376
rect 30064 9364 30070 9376
rect 31294 9364 31300 9376
rect 30064 9336 31300 9364
rect 30064 9324 30070 9336
rect 31294 9324 31300 9336
rect 31352 9324 31358 9376
rect 31386 9324 31392 9376
rect 31444 9364 31450 9376
rect 32582 9364 32588 9376
rect 31444 9336 32588 9364
rect 31444 9324 31450 9336
rect 32582 9324 32588 9336
rect 32640 9324 32646 9376
rect 16908 9268 17264 9296
rect 16908 9256 16914 9268
rect 18598 9256 18604 9308
rect 18656 9296 18662 9308
rect 22830 9296 22836 9308
rect 18656 9268 22836 9296
rect 18656 9256 18662 9268
rect 22830 9256 22836 9268
rect 22888 9256 22894 9308
rect 23658 9256 23664 9308
rect 23716 9256 23722 9308
rect 25406 9256 25412 9308
rect 25464 9296 25470 9308
rect 38562 9296 38568 9308
rect 25464 9268 38568 9296
rect 25464 9256 25470 9268
rect 38562 9256 38568 9268
rect 38620 9256 38626 9308
rect 2188 9200 2774 9228
rect 2188 9188 2194 9200
rect 5534 9188 5540 9240
rect 5592 9228 5598 9240
rect 11698 9228 11704 9240
rect 5592 9200 11704 9228
rect 5592 9188 5598 9200
rect 11698 9188 11704 9200
rect 11756 9188 11762 9240
rect 11790 9188 11796 9240
rect 11848 9228 11854 9240
rect 11848 9200 19334 9228
rect 11848 9188 11854 9200
rect 1854 9120 1860 9172
rect 1912 9160 1918 9172
rect 9674 9160 9680 9172
rect 1912 9132 9680 9160
rect 1912 9120 1918 9132
rect 9674 9120 9680 9132
rect 9732 9120 9738 9172
rect 11330 9120 11336 9172
rect 11388 9160 11394 9172
rect 18046 9160 18052 9172
rect 11388 9132 18052 9160
rect 11388 9120 11394 9132
rect 18046 9120 18052 9132
rect 18104 9120 18110 9172
rect 19306 9160 19334 9200
rect 26142 9188 26148 9240
rect 26200 9228 26206 9240
rect 28810 9228 28816 9240
rect 26200 9200 28816 9228
rect 26200 9188 26206 9200
rect 28810 9188 28816 9200
rect 28868 9188 28874 9240
rect 29730 9188 29736 9240
rect 29788 9228 29794 9240
rect 31570 9228 31576 9240
rect 29788 9200 31576 9228
rect 29788 9188 29794 9200
rect 31570 9188 31576 9200
rect 31628 9188 31634 9240
rect 31938 9188 31944 9240
rect 31996 9228 32002 9240
rect 33962 9228 33968 9240
rect 31996 9200 33968 9228
rect 31996 9188 32002 9200
rect 33962 9188 33968 9200
rect 34020 9188 34026 9240
rect 26326 9160 26332 9172
rect 19306 9132 26332 9160
rect 26326 9120 26332 9132
rect 26384 9120 26390 9172
rect 27798 9120 27804 9172
rect 27856 9160 27862 9172
rect 30926 9160 30932 9172
rect 27856 9132 30932 9160
rect 27856 9120 27862 9132
rect 30926 9120 30932 9132
rect 30984 9120 30990 9172
rect 5442 9052 5448 9104
rect 5500 9092 5506 9104
rect 16850 9092 16856 9104
rect 5500 9064 16856 9092
rect 5500 9052 5506 9064
rect 16850 9052 16856 9064
rect 16908 9052 16914 9104
rect 23842 9052 23848 9104
rect 23900 9092 23906 9104
rect 27890 9092 27896 9104
rect 23900 9064 27896 9092
rect 23900 9052 23906 9064
rect 3602 8984 3608 9036
rect 3660 9024 3666 9036
rect 5994 9024 6000 9036
rect 3660 8996 6000 9024
rect 3660 8984 3666 8996
rect 5994 8984 6000 8996
rect 6052 8984 6058 9036
rect 8018 8984 8024 9036
rect 8076 9024 8082 9036
rect 12066 9024 12072 9036
rect 8076 8996 12072 9024
rect 8076 8984 8082 8996
rect 12066 8984 12072 8996
rect 12124 8984 12130 9036
rect 13078 8984 13084 9036
rect 13136 9024 13142 9036
rect 20530 9024 20536 9036
rect 13136 8996 20536 9024
rect 13136 8984 13142 8996
rect 20530 8984 20536 8996
rect 20588 8984 20594 9036
rect 1394 8916 1400 8968
rect 1452 8956 1458 8968
rect 6914 8956 6920 8968
rect 1452 8928 6920 8956
rect 1452 8916 1458 8928
rect 6914 8916 6920 8928
rect 6972 8916 6978 8968
rect 7742 8916 7748 8968
rect 7800 8956 7806 8968
rect 7800 8928 8791 8956
rect 7800 8916 7806 8928
rect 1578 8848 1584 8900
rect 1636 8888 1642 8900
rect 8110 8888 8116 8900
rect 1636 8860 8116 8888
rect 1636 8848 1642 8860
rect 8110 8848 8116 8860
rect 8168 8848 8174 8900
rect 8763 8888 8791 8928
rect 8846 8916 8852 8968
rect 8904 8956 8910 8968
rect 8904 8928 16620 8956
rect 8904 8916 8910 8928
rect 13078 8888 13084 8900
rect 8763 8860 13084 8888
rect 13078 8848 13084 8860
rect 13136 8848 13142 8900
rect 13262 8848 13268 8900
rect 13320 8888 13326 8900
rect 15194 8888 15200 8900
rect 13320 8860 15200 8888
rect 13320 8848 13326 8860
rect 15194 8848 15200 8860
rect 15252 8848 15258 8900
rect 3878 8780 3884 8832
rect 3936 8820 3942 8832
rect 9030 8820 9036 8832
rect 3936 8792 9036 8820
rect 3936 8780 3942 8792
rect 9030 8780 9036 8792
rect 9088 8780 9094 8832
rect 11790 8780 11796 8832
rect 11848 8820 11854 8832
rect 14734 8820 14740 8832
rect 11848 8792 14740 8820
rect 11848 8780 11854 8792
rect 14734 8780 14740 8792
rect 14792 8780 14798 8832
rect 16022 8780 16028 8832
rect 16080 8820 16086 8832
rect 16482 8820 16488 8832
rect 16080 8792 16488 8820
rect 16080 8780 16086 8792
rect 16482 8780 16488 8792
rect 16540 8780 16546 8832
rect 16592 8820 16620 8928
rect 18230 8916 18236 8968
rect 18288 8956 18294 8968
rect 24026 8956 24032 8968
rect 18288 8928 24032 8956
rect 18288 8916 18294 8928
rect 24026 8916 24032 8928
rect 24084 8916 24090 8968
rect 18966 8848 18972 8900
rect 19024 8888 19030 8900
rect 24136 8888 24164 9064
rect 27890 9052 27896 9064
rect 27948 9052 27954 9104
rect 29362 9052 29368 9104
rect 29420 9092 29426 9104
rect 34974 9092 34980 9104
rect 29420 9064 34980 9092
rect 29420 9052 29426 9064
rect 34974 9052 34980 9064
rect 35032 9052 35038 9104
rect 24302 8984 24308 9036
rect 24360 9024 24366 9036
rect 30098 9024 30104 9036
rect 24360 8996 30104 9024
rect 24360 8984 24366 8996
rect 30098 8984 30104 8996
rect 30156 8984 30162 9036
rect 32214 8984 32220 9036
rect 32272 9024 32278 9036
rect 34790 9024 34796 9036
rect 32272 8996 34796 9024
rect 32272 8984 32278 8996
rect 34790 8984 34796 8996
rect 34848 8984 34854 9036
rect 26510 8916 26516 8968
rect 26568 8956 26574 8968
rect 31754 8956 31760 8968
rect 26568 8928 31760 8956
rect 26568 8916 26574 8928
rect 31754 8916 31760 8928
rect 31812 8916 31818 8968
rect 33042 8916 33048 8968
rect 33100 8956 33106 8968
rect 34514 8956 34520 8968
rect 33100 8928 34520 8956
rect 33100 8916 33106 8928
rect 34514 8916 34520 8928
rect 34572 8916 34578 8968
rect 35342 8916 35348 8968
rect 35400 8956 35406 8968
rect 38378 8956 38384 8968
rect 35400 8928 38384 8956
rect 35400 8916 35406 8928
rect 38378 8916 38384 8928
rect 38436 8916 38442 8968
rect 19024 8860 24164 8888
rect 19024 8848 19030 8860
rect 25590 8848 25596 8900
rect 25648 8888 25654 8900
rect 26878 8888 26884 8900
rect 25648 8860 26884 8888
rect 25648 8848 25654 8860
rect 26878 8848 26884 8860
rect 26936 8848 26942 8900
rect 27522 8848 27528 8900
rect 27580 8888 27586 8900
rect 32122 8888 32128 8900
rect 27580 8860 32128 8888
rect 27580 8848 27586 8860
rect 32122 8848 32128 8860
rect 32180 8848 32186 8900
rect 34330 8848 34336 8900
rect 34388 8888 34394 8900
rect 36538 8888 36544 8900
rect 34388 8860 36544 8888
rect 34388 8848 34394 8860
rect 36538 8848 36544 8860
rect 36596 8848 36602 8900
rect 21542 8820 21548 8832
rect 16592 8792 21548 8820
rect 21542 8780 21548 8792
rect 21600 8780 21606 8832
rect 22830 8780 22836 8832
rect 22888 8820 22894 8832
rect 23842 8820 23848 8832
rect 22888 8792 23848 8820
rect 22888 8780 22894 8792
rect 23842 8780 23848 8792
rect 23900 8780 23906 8832
rect 25314 8780 25320 8832
rect 25372 8820 25378 8832
rect 30190 8820 30196 8832
rect 25372 8792 30196 8820
rect 25372 8780 25378 8792
rect 30190 8780 30196 8792
rect 30248 8780 30254 8832
rect 33318 8780 33324 8832
rect 33376 8820 33382 8832
rect 33778 8820 33784 8832
rect 33376 8792 33784 8820
rect 33376 8780 33382 8792
rect 33778 8780 33784 8792
rect 33836 8780 33842 8832
rect 35710 8780 35716 8832
rect 35768 8820 35774 8832
rect 37366 8820 37372 8832
rect 35768 8792 37372 8820
rect 35768 8780 35774 8792
rect 37366 8780 37372 8792
rect 37424 8780 37430 8832
rect 1104 8730 39836 8752
rect 1104 8678 3010 8730
rect 3062 8678 3074 8730
rect 3126 8678 3138 8730
rect 3190 8678 3202 8730
rect 3254 8678 3266 8730
rect 3318 8678 9010 8730
rect 9062 8678 9074 8730
rect 9126 8678 9138 8730
rect 9190 8678 9202 8730
rect 9254 8678 9266 8730
rect 9318 8678 15010 8730
rect 15062 8678 15074 8730
rect 15126 8678 15138 8730
rect 15190 8678 15202 8730
rect 15254 8678 15266 8730
rect 15318 8678 21010 8730
rect 21062 8678 21074 8730
rect 21126 8678 21138 8730
rect 21190 8678 21202 8730
rect 21254 8678 21266 8730
rect 21318 8678 27010 8730
rect 27062 8678 27074 8730
rect 27126 8678 27138 8730
rect 27190 8678 27202 8730
rect 27254 8678 27266 8730
rect 27318 8678 33010 8730
rect 33062 8678 33074 8730
rect 33126 8678 33138 8730
rect 33190 8678 33202 8730
rect 33254 8678 33266 8730
rect 33318 8678 39010 8730
rect 39062 8678 39074 8730
rect 39126 8678 39138 8730
rect 39190 8678 39202 8730
rect 39254 8678 39266 8730
rect 39318 8678 39836 8730
rect 1104 8656 39836 8678
rect 1578 8576 1584 8628
rect 1636 8576 1642 8628
rect 3510 8576 3516 8628
rect 3568 8576 3574 8628
rect 3881 8619 3939 8625
rect 3881 8585 3893 8619
rect 3927 8616 3939 8619
rect 4430 8616 4436 8628
rect 3927 8588 4436 8616
rect 3927 8585 3939 8588
rect 3881 8579 3939 8585
rect 4430 8576 4436 8588
rect 4488 8576 4494 8628
rect 5442 8576 5448 8628
rect 5500 8576 5506 8628
rect 5721 8619 5779 8625
rect 5721 8585 5733 8619
rect 5767 8616 5779 8619
rect 5810 8616 5816 8628
rect 5767 8588 5816 8616
rect 5767 8585 5779 8588
rect 5721 8579 5779 8585
rect 5810 8576 5816 8588
rect 5868 8576 5874 8628
rect 6086 8576 6092 8628
rect 6144 8576 6150 8628
rect 6549 8619 6607 8625
rect 6549 8585 6561 8619
rect 6595 8616 6607 8619
rect 6638 8616 6644 8628
rect 6595 8588 6644 8616
rect 6595 8585 6607 8588
rect 6549 8579 6607 8585
rect 6638 8576 6644 8588
rect 6696 8576 6702 8628
rect 6917 8619 6975 8625
rect 6917 8585 6929 8619
rect 6963 8616 6975 8619
rect 7006 8616 7012 8628
rect 6963 8588 7012 8616
rect 6963 8585 6975 8588
rect 6917 8579 6975 8585
rect 7006 8576 7012 8588
rect 7064 8576 7070 8628
rect 7101 8619 7159 8625
rect 7101 8585 7113 8619
rect 7147 8616 7159 8619
rect 7190 8616 7196 8628
rect 7147 8588 7196 8616
rect 7147 8585 7159 8588
rect 7101 8579 7159 8585
rect 7190 8576 7196 8588
rect 7248 8576 7254 8628
rect 7469 8619 7527 8625
rect 7469 8585 7481 8619
rect 7515 8616 7527 8619
rect 7742 8616 7748 8628
rect 7515 8588 7748 8616
rect 7515 8585 7527 8588
rect 7469 8579 7527 8585
rect 7742 8576 7748 8588
rect 7800 8576 7806 8628
rect 8297 8619 8355 8625
rect 8297 8585 8309 8619
rect 8343 8616 8355 8619
rect 8386 8616 8392 8628
rect 8343 8588 8392 8616
rect 8343 8585 8355 8588
rect 8297 8579 8355 8585
rect 8386 8576 8392 8588
rect 8444 8576 8450 8628
rect 8570 8576 8576 8628
rect 8628 8576 8634 8628
rect 9125 8619 9183 8625
rect 9125 8585 9137 8619
rect 9171 8616 9183 8619
rect 9582 8616 9588 8628
rect 9171 8588 9588 8616
rect 9171 8585 9183 8588
rect 9125 8579 9183 8585
rect 9582 8576 9588 8588
rect 9640 8576 9646 8628
rect 10505 8619 10563 8625
rect 10505 8585 10517 8619
rect 10551 8585 10563 8619
rect 10505 8579 10563 8585
rect 3970 8548 3976 8560
rect 1964 8520 3976 8548
rect 1394 8440 1400 8492
rect 1452 8440 1458 8492
rect 1670 8440 1676 8492
rect 1728 8440 1734 8492
rect 1854 8440 1860 8492
rect 1912 8440 1918 8492
rect 1964 8489 1992 8520
rect 3970 8508 3976 8520
rect 4028 8508 4034 8560
rect 9490 8548 9496 8560
rect 4080 8520 9496 8548
rect 1949 8483 2007 8489
rect 1949 8449 1961 8483
rect 1995 8449 2007 8483
rect 1949 8443 2007 8449
rect 2130 8440 2136 8492
rect 2188 8440 2194 8492
rect 2498 8440 2504 8492
rect 2556 8440 2562 8492
rect 3237 8483 3295 8489
rect 3237 8449 3249 8483
rect 3283 8480 3295 8483
rect 3329 8483 3387 8489
rect 3329 8480 3341 8483
rect 3283 8452 3341 8480
rect 3283 8449 3295 8452
rect 3237 8443 3295 8449
rect 3329 8449 3341 8452
rect 3375 8480 3387 8483
rect 3878 8480 3884 8492
rect 3375 8452 3884 8480
rect 3375 8449 3387 8452
rect 3329 8443 3387 8449
rect 3878 8440 3884 8452
rect 3936 8440 3942 8492
rect 1118 8372 1124 8424
rect 1176 8412 1182 8424
rect 2225 8415 2283 8421
rect 2225 8412 2237 8415
rect 1176 8384 2237 8412
rect 1176 8372 1182 8384
rect 2225 8381 2237 8384
rect 2271 8381 2283 8415
rect 4080 8412 4108 8520
rect 9490 8508 9496 8520
rect 9548 8508 9554 8560
rect 10520 8548 10548 8579
rect 11238 8576 11244 8628
rect 11296 8616 11302 8628
rect 11606 8616 11612 8628
rect 11296 8588 11612 8616
rect 11296 8576 11302 8588
rect 11606 8576 11612 8588
rect 11664 8576 11670 8628
rect 11790 8576 11796 8628
rect 11848 8576 11854 8628
rect 12986 8616 12992 8628
rect 11900 8588 12992 8616
rect 11900 8548 11928 8588
rect 12986 8576 12992 8588
rect 13044 8576 13050 8628
rect 13081 8619 13139 8625
rect 13081 8585 13093 8619
rect 13127 8616 13139 8619
rect 14918 8616 14924 8628
rect 13127 8588 14924 8616
rect 13127 8585 13139 8588
rect 13081 8579 13139 8585
rect 14918 8576 14924 8588
rect 14976 8576 14982 8628
rect 15197 8619 15255 8625
rect 15197 8585 15209 8619
rect 15243 8585 15255 8619
rect 15197 8579 15255 8585
rect 15565 8619 15623 8625
rect 15565 8585 15577 8619
rect 15611 8616 15623 8619
rect 16206 8616 16212 8628
rect 15611 8588 16212 8616
rect 15611 8585 15623 8588
rect 15565 8579 15623 8585
rect 10520 8520 11928 8548
rect 12066 8508 12072 8560
rect 12124 8548 12130 8560
rect 12124 8520 13676 8548
rect 12124 8508 12130 8520
rect 4798 8440 4804 8492
rect 4856 8480 4862 8492
rect 4985 8483 5043 8489
rect 4985 8480 4997 8483
rect 4856 8452 4997 8480
rect 4856 8440 4862 8452
rect 4985 8449 4997 8452
rect 5031 8449 5043 8483
rect 4985 8443 5043 8449
rect 5445 8483 5503 8489
rect 5445 8449 5457 8483
rect 5491 8480 5503 8483
rect 5537 8483 5595 8489
rect 5537 8480 5549 8483
rect 5491 8452 5549 8480
rect 5491 8449 5503 8452
rect 5445 8443 5503 8449
rect 5537 8449 5549 8452
rect 5583 8449 5595 8483
rect 5537 8443 5595 8449
rect 5905 8483 5963 8489
rect 5905 8449 5917 8483
rect 5951 8480 5963 8483
rect 5994 8480 6000 8492
rect 5951 8452 6000 8480
rect 5951 8449 5963 8452
rect 5905 8443 5963 8449
rect 5994 8440 6000 8452
rect 6052 8440 6058 8492
rect 6733 8483 6791 8489
rect 6733 8449 6745 8483
rect 6779 8480 6791 8483
rect 6825 8483 6883 8489
rect 6825 8480 6837 8483
rect 6779 8452 6837 8480
rect 6779 8449 6791 8452
rect 6733 8443 6791 8449
rect 6825 8449 6837 8452
rect 6871 8449 6883 8483
rect 6825 8443 6883 8449
rect 7285 8483 7343 8489
rect 7285 8449 7297 8483
rect 7331 8480 7343 8483
rect 7377 8483 7435 8489
rect 7377 8480 7389 8483
rect 7331 8452 7389 8480
rect 7331 8449 7343 8452
rect 7285 8443 7343 8449
rect 7377 8449 7389 8452
rect 7423 8449 7435 8483
rect 7377 8443 7435 8449
rect 7650 8440 7656 8492
rect 7708 8480 7714 8492
rect 7745 8483 7803 8489
rect 7745 8480 7757 8483
rect 7708 8452 7757 8480
rect 7708 8440 7714 8452
rect 7745 8449 7757 8452
rect 7791 8449 7803 8483
rect 7745 8443 7803 8449
rect 8110 8440 8116 8492
rect 8168 8440 8174 8492
rect 8754 8440 8760 8492
rect 8812 8440 8818 8492
rect 9309 8483 9367 8489
rect 9309 8449 9321 8483
rect 9355 8480 9367 8483
rect 9355 8452 10272 8480
rect 9355 8449 9367 8452
rect 9309 8443 9367 8449
rect 2225 8375 2283 8381
rect 2746 8384 4108 8412
rect 4525 8415 4583 8421
rect 2041 8347 2099 8353
rect 2041 8313 2053 8347
rect 2087 8344 2099 8347
rect 2746 8344 2774 8384
rect 4525 8381 4537 8415
rect 4571 8381 4583 8415
rect 4525 8375 4583 8381
rect 4065 8347 4123 8353
rect 4065 8344 4077 8347
rect 2087 8316 2774 8344
rect 2884 8316 4077 8344
rect 2087 8313 2099 8316
rect 2041 8307 2099 8313
rect 1765 8279 1823 8285
rect 1765 8245 1777 8279
rect 1811 8276 1823 8279
rect 2590 8276 2596 8288
rect 1811 8248 2596 8276
rect 1811 8245 1823 8248
rect 1765 8239 1823 8245
rect 2590 8236 2596 8248
rect 2648 8236 2654 8288
rect 2682 8236 2688 8288
rect 2740 8276 2746 8288
rect 2884 8276 2912 8316
rect 4065 8313 4077 8316
rect 4111 8313 4123 8347
rect 4540 8344 4568 8375
rect 4706 8372 4712 8424
rect 4764 8372 4770 8424
rect 5184 8384 8340 8412
rect 5184 8353 5212 8384
rect 5169 8347 5227 8353
rect 4540 8316 5120 8344
rect 4065 8307 4123 8313
rect 2740 8248 2912 8276
rect 5092 8276 5120 8316
rect 5169 8313 5181 8347
rect 5215 8313 5227 8347
rect 6086 8344 6092 8356
rect 5169 8307 5227 8313
rect 5276 8316 6092 8344
rect 5276 8276 5304 8316
rect 6086 8304 6092 8316
rect 6144 8344 6150 8356
rect 6144 8316 7604 8344
rect 6144 8304 6150 8316
rect 5092 8248 5304 8276
rect 2740 8236 2746 8248
rect 6638 8236 6644 8288
rect 6696 8276 6702 8288
rect 7466 8276 7472 8288
rect 6696 8248 7472 8276
rect 6696 8236 6702 8248
rect 7466 8236 7472 8248
rect 7524 8236 7530 8288
rect 7576 8276 7604 8316
rect 7926 8304 7932 8356
rect 7984 8304 7990 8356
rect 8312 8344 8340 8384
rect 8386 8372 8392 8424
rect 8444 8412 8450 8424
rect 8938 8412 8944 8424
rect 8444 8384 8944 8412
rect 8444 8372 8450 8384
rect 8938 8372 8944 8384
rect 8996 8372 9002 8424
rect 9214 8372 9220 8424
rect 9272 8412 9278 8424
rect 9401 8415 9459 8421
rect 9401 8412 9413 8415
rect 9272 8384 9413 8412
rect 9272 8372 9278 8384
rect 9401 8381 9413 8384
rect 9447 8412 9459 8415
rect 9582 8412 9588 8424
rect 9447 8384 9588 8412
rect 9447 8381 9459 8384
rect 9401 8375 9459 8381
rect 9582 8372 9588 8384
rect 9640 8372 9646 8424
rect 9950 8372 9956 8424
rect 10008 8372 10014 8424
rect 10244 8412 10272 8452
rect 10318 8440 10324 8492
rect 10376 8440 10382 8492
rect 10962 8440 10968 8492
rect 11020 8480 11026 8492
rect 11609 8483 11667 8489
rect 11020 8452 11560 8480
rect 11020 8440 11026 8452
rect 11238 8412 11244 8424
rect 10244 8384 11244 8412
rect 11238 8372 11244 8384
rect 11296 8372 11302 8424
rect 11333 8415 11391 8421
rect 11333 8381 11345 8415
rect 11379 8412 11391 8415
rect 11422 8412 11428 8424
rect 11379 8384 11428 8412
rect 11379 8381 11391 8384
rect 11333 8375 11391 8381
rect 11422 8372 11428 8384
rect 11480 8372 11486 8424
rect 11532 8412 11560 8452
rect 11609 8449 11621 8483
rect 11655 8480 11667 8483
rect 11698 8480 11704 8492
rect 11655 8452 11704 8480
rect 11655 8449 11667 8452
rect 11609 8443 11667 8449
rect 11698 8440 11704 8452
rect 11756 8440 11762 8492
rect 11974 8440 11980 8492
rect 12032 8440 12038 8492
rect 12161 8483 12219 8489
rect 12161 8449 12173 8483
rect 12207 8449 12219 8483
rect 12161 8443 12219 8449
rect 12253 8483 12311 8489
rect 12253 8449 12265 8483
rect 12299 8449 12311 8483
rect 12253 8443 12311 8449
rect 12345 8483 12403 8489
rect 12345 8449 12357 8483
rect 12391 8480 12403 8483
rect 12710 8480 12716 8492
rect 12391 8452 12716 8480
rect 12391 8449 12403 8452
rect 12345 8443 12403 8449
rect 12176 8412 12204 8443
rect 11532 8384 12204 8412
rect 12268 8412 12296 8443
rect 12710 8440 12716 8452
rect 12768 8440 12774 8492
rect 12802 8440 12808 8492
rect 12860 8480 12866 8492
rect 12897 8483 12955 8489
rect 12897 8480 12909 8483
rect 12860 8452 12909 8480
rect 12860 8440 12866 8452
rect 12897 8449 12909 8452
rect 12943 8449 12955 8483
rect 12897 8443 12955 8449
rect 13538 8440 13544 8492
rect 13596 8440 13602 8492
rect 13648 8489 13676 8520
rect 13722 8508 13728 8560
rect 13780 8548 13786 8560
rect 14642 8548 14648 8560
rect 13780 8520 14648 8548
rect 13780 8508 13786 8520
rect 14642 8508 14648 8520
rect 14700 8508 14706 8560
rect 14734 8508 14740 8560
rect 14792 8508 14798 8560
rect 15212 8548 15240 8579
rect 16206 8576 16212 8588
rect 16264 8576 16270 8628
rect 16301 8619 16359 8625
rect 16301 8585 16313 8619
rect 16347 8616 16359 8619
rect 16758 8616 16764 8628
rect 16347 8588 16764 8616
rect 16347 8585 16359 8588
rect 16301 8579 16359 8585
rect 16758 8576 16764 8588
rect 16816 8576 16822 8628
rect 17034 8576 17040 8628
rect 17092 8616 17098 8628
rect 18049 8619 18107 8625
rect 18049 8616 18061 8619
rect 17092 8588 18061 8616
rect 17092 8576 17098 8588
rect 18049 8585 18061 8588
rect 18095 8585 18107 8619
rect 18049 8579 18107 8585
rect 18322 8576 18328 8628
rect 18380 8576 18386 8628
rect 18414 8576 18420 8628
rect 18472 8616 18478 8628
rect 20625 8619 20683 8625
rect 20625 8616 20637 8619
rect 18472 8588 20637 8616
rect 18472 8576 18478 8588
rect 20625 8585 20637 8588
rect 20671 8585 20683 8619
rect 23845 8619 23903 8625
rect 23845 8616 23857 8619
rect 20625 8579 20683 8585
rect 23676 8588 23857 8616
rect 15930 8548 15936 8560
rect 15212 8520 15936 8548
rect 15930 8508 15936 8520
rect 15988 8508 15994 8560
rect 16669 8551 16727 8557
rect 16669 8548 16681 8551
rect 16040 8520 16681 8548
rect 13633 8483 13691 8489
rect 13633 8449 13645 8483
rect 13679 8449 13691 8483
rect 13633 8443 13691 8449
rect 14016 8452 14412 8480
rect 12986 8412 12992 8424
rect 12268 8384 12992 8412
rect 12986 8372 12992 8384
rect 13044 8372 13050 8424
rect 14016 8412 14044 8452
rect 13372 8384 14044 8412
rect 11514 8344 11520 8356
rect 8312 8316 11520 8344
rect 11514 8304 11520 8316
rect 11572 8304 11578 8356
rect 11974 8304 11980 8356
rect 12032 8344 12038 8356
rect 13372 8353 13400 8384
rect 14090 8372 14096 8424
rect 14148 8372 14154 8424
rect 14384 8412 14412 8452
rect 14826 8440 14832 8492
rect 14884 8480 14890 8492
rect 15013 8483 15071 8489
rect 15013 8480 15025 8483
rect 14884 8452 15025 8480
rect 14884 8440 14890 8452
rect 15013 8449 15025 8452
rect 15059 8449 15071 8483
rect 15013 8443 15071 8449
rect 15286 8440 15292 8492
rect 15344 8440 15350 8492
rect 15381 8483 15439 8489
rect 15381 8449 15393 8483
rect 15427 8480 15439 8483
rect 15562 8480 15568 8492
rect 15427 8452 15568 8480
rect 15427 8449 15439 8452
rect 15381 8443 15439 8449
rect 15562 8440 15568 8452
rect 15620 8440 15626 8492
rect 15746 8440 15752 8492
rect 15804 8440 15810 8492
rect 15304 8412 15332 8440
rect 16040 8412 16068 8520
rect 16669 8517 16681 8520
rect 16715 8517 16727 8551
rect 16669 8511 16727 8517
rect 16850 8508 16856 8560
rect 16908 8548 16914 8560
rect 19705 8551 19763 8557
rect 19705 8548 19717 8551
rect 16908 8520 17632 8548
rect 16908 8508 16914 8520
rect 16117 8483 16175 8489
rect 16117 8449 16129 8483
rect 16163 8449 16175 8483
rect 16117 8443 16175 8449
rect 16485 8483 16543 8489
rect 16485 8449 16497 8483
rect 16531 8480 16543 8483
rect 17494 8480 17500 8492
rect 16531 8452 17500 8480
rect 16531 8449 16543 8452
rect 16485 8443 16543 8449
rect 14384 8384 15332 8412
rect 15764 8384 16068 8412
rect 16132 8412 16160 8443
rect 17494 8440 17500 8452
rect 17552 8440 17558 8492
rect 17604 8489 17632 8520
rect 17880 8520 19717 8548
rect 17880 8489 17908 8520
rect 19705 8517 19717 8520
rect 19751 8517 19763 8551
rect 19705 8511 19763 8517
rect 22572 8520 23152 8548
rect 17589 8483 17647 8489
rect 17589 8449 17601 8483
rect 17635 8449 17647 8483
rect 17589 8443 17647 8449
rect 17865 8483 17923 8489
rect 17865 8449 17877 8483
rect 17911 8449 17923 8483
rect 17865 8443 17923 8449
rect 16132 8384 16344 8412
rect 13357 8347 13415 8353
rect 12032 8316 12756 8344
rect 12032 8304 12038 8316
rect 8386 8276 8392 8288
rect 7576 8248 8392 8276
rect 8386 8236 8392 8248
rect 8444 8236 8450 8288
rect 8754 8236 8760 8288
rect 8812 8276 8818 8288
rect 9398 8276 9404 8288
rect 8812 8248 9404 8276
rect 8812 8236 8818 8248
rect 9398 8236 9404 8248
rect 9456 8236 9462 8288
rect 9766 8236 9772 8288
rect 9824 8276 9830 8288
rect 10502 8276 10508 8288
rect 9824 8248 10508 8276
rect 9824 8236 9830 8248
rect 10502 8236 10508 8248
rect 10560 8236 10566 8288
rect 10689 8279 10747 8285
rect 10689 8245 10701 8279
rect 10735 8276 10747 8279
rect 10778 8276 10784 8288
rect 10735 8248 10784 8276
rect 10735 8245 10747 8248
rect 10689 8239 10747 8245
rect 10778 8236 10784 8248
rect 10836 8236 10842 8288
rect 11054 8236 11060 8288
rect 11112 8276 11118 8288
rect 11882 8276 11888 8288
rect 11112 8248 11888 8276
rect 11112 8236 11118 8248
rect 11882 8236 11888 8248
rect 11940 8236 11946 8288
rect 12618 8236 12624 8288
rect 12676 8236 12682 8288
rect 12728 8276 12756 8316
rect 13357 8313 13369 8347
rect 13403 8313 13415 8347
rect 13357 8307 13415 8313
rect 13817 8347 13875 8353
rect 13817 8313 13829 8347
rect 13863 8344 13875 8347
rect 15654 8344 15660 8356
rect 13863 8316 15660 8344
rect 13863 8313 13875 8316
rect 13817 8307 13875 8313
rect 15654 8304 15660 8316
rect 15712 8304 15718 8356
rect 14458 8276 14464 8288
rect 12728 8248 14464 8276
rect 14458 8236 14464 8248
rect 14516 8236 14522 8288
rect 14826 8236 14832 8288
rect 14884 8236 14890 8288
rect 14918 8236 14924 8288
rect 14976 8276 14982 8288
rect 15764 8276 15792 8384
rect 15933 8347 15991 8353
rect 15933 8313 15945 8347
rect 15979 8344 15991 8347
rect 16022 8344 16028 8356
rect 15979 8316 16028 8344
rect 15979 8313 15991 8316
rect 15933 8307 15991 8313
rect 16022 8304 16028 8316
rect 16080 8304 16086 8356
rect 14976 8248 15792 8276
rect 16316 8276 16344 8384
rect 16390 8372 16396 8424
rect 16448 8412 16454 8424
rect 16448 8384 16620 8412
rect 16448 8372 16454 8384
rect 16592 8344 16620 8384
rect 16666 8372 16672 8424
rect 16724 8412 16730 8424
rect 17221 8415 17279 8421
rect 17221 8412 17233 8415
rect 16724 8384 17233 8412
rect 16724 8372 16730 8384
rect 17221 8381 17233 8384
rect 17267 8381 17279 8415
rect 17221 8375 17279 8381
rect 17402 8372 17408 8424
rect 17460 8372 17466 8424
rect 17604 8412 17632 8443
rect 18230 8440 18236 8492
rect 18288 8440 18294 8492
rect 18509 8483 18567 8489
rect 18509 8449 18521 8483
rect 18555 8480 18567 8483
rect 18555 8452 18920 8480
rect 18555 8449 18567 8452
rect 18509 8443 18567 8449
rect 17604 8384 18644 8412
rect 18616 8356 18644 8384
rect 18690 8372 18696 8424
rect 18748 8372 18754 8424
rect 18785 8415 18843 8421
rect 18785 8381 18797 8415
rect 18831 8381 18843 8415
rect 18892 8412 18920 8452
rect 18966 8440 18972 8492
rect 19024 8440 19030 8492
rect 19058 8440 19064 8492
rect 19116 8440 19122 8492
rect 19429 8483 19487 8489
rect 19429 8449 19441 8483
rect 19475 8480 19487 8483
rect 20898 8480 20904 8492
rect 19475 8452 20904 8480
rect 19475 8449 19487 8452
rect 19429 8443 19487 8449
rect 20898 8440 20904 8452
rect 20956 8440 20962 8492
rect 21450 8440 21456 8492
rect 21508 8440 21514 8492
rect 18892 8384 20300 8412
rect 18785 8375 18843 8381
rect 17773 8347 17831 8353
rect 17773 8344 17785 8347
rect 16592 8316 17785 8344
rect 17773 8313 17785 8316
rect 17819 8313 17831 8347
rect 17773 8307 17831 8313
rect 17880 8316 18552 8344
rect 17880 8276 17908 8316
rect 16316 8248 17908 8276
rect 18524 8276 18552 8316
rect 18598 8304 18604 8356
rect 18656 8344 18662 8356
rect 18800 8344 18828 8375
rect 18656 8316 18828 8344
rect 18877 8347 18935 8353
rect 18656 8304 18662 8316
rect 18877 8313 18889 8347
rect 18923 8344 18935 8347
rect 18966 8344 18972 8356
rect 18923 8316 18972 8344
rect 18923 8313 18935 8316
rect 18877 8307 18935 8313
rect 18966 8304 18972 8316
rect 19024 8304 19030 8356
rect 19518 8344 19524 8356
rect 19168 8316 19524 8344
rect 19168 8276 19196 8316
rect 19518 8304 19524 8316
rect 19576 8304 19582 8356
rect 19613 8347 19671 8353
rect 19613 8313 19625 8347
rect 19659 8344 19671 8347
rect 20272 8344 20300 8384
rect 20346 8372 20352 8424
rect 20404 8412 20410 8424
rect 21082 8412 21088 8424
rect 20404 8384 21088 8412
rect 20404 8372 20410 8384
rect 21082 8372 21088 8384
rect 21140 8372 21146 8424
rect 21269 8415 21327 8421
rect 21269 8381 21281 8415
rect 21315 8412 21327 8415
rect 21358 8412 21364 8424
rect 21315 8384 21364 8412
rect 21315 8381 21327 8384
rect 21269 8375 21327 8381
rect 21358 8372 21364 8384
rect 21416 8372 21422 8424
rect 21634 8372 21640 8424
rect 21692 8412 21698 8424
rect 22005 8415 22063 8421
rect 22005 8412 22017 8415
rect 21692 8384 22017 8412
rect 21692 8372 21698 8384
rect 22005 8381 22017 8384
rect 22051 8412 22063 8415
rect 22572 8412 22600 8520
rect 22830 8440 22836 8492
rect 22888 8480 22894 8492
rect 23017 8483 23075 8489
rect 23017 8480 23029 8483
rect 22888 8452 23029 8480
rect 22888 8440 22894 8452
rect 23017 8449 23029 8452
rect 23063 8449 23075 8483
rect 23124 8480 23152 8520
rect 23198 8508 23204 8560
rect 23256 8548 23262 8560
rect 23676 8548 23704 8588
rect 23845 8585 23857 8588
rect 23891 8585 23903 8619
rect 23845 8579 23903 8585
rect 24118 8576 24124 8628
rect 24176 8616 24182 8628
rect 24765 8619 24823 8625
rect 24765 8616 24777 8619
rect 24176 8588 24777 8616
rect 24176 8576 24182 8588
rect 24765 8585 24777 8588
rect 24811 8585 24823 8619
rect 24765 8579 24823 8585
rect 25222 8576 25228 8628
rect 25280 8576 25286 8628
rect 27801 8619 27859 8625
rect 25608 8588 27752 8616
rect 23256 8520 23704 8548
rect 23256 8508 23262 8520
rect 23750 8508 23756 8560
rect 23808 8548 23814 8560
rect 23997 8551 24055 8557
rect 23997 8548 24009 8551
rect 23808 8520 24009 8548
rect 23808 8508 23814 8520
rect 23997 8517 24009 8520
rect 24043 8517 24055 8551
rect 23997 8511 24055 8517
rect 24213 8551 24271 8557
rect 24213 8517 24225 8551
rect 24259 8548 24271 8551
rect 24486 8548 24492 8560
rect 24259 8520 24492 8548
rect 24259 8517 24271 8520
rect 24213 8511 24271 8517
rect 24486 8508 24492 8520
rect 24544 8508 24550 8560
rect 24578 8508 24584 8560
rect 24636 8548 24642 8560
rect 24673 8551 24731 8557
rect 24673 8548 24685 8551
rect 24636 8520 24685 8548
rect 24636 8508 24642 8520
rect 24673 8517 24685 8520
rect 24719 8517 24731 8551
rect 24673 8511 24731 8517
rect 25608 8489 25636 8588
rect 25866 8508 25872 8560
rect 25924 8548 25930 8560
rect 25924 8520 27660 8548
rect 25924 8508 25930 8520
rect 25439 8483 25497 8489
rect 25439 8480 25451 8483
rect 23124 8452 25451 8480
rect 23017 8443 23075 8449
rect 25439 8449 25451 8452
rect 25485 8449 25497 8483
rect 25439 8443 25497 8449
rect 25593 8483 25651 8489
rect 25593 8449 25605 8483
rect 25639 8449 25651 8483
rect 25593 8443 25651 8449
rect 22051 8384 22600 8412
rect 22649 8415 22707 8421
rect 22051 8381 22063 8384
rect 22005 8375 22063 8381
rect 22649 8381 22661 8415
rect 22695 8412 22707 8415
rect 22741 8415 22799 8421
rect 22741 8412 22753 8415
rect 22695 8384 22753 8412
rect 22695 8381 22707 8384
rect 22649 8375 22707 8381
rect 22741 8381 22753 8384
rect 22787 8381 22799 8415
rect 22741 8375 22799 8381
rect 22922 8372 22928 8424
rect 22980 8412 22986 8424
rect 23198 8412 23204 8424
rect 22980 8384 23204 8412
rect 22980 8372 22986 8384
rect 23198 8372 23204 8384
rect 23256 8372 23262 8424
rect 23566 8372 23572 8424
rect 23624 8412 23630 8424
rect 23753 8415 23811 8421
rect 23753 8412 23765 8415
rect 23624 8384 23765 8412
rect 23624 8372 23630 8384
rect 23753 8381 23765 8384
rect 23799 8412 23811 8415
rect 24302 8412 24308 8424
rect 23799 8384 24308 8412
rect 23799 8381 23811 8384
rect 23753 8375 23811 8381
rect 24302 8372 24308 8384
rect 24360 8372 24366 8424
rect 24581 8415 24639 8421
rect 24581 8381 24593 8415
rect 24627 8381 24639 8415
rect 24581 8375 24639 8381
rect 21726 8344 21732 8356
rect 19659 8316 20208 8344
rect 20272 8316 21732 8344
rect 19659 8313 19671 8316
rect 19613 8307 19671 8313
rect 18524 8248 19196 8276
rect 20180 8276 20208 8316
rect 21726 8304 21732 8316
rect 21784 8304 21790 8356
rect 22833 8347 22891 8353
rect 22833 8313 22845 8347
rect 22879 8344 22891 8347
rect 23293 8347 23351 8353
rect 23293 8344 23305 8347
rect 22879 8316 23305 8344
rect 22879 8313 22891 8316
rect 22833 8307 22891 8313
rect 23293 8313 23305 8316
rect 23339 8313 23351 8347
rect 23293 8307 23351 8313
rect 23382 8304 23388 8356
rect 23440 8344 23446 8356
rect 23477 8347 23535 8353
rect 23477 8344 23489 8347
rect 23440 8316 23489 8344
rect 23440 8304 23446 8316
rect 23477 8313 23489 8316
rect 23523 8344 23535 8347
rect 24596 8344 24624 8375
rect 24670 8372 24676 8424
rect 24728 8412 24734 8424
rect 25608 8412 25636 8443
rect 25682 8440 25688 8492
rect 25740 8480 25746 8492
rect 26053 8483 26111 8489
rect 26053 8480 26065 8483
rect 25740 8452 26065 8480
rect 25740 8440 25746 8452
rect 26053 8449 26065 8452
rect 26099 8449 26111 8483
rect 26053 8443 26111 8449
rect 27062 8440 27068 8492
rect 27120 8440 27126 8492
rect 27632 8489 27660 8520
rect 27617 8483 27675 8489
rect 27617 8449 27629 8483
rect 27663 8449 27675 8483
rect 27617 8443 27675 8449
rect 24728 8384 25636 8412
rect 24728 8372 24734 8384
rect 25774 8372 25780 8424
rect 25832 8372 25838 8424
rect 26878 8372 26884 8424
rect 26936 8412 26942 8424
rect 27246 8412 27252 8424
rect 26936 8384 27252 8412
rect 26936 8372 26942 8384
rect 27246 8372 27252 8384
rect 27304 8372 27310 8424
rect 27724 8412 27752 8588
rect 27801 8585 27813 8619
rect 27847 8616 27859 8619
rect 28258 8616 28264 8628
rect 27847 8588 28264 8616
rect 27847 8585 27859 8588
rect 27801 8579 27859 8585
rect 28258 8576 28264 8588
rect 28316 8576 28322 8628
rect 28902 8576 28908 8628
rect 28960 8616 28966 8628
rect 28994 8616 29000 8628
rect 28960 8588 29000 8616
rect 28960 8576 28966 8588
rect 28994 8576 29000 8588
rect 29052 8576 29058 8628
rect 32769 8619 32827 8625
rect 29104 8588 29960 8616
rect 28074 8508 28080 8560
rect 28132 8548 28138 8560
rect 28629 8551 28687 8557
rect 28132 8520 28212 8548
rect 28132 8508 28138 8520
rect 28184 8489 28212 8520
rect 28399 8517 28457 8523
rect 28399 8514 28411 8517
rect 28322 8492 28411 8514
rect 28169 8483 28227 8489
rect 28169 8449 28181 8483
rect 28215 8449 28227 8483
rect 28169 8443 28227 8449
rect 28258 8440 28264 8492
rect 28316 8486 28411 8492
rect 28316 8452 28350 8486
rect 28399 8483 28411 8486
rect 28445 8483 28457 8517
rect 28629 8517 28641 8551
rect 28675 8548 28687 8551
rect 29104 8548 29132 8588
rect 28675 8520 29132 8548
rect 29717 8551 29775 8557
rect 28675 8517 28687 8520
rect 28629 8511 28687 8517
rect 29717 8517 29729 8551
rect 29763 8548 29775 8551
rect 29822 8548 29828 8560
rect 29763 8520 29828 8548
rect 29763 8517 29775 8520
rect 29717 8511 29775 8517
rect 28399 8477 28457 8483
rect 28316 8440 28322 8452
rect 28644 8412 28672 8511
rect 29822 8508 29828 8520
rect 29880 8508 29886 8560
rect 29932 8557 29960 8588
rect 32769 8585 32781 8619
rect 32815 8585 32827 8619
rect 32769 8579 32827 8585
rect 29917 8551 29975 8557
rect 29917 8517 29929 8551
rect 29963 8517 29975 8551
rect 29917 8511 29975 8517
rect 28905 8483 28963 8489
rect 28905 8449 28917 8483
rect 28951 8466 28963 8483
rect 28994 8466 29000 8492
rect 28951 8449 29000 8466
rect 28905 8443 29000 8449
rect 28920 8440 29000 8443
rect 29052 8440 29058 8492
rect 29086 8440 29092 8492
rect 29144 8440 29150 8492
rect 29207 8483 29265 8489
rect 29207 8449 29219 8483
rect 29253 8480 29265 8483
rect 29546 8480 29552 8492
rect 29253 8452 29552 8480
rect 29253 8449 29265 8452
rect 29207 8443 29265 8449
rect 29546 8440 29552 8452
rect 29604 8440 29610 8492
rect 28920 8438 29040 8440
rect 28966 8436 29040 8438
rect 27724 8384 28672 8412
rect 24854 8344 24860 8356
rect 23523 8316 24164 8344
rect 24596 8316 24860 8344
rect 23523 8313 23535 8316
rect 23477 8307 23535 8313
rect 20898 8276 20904 8288
rect 20180 8248 20904 8276
rect 14976 8236 14982 8248
rect 20898 8236 20904 8248
rect 20956 8236 20962 8288
rect 21637 8279 21695 8285
rect 21637 8245 21649 8279
rect 21683 8276 21695 8279
rect 23106 8276 23112 8288
rect 21683 8248 23112 8276
rect 21683 8245 21695 8248
rect 21637 8239 21695 8245
rect 23106 8236 23112 8248
rect 23164 8236 23170 8288
rect 23198 8236 23204 8288
rect 23256 8236 23262 8288
rect 23842 8236 23848 8288
rect 23900 8276 23906 8288
rect 24029 8279 24087 8285
rect 24029 8276 24041 8279
rect 23900 8248 24041 8276
rect 23900 8236 23906 8248
rect 24029 8245 24041 8248
rect 24075 8245 24087 8279
rect 24136 8276 24164 8316
rect 24854 8304 24860 8316
rect 24912 8304 24918 8356
rect 25133 8347 25191 8353
rect 25133 8313 25145 8347
rect 25179 8344 25191 8347
rect 25222 8344 25228 8356
rect 25179 8316 25228 8344
rect 25179 8313 25191 8316
rect 25133 8307 25191 8313
rect 25222 8304 25228 8316
rect 25280 8304 25286 8356
rect 25314 8304 25320 8356
rect 25372 8344 25378 8356
rect 27985 8347 28043 8353
rect 27985 8344 27997 8347
rect 25372 8316 25912 8344
rect 25372 8304 25378 8316
rect 24670 8276 24676 8288
rect 24136 8248 24676 8276
rect 24029 8239 24087 8245
rect 24670 8236 24676 8248
rect 24728 8236 24734 8288
rect 24762 8236 24768 8288
rect 24820 8276 24826 8288
rect 25682 8276 25688 8288
rect 24820 8248 25688 8276
rect 24820 8236 24826 8248
rect 25682 8236 25688 8248
rect 25740 8236 25746 8288
rect 25884 8276 25912 8316
rect 26436 8316 27997 8344
rect 26436 8276 26464 8316
rect 27985 8313 27997 8316
rect 28031 8313 28043 8347
rect 27985 8307 28043 8313
rect 28258 8304 28264 8356
rect 28316 8304 28322 8356
rect 28902 8304 28908 8356
rect 28960 8344 28966 8356
rect 29086 8344 29092 8356
rect 28960 8316 29092 8344
rect 28960 8304 28966 8316
rect 29086 8304 29092 8316
rect 29144 8304 29150 8356
rect 29362 8304 29368 8356
rect 29420 8304 29426 8356
rect 29932 8344 29960 8511
rect 30098 8508 30104 8560
rect 30156 8548 30162 8560
rect 30469 8551 30527 8557
rect 30469 8548 30481 8551
rect 30156 8520 30481 8548
rect 30156 8508 30162 8520
rect 30469 8517 30481 8520
rect 30515 8517 30527 8551
rect 30469 8511 30527 8517
rect 30650 8508 30656 8560
rect 30708 8508 30714 8560
rect 30926 8508 30932 8560
rect 30984 8548 30990 8560
rect 30984 8520 32536 8548
rect 30984 8508 30990 8520
rect 30190 8440 30196 8492
rect 30248 8440 30254 8492
rect 30374 8440 30380 8492
rect 30432 8480 30438 8492
rect 30745 8483 30803 8489
rect 30745 8480 30757 8483
rect 30432 8452 30757 8480
rect 30432 8440 30438 8452
rect 30745 8449 30757 8452
rect 30791 8449 30803 8483
rect 30745 8443 30803 8449
rect 30837 8483 30895 8489
rect 30837 8449 30849 8483
rect 30883 8449 30895 8483
rect 30837 8443 30895 8449
rect 30006 8372 30012 8424
rect 30064 8412 30070 8424
rect 30852 8412 30880 8443
rect 31386 8440 31392 8492
rect 31444 8480 31450 8492
rect 31481 8483 31539 8489
rect 31481 8480 31493 8483
rect 31444 8452 31493 8480
rect 31444 8440 31450 8452
rect 31481 8449 31493 8452
rect 31527 8449 31539 8483
rect 31481 8443 31539 8449
rect 31570 8440 31576 8492
rect 31628 8440 31634 8492
rect 31665 8483 31723 8489
rect 31665 8449 31677 8483
rect 31711 8480 31723 8483
rect 31754 8480 31760 8492
rect 31711 8452 31760 8480
rect 31711 8449 31723 8452
rect 31665 8443 31723 8449
rect 31754 8440 31760 8452
rect 31812 8440 31818 8492
rect 32122 8440 32128 8492
rect 32180 8440 32186 8492
rect 32508 8484 32536 8520
rect 32591 8484 32649 8489
rect 32508 8483 32649 8484
rect 32508 8456 32603 8483
rect 32591 8449 32603 8456
rect 32637 8449 32649 8483
rect 32591 8443 32649 8449
rect 31110 8412 31116 8424
rect 30064 8384 30880 8412
rect 30944 8384 31116 8412
rect 30064 8372 30070 8384
rect 30944 8344 30972 8384
rect 31110 8372 31116 8384
rect 31168 8372 31174 8424
rect 31297 8415 31355 8421
rect 31297 8381 31309 8415
rect 31343 8412 31355 8415
rect 32398 8412 32404 8424
rect 31343 8384 32076 8412
rect 31343 8381 31355 8384
rect 31297 8375 31355 8381
rect 29932 8316 30972 8344
rect 31018 8304 31024 8356
rect 31076 8304 31082 8356
rect 31202 8304 31208 8356
rect 31260 8344 31266 8356
rect 31938 8344 31944 8356
rect 31260 8316 31944 8344
rect 31260 8304 31266 8316
rect 31938 8304 31944 8316
rect 31996 8304 32002 8356
rect 25884 8248 26464 8276
rect 26786 8236 26792 8288
rect 26844 8236 26850 8288
rect 27706 8236 27712 8288
rect 27764 8276 27770 8288
rect 28445 8279 28503 8285
rect 28445 8276 28457 8279
rect 27764 8248 28457 8276
rect 27764 8236 27770 8248
rect 28445 8245 28457 8248
rect 28491 8245 28503 8279
rect 28445 8239 28503 8245
rect 28718 8236 28724 8288
rect 28776 8236 28782 8288
rect 29546 8236 29552 8288
rect 29604 8236 29610 8288
rect 29730 8236 29736 8288
rect 29788 8236 29794 8288
rect 29914 8236 29920 8288
rect 29972 8276 29978 8288
rect 30009 8279 30067 8285
rect 30009 8276 30021 8279
rect 29972 8248 30021 8276
rect 29972 8236 29978 8248
rect 30009 8245 30021 8248
rect 30055 8245 30067 8279
rect 30009 8239 30067 8245
rect 31754 8236 31760 8288
rect 31812 8276 31818 8288
rect 31849 8279 31907 8285
rect 31849 8276 31861 8279
rect 31812 8248 31861 8276
rect 31812 8236 31818 8248
rect 31849 8245 31861 8248
rect 31895 8245 31907 8279
rect 32048 8276 32076 8384
rect 32232 8384 32404 8412
rect 32232 8276 32260 8384
rect 32398 8372 32404 8384
rect 32456 8372 32462 8424
rect 32490 8372 32496 8424
rect 32548 8412 32554 8424
rect 32784 8412 32812 8579
rect 32858 8576 32864 8628
rect 32916 8616 32922 8628
rect 33505 8619 33563 8625
rect 32916 8588 32996 8616
rect 32916 8576 32922 8588
rect 32968 8489 32996 8588
rect 33505 8585 33517 8619
rect 33551 8616 33563 8619
rect 34514 8616 34520 8628
rect 33551 8588 34520 8616
rect 33551 8585 33563 8588
rect 33505 8579 33563 8585
rect 34514 8576 34520 8588
rect 34572 8576 34578 8628
rect 34793 8619 34851 8625
rect 34793 8585 34805 8619
rect 34839 8585 34851 8619
rect 35161 8619 35219 8625
rect 35161 8616 35173 8619
rect 34793 8579 34851 8585
rect 35084 8588 35173 8616
rect 33870 8508 33876 8560
rect 33928 8548 33934 8560
rect 34808 8548 34836 8579
rect 33928 8520 34836 8548
rect 33928 8508 33934 8520
rect 32953 8483 33011 8489
rect 32953 8449 32965 8483
rect 32999 8449 33011 8483
rect 32953 8443 33011 8449
rect 33042 8440 33048 8492
rect 33100 8480 33106 8492
rect 33321 8483 33379 8489
rect 33321 8480 33333 8483
rect 33100 8452 33333 8480
rect 33100 8440 33106 8452
rect 33321 8449 33333 8452
rect 33367 8449 33379 8483
rect 33321 8443 33379 8449
rect 33965 8483 34023 8489
rect 33965 8449 33977 8483
rect 34011 8449 34023 8483
rect 33965 8443 34023 8449
rect 32548 8384 32812 8412
rect 32548 8372 32554 8384
rect 33870 8372 33876 8424
rect 33928 8412 33934 8424
rect 33980 8412 34008 8443
rect 34146 8440 34152 8492
rect 34204 8480 34210 8492
rect 34204 8452 34284 8480
rect 34204 8440 34210 8452
rect 33928 8384 34008 8412
rect 34256 8412 34284 8452
rect 34330 8440 34336 8492
rect 34388 8440 34394 8492
rect 34882 8440 34888 8492
rect 34940 8480 34946 8492
rect 34977 8483 35035 8489
rect 34977 8480 34989 8483
rect 34940 8452 34989 8480
rect 34940 8440 34946 8452
rect 34977 8449 34989 8452
rect 35023 8449 35035 8483
rect 34977 8443 35035 8449
rect 35084 8412 35112 8588
rect 35161 8585 35173 8588
rect 35207 8585 35219 8619
rect 35161 8579 35219 8585
rect 35802 8576 35808 8628
rect 35860 8616 35866 8628
rect 36633 8619 36691 8625
rect 36633 8616 36645 8619
rect 35860 8588 36645 8616
rect 35860 8576 35866 8588
rect 36633 8585 36645 8588
rect 36679 8585 36691 8619
rect 36633 8579 36691 8585
rect 36906 8576 36912 8628
rect 36964 8616 36970 8628
rect 37737 8619 37795 8625
rect 37737 8616 37749 8619
rect 36964 8588 37749 8616
rect 36964 8576 36970 8588
rect 37737 8585 37749 8588
rect 37783 8585 37795 8619
rect 37737 8579 37795 8585
rect 38473 8619 38531 8625
rect 38473 8585 38485 8619
rect 38519 8585 38531 8619
rect 38473 8579 38531 8585
rect 37458 8508 37464 8560
rect 37516 8548 37522 8560
rect 38488 8548 38516 8579
rect 37516 8520 38516 8548
rect 37516 8508 37522 8520
rect 38562 8508 38568 8560
rect 38620 8548 38626 8560
rect 38620 8520 39252 8548
rect 38620 8508 38626 8520
rect 35342 8440 35348 8492
rect 35400 8440 35406 8492
rect 35710 8440 35716 8492
rect 35768 8440 35774 8492
rect 35894 8440 35900 8492
rect 35952 8480 35958 8492
rect 36081 8483 36139 8489
rect 36081 8480 36093 8483
rect 35952 8452 36093 8480
rect 35952 8440 35958 8452
rect 36081 8449 36093 8452
rect 36127 8449 36139 8483
rect 36081 8443 36139 8449
rect 36449 8483 36507 8489
rect 36449 8449 36461 8483
rect 36495 8480 36507 8483
rect 36722 8480 36728 8492
rect 36495 8452 36728 8480
rect 36495 8449 36507 8452
rect 36449 8443 36507 8449
rect 36722 8440 36728 8452
rect 36780 8440 36786 8492
rect 36814 8440 36820 8492
rect 36872 8440 36878 8492
rect 37274 8440 37280 8492
rect 37332 8440 37338 8492
rect 37642 8440 37648 8492
rect 37700 8480 37706 8492
rect 37921 8483 37979 8489
rect 37921 8480 37933 8483
rect 37700 8452 37933 8480
rect 37700 8440 37706 8452
rect 37921 8449 37933 8452
rect 37967 8449 37979 8483
rect 37921 8443 37979 8449
rect 38013 8483 38071 8489
rect 38013 8449 38025 8483
rect 38059 8449 38071 8483
rect 38013 8443 38071 8449
rect 38657 8483 38715 8489
rect 38657 8449 38669 8483
rect 38703 8480 38715 8483
rect 38746 8480 38752 8492
rect 38703 8452 38752 8480
rect 38703 8449 38715 8452
rect 38657 8443 38715 8449
rect 34256 8384 35112 8412
rect 33928 8372 33934 8384
rect 35158 8372 35164 8424
rect 35216 8412 35222 8424
rect 35216 8384 35940 8412
rect 35216 8372 35222 8384
rect 32766 8304 32772 8356
rect 32824 8344 32830 8356
rect 33137 8347 33195 8353
rect 33137 8344 33149 8347
rect 32824 8316 33149 8344
rect 32824 8304 32830 8316
rect 33137 8313 33149 8316
rect 33183 8313 33195 8347
rect 33137 8307 33195 8313
rect 33594 8304 33600 8356
rect 33652 8344 33658 8356
rect 34149 8347 34207 8353
rect 34149 8344 34161 8347
rect 33652 8316 34161 8344
rect 33652 8304 33658 8316
rect 34149 8313 34161 8316
rect 34195 8313 34207 8347
rect 34149 8307 34207 8313
rect 34698 8304 34704 8356
rect 34756 8344 34762 8356
rect 35912 8353 35940 8384
rect 37826 8372 37832 8424
rect 37884 8412 37890 8424
rect 38028 8412 38056 8443
rect 38746 8440 38752 8452
rect 38804 8440 38810 8492
rect 38838 8440 38844 8492
rect 38896 8440 38902 8492
rect 39224 8489 39252 8520
rect 39209 8483 39267 8489
rect 39209 8449 39221 8483
rect 39255 8449 39267 8483
rect 39209 8443 39267 8449
rect 37884 8384 38056 8412
rect 37884 8372 37890 8384
rect 35529 8347 35587 8353
rect 35529 8344 35541 8347
rect 34756 8316 35541 8344
rect 34756 8304 34762 8316
rect 35529 8313 35541 8316
rect 35575 8313 35587 8347
rect 35529 8307 35587 8313
rect 35897 8347 35955 8353
rect 35897 8313 35909 8347
rect 35943 8313 35955 8347
rect 35897 8307 35955 8313
rect 36354 8304 36360 8356
rect 36412 8344 36418 8356
rect 36412 8316 37136 8344
rect 36412 8304 36418 8316
rect 32048 8248 32260 8276
rect 32309 8279 32367 8285
rect 31849 8239 31907 8245
rect 32309 8245 32321 8279
rect 32355 8276 32367 8279
rect 32858 8276 32864 8288
rect 32355 8248 32864 8276
rect 32355 8245 32367 8248
rect 32309 8239 32367 8245
rect 32858 8236 32864 8248
rect 32916 8236 32922 8288
rect 33778 8236 33784 8288
rect 33836 8236 33842 8288
rect 35250 8236 35256 8288
rect 35308 8276 35314 8288
rect 36265 8279 36323 8285
rect 36265 8276 36277 8279
rect 35308 8248 36277 8276
rect 35308 8236 35314 8248
rect 36265 8245 36277 8248
rect 36311 8245 36323 8279
rect 37108 8276 37136 8316
rect 37182 8304 37188 8356
rect 37240 8344 37246 8356
rect 38197 8347 38255 8353
rect 38197 8344 38209 8347
rect 37240 8316 38209 8344
rect 37240 8304 37246 8316
rect 38197 8313 38209 8316
rect 38243 8313 38255 8347
rect 38197 8307 38255 8313
rect 39022 8304 39028 8356
rect 39080 8304 39086 8356
rect 39390 8304 39396 8356
rect 39448 8304 39454 8356
rect 37461 8279 37519 8285
rect 37461 8276 37473 8279
rect 37108 8248 37473 8276
rect 36265 8239 36323 8245
rect 37461 8245 37473 8248
rect 37507 8245 37519 8279
rect 37461 8239 37519 8245
rect 1104 8186 39836 8208
rect 1104 8134 1950 8186
rect 2002 8134 2014 8186
rect 2066 8134 2078 8186
rect 2130 8134 2142 8186
rect 2194 8134 2206 8186
rect 2258 8134 7950 8186
rect 8002 8134 8014 8186
rect 8066 8134 8078 8186
rect 8130 8134 8142 8186
rect 8194 8134 8206 8186
rect 8258 8134 13950 8186
rect 14002 8134 14014 8186
rect 14066 8134 14078 8186
rect 14130 8134 14142 8186
rect 14194 8134 14206 8186
rect 14258 8134 19950 8186
rect 20002 8134 20014 8186
rect 20066 8134 20078 8186
rect 20130 8134 20142 8186
rect 20194 8134 20206 8186
rect 20258 8134 25950 8186
rect 26002 8134 26014 8186
rect 26066 8134 26078 8186
rect 26130 8134 26142 8186
rect 26194 8134 26206 8186
rect 26258 8134 31950 8186
rect 32002 8134 32014 8186
rect 32066 8134 32078 8186
rect 32130 8134 32142 8186
rect 32194 8134 32206 8186
rect 32258 8134 37950 8186
rect 38002 8134 38014 8186
rect 38066 8134 38078 8186
rect 38130 8134 38142 8186
rect 38194 8134 38206 8186
rect 38258 8134 39836 8186
rect 1104 8112 39836 8134
rect 3513 8075 3571 8081
rect 3513 8041 3525 8075
rect 3559 8072 3571 8075
rect 3559 8044 4476 8072
rect 3559 8041 3571 8044
rect 3513 8035 3571 8041
rect 4448 8004 4476 8044
rect 4706 8032 4712 8084
rect 4764 8072 4770 8084
rect 4801 8075 4859 8081
rect 4801 8072 4813 8075
rect 4764 8044 4813 8072
rect 4764 8032 4770 8044
rect 4801 8041 4813 8044
rect 4847 8041 4859 8075
rect 4801 8035 4859 8041
rect 6914 8032 6920 8084
rect 6972 8032 6978 8084
rect 7837 8075 7895 8081
rect 7837 8041 7849 8075
rect 7883 8072 7895 8075
rect 11054 8072 11060 8084
rect 7883 8044 11060 8072
rect 7883 8041 7895 8044
rect 7837 8035 7895 8041
rect 11054 8032 11060 8044
rect 11112 8032 11118 8084
rect 11146 8032 11152 8084
rect 11204 8072 11210 8084
rect 12161 8075 12219 8081
rect 12161 8072 12173 8075
rect 11204 8044 12173 8072
rect 11204 8032 11210 8044
rect 12161 8041 12173 8044
rect 12207 8041 12219 8075
rect 12161 8035 12219 8041
rect 12342 8032 12348 8084
rect 12400 8072 12406 8084
rect 16574 8072 16580 8084
rect 12400 8044 16580 8072
rect 12400 8032 12406 8044
rect 16574 8032 16580 8044
rect 16632 8032 16638 8084
rect 16666 8032 16672 8084
rect 16724 8032 16730 8084
rect 17310 8032 17316 8084
rect 17368 8072 17374 8084
rect 18233 8075 18291 8081
rect 18233 8072 18245 8075
rect 17368 8044 18245 8072
rect 17368 8032 17374 8044
rect 18233 8041 18245 8044
rect 18279 8041 18291 8075
rect 18233 8035 18291 8041
rect 18322 8032 18328 8084
rect 18380 8072 18386 8084
rect 18598 8072 18604 8084
rect 18380 8044 18604 8072
rect 18380 8032 18386 8044
rect 18598 8032 18604 8044
rect 18656 8072 18662 8084
rect 20162 8072 20168 8084
rect 18656 8044 20168 8072
rect 18656 8032 18662 8044
rect 20162 8032 20168 8044
rect 20220 8032 20226 8084
rect 22066 8044 24992 8072
rect 4890 8004 4896 8016
rect 4448 7976 4896 8004
rect 4890 7964 4896 7976
rect 4948 7964 4954 8016
rect 6733 8007 6791 8013
rect 5092 7976 5764 8004
rect 1210 7896 1216 7948
rect 1268 7936 1274 7948
rect 2317 7939 2375 7945
rect 2317 7936 2329 7939
rect 1268 7908 2329 7936
rect 1268 7896 1274 7908
rect 2317 7905 2329 7908
rect 2363 7905 2375 7939
rect 2317 7899 2375 7905
rect 750 7828 756 7880
rect 808 7868 814 7880
rect 1397 7871 1455 7877
rect 1397 7868 1409 7871
rect 808 7840 1409 7868
rect 808 7828 814 7840
rect 1397 7837 1409 7840
rect 1443 7837 1455 7871
rect 1397 7831 1455 7837
rect 1673 7871 1731 7877
rect 1673 7837 1685 7871
rect 1719 7868 1731 7871
rect 2406 7868 2412 7880
rect 1719 7840 2412 7868
rect 1719 7837 1731 7840
rect 1673 7831 1731 7837
rect 2406 7828 2412 7840
rect 2464 7828 2470 7880
rect 2590 7828 2596 7880
rect 2648 7828 2654 7880
rect 3329 7871 3387 7877
rect 3329 7868 3341 7871
rect 2746 7840 3341 7868
rect 2498 7760 2504 7812
rect 2556 7800 2562 7812
rect 2746 7800 2774 7840
rect 3329 7837 3341 7840
rect 3375 7837 3387 7871
rect 3329 7831 3387 7837
rect 3789 7871 3847 7877
rect 3789 7837 3801 7871
rect 3835 7837 3847 7871
rect 3789 7831 3847 7837
rect 2556 7772 2774 7800
rect 3804 7800 3832 7831
rect 4062 7828 4068 7880
rect 4120 7828 4126 7880
rect 5092 7868 5120 7976
rect 5166 7896 5172 7948
rect 5224 7936 5230 7948
rect 5736 7945 5764 7976
rect 6733 7973 6745 8007
rect 6779 8004 6791 8007
rect 6779 7976 7512 8004
rect 6779 7973 6791 7976
rect 6733 7967 6791 7973
rect 7484 7945 7512 7976
rect 7650 7964 7656 8016
rect 7708 8004 7714 8016
rect 14277 8007 14335 8013
rect 7708 7976 8248 8004
rect 7708 7964 7714 7976
rect 5445 7939 5503 7945
rect 5445 7936 5457 7939
rect 5224 7908 5457 7936
rect 5224 7896 5230 7908
rect 5445 7905 5457 7908
rect 5491 7905 5503 7939
rect 5445 7899 5503 7905
rect 5721 7939 5779 7945
rect 5721 7905 5733 7939
rect 5767 7905 5779 7939
rect 5721 7899 5779 7905
rect 7469 7939 7527 7945
rect 7469 7905 7481 7939
rect 7515 7905 7527 7939
rect 7926 7936 7932 7948
rect 7469 7899 7527 7905
rect 7668 7908 7932 7936
rect 4724 7840 5120 7868
rect 5261 7871 5319 7877
rect 3878 7800 3884 7812
rect 3804 7772 3884 7800
rect 2556 7760 2562 7772
rect 3878 7760 3884 7772
rect 3936 7800 3942 7812
rect 4724 7800 4752 7840
rect 5261 7837 5273 7871
rect 5307 7868 5319 7871
rect 5626 7868 5632 7880
rect 5307 7840 5632 7868
rect 5307 7837 5319 7840
rect 5261 7831 5319 7837
rect 5626 7828 5632 7840
rect 5684 7828 5690 7880
rect 5902 7828 5908 7880
rect 5960 7868 5966 7880
rect 5997 7871 6055 7877
rect 5997 7868 6009 7871
rect 5960 7840 6009 7868
rect 5960 7828 5966 7840
rect 5997 7837 6009 7840
rect 6043 7837 6055 7871
rect 5997 7831 6055 7837
rect 7285 7871 7343 7877
rect 7285 7837 7297 7871
rect 7331 7868 7343 7871
rect 7668 7868 7696 7908
rect 7926 7896 7932 7908
rect 7984 7896 7990 7948
rect 7331 7840 7696 7868
rect 7331 7837 7343 7840
rect 7285 7831 7343 7837
rect 7742 7828 7748 7880
rect 7800 7868 7806 7880
rect 8021 7871 8079 7877
rect 8021 7868 8033 7871
rect 7800 7840 8033 7868
rect 7800 7828 7806 7840
rect 8021 7837 8033 7840
rect 8067 7837 8079 7871
rect 8021 7831 8079 7837
rect 8110 7828 8116 7880
rect 8168 7828 8174 7880
rect 8220 7868 8248 7976
rect 14277 7973 14289 8007
rect 14323 7973 14335 8007
rect 14277 7967 14335 7973
rect 8757 7939 8815 7945
rect 8757 7905 8769 7939
rect 8803 7905 8815 7939
rect 8757 7899 8815 7905
rect 8297 7871 8355 7877
rect 8297 7868 8309 7871
rect 8220 7840 8309 7868
rect 8297 7837 8309 7840
rect 8343 7837 8355 7871
rect 8297 7831 8355 7837
rect 8386 7828 8392 7880
rect 8444 7828 8450 7880
rect 8527 7871 8585 7877
rect 8527 7837 8539 7871
rect 8573 7868 8585 7871
rect 8772 7868 8800 7899
rect 8938 7896 8944 7948
rect 8996 7896 9002 7948
rect 13446 7896 13452 7948
rect 13504 7936 13510 7948
rect 14292 7936 14320 7967
rect 14642 7964 14648 8016
rect 14700 8004 14706 8016
rect 16485 8007 16543 8013
rect 16485 8004 16497 8007
rect 14700 7976 14780 8004
rect 14700 7964 14706 7976
rect 14752 7936 14780 7976
rect 16132 7976 16497 8004
rect 13504 7908 14228 7936
rect 14292 7908 14688 7936
rect 13504 7896 13510 7908
rect 9208 7871 9266 7877
rect 8573 7837 8596 7868
rect 8772 7865 9168 7868
rect 9208 7865 9220 7871
rect 8772 7840 9220 7865
rect 9140 7837 9220 7840
rect 9254 7837 9266 7871
rect 8527 7831 8596 7837
rect 9208 7831 9266 7837
rect 6638 7800 6644 7812
rect 3936 7772 4752 7800
rect 4816 7772 6644 7800
rect 3936 7760 3942 7772
rect 2774 7692 2780 7744
rect 2832 7732 2838 7744
rect 4816 7732 4844 7772
rect 6638 7760 6644 7772
rect 6696 7760 6702 7812
rect 7300 7772 8248 7800
rect 2832 7704 4844 7732
rect 2832 7692 2838 7704
rect 4890 7692 4896 7744
rect 4948 7692 4954 7744
rect 5353 7735 5411 7741
rect 5353 7701 5365 7735
rect 5399 7732 5411 7735
rect 6546 7732 6552 7744
rect 5399 7704 6552 7732
rect 5399 7701 5411 7704
rect 5353 7695 5411 7701
rect 6546 7692 6552 7704
rect 6604 7732 6610 7744
rect 7300 7732 7328 7772
rect 6604 7704 7328 7732
rect 7377 7735 7435 7741
rect 6604 7692 6610 7704
rect 7377 7701 7389 7735
rect 7423 7732 7435 7735
rect 7742 7732 7748 7744
rect 7423 7704 7748 7732
rect 7423 7701 7435 7704
rect 7377 7695 7435 7701
rect 7742 7692 7748 7704
rect 7800 7692 7806 7744
rect 8220 7732 8248 7772
rect 8568 7732 8596 7831
rect 10502 7828 10508 7880
rect 10560 7828 10566 7880
rect 10594 7828 10600 7880
rect 10652 7868 10658 7880
rect 10689 7871 10747 7877
rect 10689 7868 10701 7871
rect 10652 7840 10701 7868
rect 10652 7828 10658 7840
rect 10689 7837 10701 7840
rect 10735 7837 10747 7871
rect 10689 7831 10747 7837
rect 10781 7871 10839 7877
rect 10781 7837 10793 7871
rect 10827 7868 10839 7871
rect 12345 7871 12403 7877
rect 12345 7868 12357 7871
rect 10827 7840 12357 7868
rect 10827 7837 10839 7840
rect 10781 7831 10839 7837
rect 12345 7837 12357 7840
rect 12391 7868 12403 7871
rect 12434 7868 12440 7880
rect 12391 7840 12440 7868
rect 12391 7837 12403 7840
rect 12345 7831 12403 7837
rect 8938 7760 8944 7812
rect 8996 7800 9002 7812
rect 9674 7800 9680 7812
rect 8996 7772 9680 7800
rect 8996 7760 9002 7772
rect 9674 7760 9680 7772
rect 9732 7800 9738 7812
rect 10796 7800 10824 7831
rect 12434 7828 12440 7840
rect 12492 7828 12498 7880
rect 12618 7877 12624 7880
rect 12612 7868 12624 7877
rect 12579 7840 12624 7868
rect 12612 7831 12624 7840
rect 12618 7828 12624 7831
rect 12676 7828 12682 7880
rect 13170 7828 13176 7880
rect 13228 7868 13234 7880
rect 13722 7868 13728 7880
rect 13228 7840 13728 7868
rect 13228 7828 13234 7840
rect 13722 7828 13728 7840
rect 13780 7828 13786 7880
rect 14093 7871 14151 7877
rect 14093 7837 14105 7871
rect 14139 7837 14151 7871
rect 14200 7868 14228 7908
rect 14660 7880 14688 7908
rect 14752 7908 15240 7936
rect 14277 7871 14335 7877
rect 14277 7868 14289 7871
rect 14200 7840 14289 7868
rect 14093 7831 14151 7837
rect 14277 7837 14289 7840
rect 14323 7837 14335 7871
rect 14277 7831 14335 7837
rect 14369 7871 14427 7877
rect 14369 7837 14381 7871
rect 14415 7837 14427 7871
rect 14369 7831 14427 7837
rect 11054 7809 11060 7812
rect 9732 7772 10824 7800
rect 9732 7760 9738 7772
rect 11048 7763 11060 7809
rect 11054 7760 11060 7763
rect 11112 7760 11118 7812
rect 13906 7800 13912 7812
rect 12360 7772 13912 7800
rect 10318 7732 10324 7744
rect 8220 7704 10324 7732
rect 10318 7692 10324 7704
rect 10376 7692 10382 7744
rect 10689 7735 10747 7741
rect 10689 7701 10701 7735
rect 10735 7732 10747 7735
rect 12360 7732 12388 7772
rect 13906 7760 13912 7772
rect 13964 7760 13970 7812
rect 10735 7704 12388 7732
rect 10735 7701 10747 7704
rect 10689 7695 10747 7701
rect 13722 7692 13728 7744
rect 13780 7692 13786 7744
rect 14108 7732 14136 7831
rect 14182 7760 14188 7812
rect 14240 7800 14246 7812
rect 14384 7800 14412 7831
rect 14458 7828 14464 7880
rect 14516 7868 14522 7880
rect 14553 7871 14611 7877
rect 14553 7868 14565 7871
rect 14516 7840 14565 7868
rect 14516 7828 14522 7840
rect 14553 7837 14565 7840
rect 14599 7837 14611 7871
rect 14553 7831 14611 7837
rect 14642 7828 14648 7880
rect 14700 7828 14706 7880
rect 14752 7877 14780 7908
rect 14737 7871 14795 7877
rect 14737 7837 14749 7871
rect 14783 7837 14795 7871
rect 14737 7831 14795 7837
rect 15102 7828 15108 7880
rect 15160 7828 15166 7880
rect 15212 7868 15240 7908
rect 15746 7868 15752 7880
rect 15212 7840 15752 7868
rect 15746 7828 15752 7840
rect 15804 7868 15810 7880
rect 16132 7868 16160 7976
rect 16485 7973 16497 7976
rect 16531 8004 16543 8007
rect 17034 8004 17040 8016
rect 16531 7976 17040 8004
rect 16531 7973 16543 7976
rect 16485 7967 16543 7973
rect 17034 7964 17040 7976
rect 17092 7964 17098 8016
rect 22066 8004 22094 8044
rect 18432 7976 22094 8004
rect 15804 7840 16160 7868
rect 15804 7828 15810 7840
rect 17402 7828 17408 7880
rect 17460 7868 17466 7880
rect 17782 7871 17840 7877
rect 17782 7868 17794 7871
rect 17460 7840 17794 7868
rect 17460 7828 17466 7840
rect 17782 7837 17794 7840
rect 17828 7837 17840 7871
rect 17782 7831 17840 7837
rect 18046 7828 18052 7880
rect 18104 7828 18110 7880
rect 18432 7877 18460 7976
rect 22370 7964 22376 8016
rect 22428 8004 22434 8016
rect 23014 8004 23020 8016
rect 22428 7976 23020 8004
rect 22428 7964 22434 7976
rect 23014 7964 23020 7976
rect 23072 7964 23078 8016
rect 18506 7896 18512 7948
rect 18564 7936 18570 7948
rect 19889 7939 19947 7945
rect 19889 7936 19901 7939
rect 18564 7908 19901 7936
rect 18564 7896 18570 7908
rect 19889 7905 19901 7908
rect 19935 7936 19947 7939
rect 21450 7936 21456 7948
rect 19935 7908 21456 7936
rect 19935 7905 19947 7908
rect 19889 7899 19947 7905
rect 21450 7896 21456 7908
rect 21508 7896 21514 7948
rect 24578 7936 24584 7948
rect 23952 7908 24584 7936
rect 18417 7871 18475 7877
rect 18417 7837 18429 7871
rect 18463 7837 18475 7871
rect 18417 7831 18475 7837
rect 18598 7828 18604 7880
rect 18656 7828 18662 7880
rect 18693 7871 18751 7877
rect 18693 7837 18705 7871
rect 18739 7837 18751 7871
rect 18693 7831 18751 7837
rect 14240 7772 14412 7800
rect 15013 7803 15071 7809
rect 14240 7760 14246 7772
rect 15013 7769 15025 7803
rect 15059 7800 15071 7803
rect 15350 7803 15408 7809
rect 15350 7800 15362 7803
rect 15059 7772 15362 7800
rect 15059 7769 15071 7772
rect 15013 7763 15071 7769
rect 15350 7769 15362 7772
rect 15396 7769 15408 7803
rect 15350 7763 15408 7769
rect 15838 7760 15844 7812
rect 15896 7800 15902 7812
rect 18708 7800 18736 7831
rect 18874 7828 18880 7880
rect 18932 7828 18938 7880
rect 20254 7828 20260 7880
rect 20312 7868 20318 7880
rect 20441 7871 20499 7877
rect 20441 7868 20453 7871
rect 20312 7840 20453 7868
rect 20312 7828 20318 7840
rect 20441 7837 20453 7840
rect 20487 7837 20499 7871
rect 20441 7831 20499 7837
rect 21910 7828 21916 7880
rect 21968 7868 21974 7880
rect 23952 7868 23980 7908
rect 24578 7896 24584 7908
rect 24636 7896 24642 7948
rect 24964 7936 24992 8044
rect 25038 8032 25044 8084
rect 25096 8072 25102 8084
rect 28902 8072 28908 8084
rect 25096 8044 28908 8072
rect 25096 8032 25102 8044
rect 28902 8032 28908 8044
rect 28960 8032 28966 8084
rect 29549 8075 29607 8081
rect 29549 8041 29561 8075
rect 29595 8072 29607 8075
rect 29730 8072 29736 8084
rect 29595 8044 29736 8072
rect 29595 8041 29607 8044
rect 29549 8035 29607 8041
rect 29730 8032 29736 8044
rect 29788 8032 29794 8084
rect 29822 8032 29828 8084
rect 29880 8072 29886 8084
rect 30190 8072 30196 8084
rect 29880 8044 30196 8072
rect 29880 8032 29886 8044
rect 30190 8032 30196 8044
rect 30248 8032 30254 8084
rect 31202 8072 31208 8084
rect 30300 8044 31208 8072
rect 27798 7964 27804 8016
rect 27856 8004 27862 8016
rect 28445 8007 28503 8013
rect 28445 8004 28457 8007
rect 27856 7976 28457 8004
rect 27856 7964 27862 7976
rect 28445 7973 28457 7976
rect 28491 7973 28503 8007
rect 28445 7967 28503 7973
rect 28718 7964 28724 8016
rect 28776 7964 28782 8016
rect 28828 7976 29040 8004
rect 25038 7936 25044 7948
rect 24964 7908 25044 7936
rect 25038 7896 25044 7908
rect 25096 7896 25102 7948
rect 25498 7896 25504 7948
rect 25556 7936 25562 7948
rect 28077 7939 28135 7945
rect 25556 7908 28019 7936
rect 25556 7896 25562 7908
rect 21968 7840 23980 7868
rect 24029 7871 24087 7877
rect 21968 7828 21974 7840
rect 24029 7837 24041 7871
rect 24075 7868 24087 7871
rect 24118 7868 24124 7880
rect 24075 7840 24124 7868
rect 24075 7837 24087 7840
rect 24029 7831 24087 7837
rect 24118 7828 24124 7840
rect 24176 7868 24182 7880
rect 27062 7868 27068 7880
rect 24176 7840 27068 7868
rect 24176 7828 24182 7840
rect 27062 7828 27068 7840
rect 27120 7868 27126 7880
rect 27522 7868 27528 7880
rect 27120 7840 27528 7868
rect 27120 7828 27126 7840
rect 27522 7828 27528 7840
rect 27580 7868 27586 7880
rect 27893 7871 27951 7877
rect 27893 7868 27905 7871
rect 27580 7840 27905 7868
rect 27580 7828 27586 7840
rect 27893 7837 27905 7840
rect 27939 7837 27951 7871
rect 27991 7868 28019 7908
rect 28077 7905 28089 7939
rect 28123 7936 28135 7939
rect 28828 7936 28856 7976
rect 28123 7908 28856 7936
rect 29012 7936 29040 7976
rect 29178 7964 29184 8016
rect 29236 7964 29242 8016
rect 29362 7964 29368 8016
rect 29420 8004 29426 8016
rect 30300 8004 30328 8044
rect 31202 8032 31208 8044
rect 31260 8032 31266 8084
rect 31570 8032 31576 8084
rect 31628 8072 31634 8084
rect 33042 8072 33048 8084
rect 31628 8044 33048 8072
rect 31628 8032 31634 8044
rect 33042 8032 33048 8044
rect 33100 8032 33106 8084
rect 33410 8032 33416 8084
rect 33468 8072 33474 8084
rect 33873 8075 33931 8081
rect 33873 8072 33885 8075
rect 33468 8044 33885 8072
rect 33468 8032 33474 8044
rect 33873 8041 33885 8044
rect 33919 8041 33931 8075
rect 33873 8035 33931 8041
rect 34514 8032 34520 8084
rect 34572 8072 34578 8084
rect 34793 8075 34851 8081
rect 34793 8072 34805 8075
rect 34572 8044 34805 8072
rect 34572 8032 34578 8044
rect 34793 8041 34805 8044
rect 34839 8041 34851 8075
rect 34793 8035 34851 8041
rect 35526 8032 35532 8084
rect 35584 8072 35590 8084
rect 35713 8075 35771 8081
rect 35713 8072 35725 8075
rect 35584 8044 35725 8072
rect 35584 8032 35590 8044
rect 35713 8041 35725 8044
rect 35759 8041 35771 8075
rect 35713 8035 35771 8041
rect 36078 8032 36084 8084
rect 36136 8072 36142 8084
rect 36265 8075 36323 8081
rect 36265 8072 36277 8075
rect 36136 8044 36277 8072
rect 36136 8032 36142 8044
rect 36265 8041 36277 8044
rect 36311 8041 36323 8075
rect 36265 8035 36323 8041
rect 36630 8032 36636 8084
rect 36688 8072 36694 8084
rect 36817 8075 36875 8081
rect 36817 8072 36829 8075
rect 36688 8044 36829 8072
rect 36688 8032 36694 8044
rect 36817 8041 36829 8044
rect 36863 8041 36875 8075
rect 36817 8035 36875 8041
rect 37734 8032 37740 8084
rect 37792 8072 37798 8084
rect 38013 8075 38071 8081
rect 38013 8072 38025 8075
rect 37792 8044 38025 8072
rect 37792 8032 37798 8044
rect 38013 8041 38025 8044
rect 38059 8041 38071 8075
rect 38013 8035 38071 8041
rect 38654 8032 38660 8084
rect 38712 8032 38718 8084
rect 29420 7976 30328 8004
rect 29420 7964 29426 7976
rect 31754 7964 31760 8016
rect 31812 8004 31818 8016
rect 32490 8004 32496 8016
rect 31812 7976 32496 8004
rect 31812 7964 31818 7976
rect 32490 7964 32496 7976
rect 32548 7964 32554 8016
rect 32766 7964 32772 8016
rect 32824 8004 32830 8016
rect 32824 7976 38884 8004
rect 32824 7964 32830 7976
rect 30466 7936 30472 7948
rect 29012 7908 30472 7936
rect 28123 7905 28135 7908
rect 28077 7899 28135 7905
rect 30466 7896 30472 7908
rect 30524 7896 30530 7948
rect 32309 7939 32367 7945
rect 32309 7936 32321 7939
rect 31496 7908 32321 7936
rect 31496 7880 31524 7908
rect 32309 7905 32321 7908
rect 32355 7905 32367 7939
rect 32309 7899 32367 7905
rect 32953 7939 33011 7945
rect 32953 7905 32965 7939
rect 32999 7936 33011 7939
rect 33137 7939 33195 7945
rect 33137 7936 33149 7939
rect 32999 7908 33149 7936
rect 32999 7905 33011 7908
rect 32953 7899 33011 7905
rect 33137 7905 33149 7908
rect 33183 7905 33195 7939
rect 33137 7899 33195 7905
rect 27991 7840 28295 7868
rect 27893 7831 27951 7837
rect 15896 7772 18736 7800
rect 19061 7803 19119 7809
rect 15896 7760 15902 7772
rect 19061 7769 19073 7803
rect 19107 7800 19119 7803
rect 19334 7800 19340 7812
rect 19107 7772 19340 7800
rect 19107 7769 19119 7772
rect 19061 7763 19119 7769
rect 19334 7760 19340 7772
rect 19392 7760 19398 7812
rect 19426 7760 19432 7812
rect 19484 7800 19490 7812
rect 19484 7772 20116 7800
rect 19484 7760 19490 7772
rect 15470 7732 15476 7744
rect 14108 7704 15476 7732
rect 15470 7692 15476 7704
rect 15528 7692 15534 7744
rect 16574 7692 16580 7744
rect 16632 7732 16638 7744
rect 17954 7732 17960 7744
rect 16632 7704 17960 7732
rect 16632 7692 16638 7704
rect 17954 7692 17960 7704
rect 18012 7692 18018 7744
rect 18966 7692 18972 7744
rect 19024 7732 19030 7744
rect 19245 7735 19303 7741
rect 19245 7732 19257 7735
rect 19024 7704 19257 7732
rect 19024 7692 19030 7704
rect 19245 7701 19257 7704
rect 19291 7701 19303 7735
rect 19245 7695 19303 7701
rect 19794 7692 19800 7744
rect 19852 7732 19858 7744
rect 19981 7735 20039 7741
rect 19981 7732 19993 7735
rect 19852 7704 19993 7732
rect 19852 7692 19858 7704
rect 19981 7701 19993 7704
rect 20027 7701 20039 7735
rect 20088 7732 20116 7772
rect 20162 7760 20168 7812
rect 20220 7760 20226 7812
rect 20346 7760 20352 7812
rect 20404 7760 20410 7812
rect 22554 7760 22560 7812
rect 22612 7800 22618 7812
rect 23762 7803 23820 7809
rect 23762 7800 23774 7803
rect 22612 7772 23774 7800
rect 22612 7760 22618 7772
rect 23762 7769 23774 7772
rect 23808 7769 23820 7803
rect 23762 7763 23820 7769
rect 24486 7760 24492 7812
rect 24544 7760 24550 7812
rect 24946 7760 24952 7812
rect 25004 7800 25010 7812
rect 25866 7800 25872 7812
rect 25004 7772 25872 7800
rect 25004 7760 25010 7772
rect 25866 7760 25872 7772
rect 25924 7760 25930 7812
rect 26234 7760 26240 7812
rect 26292 7760 26298 7812
rect 26329 7803 26387 7809
rect 26329 7769 26341 7803
rect 26375 7769 26387 7803
rect 26329 7763 26387 7769
rect 20990 7732 20996 7744
rect 20088 7704 20996 7732
rect 19981 7695 20039 7701
rect 20990 7692 20996 7704
rect 21048 7692 21054 7744
rect 21082 7692 21088 7744
rect 21140 7732 21146 7744
rect 22649 7735 22707 7741
rect 22649 7732 22661 7735
rect 21140 7704 22661 7732
rect 21140 7692 21146 7704
rect 22649 7701 22661 7704
rect 22695 7701 22707 7735
rect 22649 7695 22707 7701
rect 22738 7692 22744 7744
rect 22796 7732 22802 7744
rect 26344 7732 26372 7763
rect 22796 7704 26372 7732
rect 22796 7692 22802 7704
rect 27982 7692 27988 7744
rect 28040 7732 28046 7744
rect 28169 7735 28227 7741
rect 28169 7732 28181 7735
rect 28040 7704 28181 7732
rect 28040 7692 28046 7704
rect 28169 7701 28181 7704
rect 28215 7701 28227 7735
rect 28267 7732 28295 7840
rect 28350 7828 28356 7880
rect 28408 7828 28414 7880
rect 28442 7828 28448 7880
rect 28500 7868 28506 7880
rect 28629 7871 28687 7877
rect 28629 7868 28641 7871
rect 28500 7840 28641 7868
rect 28500 7828 28506 7840
rect 28629 7837 28641 7840
rect 28675 7837 28687 7871
rect 28629 7831 28687 7837
rect 28902 7828 28908 7880
rect 28960 7828 28966 7880
rect 28997 7871 29055 7877
rect 28997 7837 29009 7871
rect 29043 7837 29055 7871
rect 28997 7831 29055 7837
rect 28810 7760 28816 7812
rect 28868 7800 28874 7812
rect 29012 7800 29040 7831
rect 29638 7828 29644 7880
rect 29696 7868 29702 7880
rect 29733 7871 29791 7877
rect 29733 7868 29745 7871
rect 29696 7840 29745 7868
rect 29696 7828 29702 7840
rect 29733 7837 29745 7840
rect 29779 7837 29791 7871
rect 29733 7831 29791 7837
rect 30009 7871 30067 7877
rect 30009 7837 30021 7871
rect 30055 7868 30067 7871
rect 30285 7871 30343 7877
rect 30285 7868 30297 7871
rect 30055 7840 30297 7868
rect 30055 7837 30067 7840
rect 30009 7831 30067 7837
rect 30285 7837 30297 7840
rect 30331 7837 30343 7871
rect 30285 7831 30343 7837
rect 30377 7871 30435 7877
rect 30377 7837 30389 7871
rect 30423 7868 30435 7871
rect 30558 7868 30564 7880
rect 30423 7840 30564 7868
rect 30423 7837 30435 7840
rect 30377 7831 30435 7837
rect 28868 7772 29040 7800
rect 29748 7800 29776 7831
rect 30101 7803 30159 7809
rect 30101 7800 30113 7803
rect 29748 7772 30113 7800
rect 28868 7760 28874 7772
rect 30101 7769 30113 7772
rect 30147 7769 30159 7803
rect 30300 7800 30328 7831
rect 30558 7828 30564 7840
rect 30616 7828 30622 7880
rect 31478 7868 31484 7880
rect 30668 7840 31484 7868
rect 30668 7800 30696 7840
rect 31478 7828 31484 7840
rect 31536 7828 31542 7880
rect 31754 7868 31760 7880
rect 31588 7840 31760 7868
rect 30300 7772 30696 7800
rect 30736 7803 30794 7809
rect 30101 7763 30159 7769
rect 30736 7769 30748 7803
rect 30782 7800 30794 7803
rect 31588 7800 31616 7840
rect 31754 7828 31760 7840
rect 31812 7828 31818 7880
rect 32214 7828 32220 7880
rect 32272 7828 32278 7880
rect 32582 7828 32588 7880
rect 32640 7868 32646 7880
rect 33045 7871 33103 7877
rect 33045 7868 33057 7871
rect 32640 7840 33057 7868
rect 32640 7828 32646 7840
rect 33045 7837 33057 7840
rect 33091 7837 33103 7871
rect 33045 7831 33103 7837
rect 33226 7828 33232 7880
rect 33284 7868 33290 7880
rect 33321 7871 33379 7877
rect 33321 7868 33333 7871
rect 33284 7840 33333 7868
rect 33284 7828 33290 7840
rect 33321 7837 33333 7840
rect 33367 7837 33379 7871
rect 33321 7831 33379 7837
rect 33502 7828 33508 7880
rect 33560 7868 33566 7880
rect 33781 7871 33839 7877
rect 33781 7868 33793 7871
rect 33560 7840 33793 7868
rect 33560 7828 33566 7840
rect 33781 7837 33793 7840
rect 33827 7837 33839 7871
rect 33781 7831 33839 7837
rect 34057 7871 34115 7877
rect 34057 7837 34069 7871
rect 34103 7837 34115 7871
rect 34057 7831 34115 7837
rect 34977 7871 35035 7877
rect 34977 7837 34989 7871
rect 35023 7837 35035 7871
rect 34977 7831 35035 7837
rect 35897 7871 35955 7877
rect 35897 7837 35909 7871
rect 35943 7868 35955 7871
rect 36354 7868 36360 7880
rect 35943 7840 36360 7868
rect 35943 7837 35955 7840
rect 35897 7831 35955 7837
rect 32600 7800 32628 7828
rect 30782 7772 31616 7800
rect 31680 7772 32628 7800
rect 30782 7769 30794 7772
rect 30736 7763 30794 7769
rect 29362 7732 29368 7744
rect 28267 7704 29368 7732
rect 28169 7695 28227 7701
rect 29362 7692 29368 7704
rect 29420 7692 29426 7744
rect 29917 7735 29975 7741
rect 29917 7701 29929 7735
rect 29963 7732 29975 7735
rect 30558 7732 30564 7744
rect 29963 7704 30564 7732
rect 29963 7701 29975 7704
rect 29917 7695 29975 7701
rect 30558 7692 30564 7704
rect 30616 7732 30622 7744
rect 31386 7732 31392 7744
rect 30616 7704 31392 7732
rect 30616 7692 30622 7704
rect 31386 7692 31392 7704
rect 31444 7732 31450 7744
rect 31680 7732 31708 7772
rect 31864 7741 31892 7772
rect 32766 7760 32772 7812
rect 32824 7800 32830 7812
rect 32950 7800 32956 7812
rect 32824 7772 32956 7800
rect 32824 7760 32830 7772
rect 32950 7760 32956 7772
rect 33008 7760 33014 7812
rect 33686 7760 33692 7812
rect 33744 7800 33750 7812
rect 34072 7800 34100 7831
rect 33744 7772 34100 7800
rect 34992 7800 35020 7831
rect 36354 7828 36360 7840
rect 36412 7828 36418 7880
rect 36446 7828 36452 7880
rect 36504 7828 36510 7880
rect 36998 7828 37004 7880
rect 37056 7828 37062 7880
rect 37366 7828 37372 7880
rect 37424 7868 37430 7880
rect 38856 7877 38884 7976
rect 37829 7871 37887 7877
rect 37829 7868 37841 7871
rect 37424 7840 37841 7868
rect 37424 7828 37430 7840
rect 37829 7837 37841 7840
rect 37875 7837 37887 7871
rect 37829 7831 37887 7837
rect 38473 7871 38531 7877
rect 38473 7837 38485 7871
rect 38519 7837 38531 7871
rect 38473 7831 38531 7837
rect 38841 7871 38899 7877
rect 38841 7837 38853 7871
rect 38887 7837 38899 7871
rect 38841 7831 38899 7837
rect 39209 7871 39267 7877
rect 39209 7837 39221 7871
rect 39255 7868 39267 7871
rect 39298 7868 39304 7880
rect 39255 7840 39304 7868
rect 39255 7837 39267 7840
rect 39209 7831 39267 7837
rect 37550 7800 37556 7812
rect 34992 7772 37556 7800
rect 33744 7760 33750 7772
rect 37550 7760 37556 7772
rect 37608 7760 37614 7812
rect 37734 7760 37740 7812
rect 37792 7800 37798 7812
rect 38488 7800 38516 7831
rect 39298 7828 39304 7840
rect 39356 7828 39362 7880
rect 37792 7772 38516 7800
rect 37792 7760 37798 7772
rect 31444 7704 31708 7732
rect 31849 7735 31907 7741
rect 31444 7692 31450 7704
rect 31849 7701 31861 7735
rect 31895 7701 31907 7735
rect 31849 7695 31907 7701
rect 31938 7692 31944 7744
rect 31996 7732 32002 7744
rect 32033 7735 32091 7741
rect 32033 7732 32045 7735
rect 31996 7704 32045 7732
rect 31996 7692 32002 7704
rect 32033 7701 32045 7704
rect 32079 7701 32091 7735
rect 32033 7695 32091 7701
rect 32122 7692 32128 7744
rect 32180 7732 32186 7744
rect 33505 7735 33563 7741
rect 33505 7732 33517 7735
rect 32180 7704 33517 7732
rect 32180 7692 32186 7704
rect 33505 7701 33517 7704
rect 33551 7701 33563 7735
rect 33505 7695 33563 7701
rect 33594 7692 33600 7744
rect 33652 7692 33658 7744
rect 38930 7692 38936 7744
rect 38988 7732 38994 7744
rect 39025 7735 39083 7741
rect 39025 7732 39037 7735
rect 38988 7704 39037 7732
rect 38988 7692 38994 7704
rect 39025 7701 39037 7704
rect 39071 7701 39083 7735
rect 39025 7695 39083 7701
rect 39390 7692 39396 7744
rect 39448 7692 39454 7744
rect 1104 7642 39836 7664
rect 1104 7590 3010 7642
rect 3062 7590 3074 7642
rect 3126 7590 3138 7642
rect 3190 7590 3202 7642
rect 3254 7590 3266 7642
rect 3318 7590 9010 7642
rect 9062 7590 9074 7642
rect 9126 7590 9138 7642
rect 9190 7590 9202 7642
rect 9254 7590 9266 7642
rect 9318 7590 15010 7642
rect 15062 7590 15074 7642
rect 15126 7590 15138 7642
rect 15190 7590 15202 7642
rect 15254 7590 15266 7642
rect 15318 7590 21010 7642
rect 21062 7590 21074 7642
rect 21126 7590 21138 7642
rect 21190 7590 21202 7642
rect 21254 7590 21266 7642
rect 21318 7590 27010 7642
rect 27062 7590 27074 7642
rect 27126 7590 27138 7642
rect 27190 7590 27202 7642
rect 27254 7590 27266 7642
rect 27318 7590 33010 7642
rect 33062 7590 33074 7642
rect 33126 7590 33138 7642
rect 33190 7590 33202 7642
rect 33254 7590 33266 7642
rect 33318 7590 39010 7642
rect 39062 7590 39074 7642
rect 39126 7590 39138 7642
rect 39190 7590 39202 7642
rect 39254 7590 39266 7642
rect 39318 7590 39836 7642
rect 1104 7568 39836 7590
rect 2498 7488 2504 7540
rect 2556 7488 2562 7540
rect 2682 7488 2688 7540
rect 2740 7488 2746 7540
rect 3145 7531 3203 7537
rect 3145 7497 3157 7531
rect 3191 7528 3203 7531
rect 3418 7528 3424 7540
rect 3191 7500 3424 7528
rect 3191 7497 3203 7500
rect 3145 7491 3203 7497
rect 3418 7488 3424 7500
rect 3476 7488 3482 7540
rect 4982 7488 4988 7540
rect 5040 7488 5046 7540
rect 5166 7488 5172 7540
rect 5224 7488 5230 7540
rect 6641 7531 6699 7537
rect 6641 7497 6653 7531
rect 6687 7528 6699 7531
rect 8846 7528 8852 7540
rect 6687 7500 8852 7528
rect 6687 7497 6699 7500
rect 6641 7491 6699 7497
rect 8846 7488 8852 7500
rect 8904 7488 8910 7540
rect 9490 7488 9496 7540
rect 9548 7528 9554 7540
rect 10594 7528 10600 7540
rect 9548 7500 10600 7528
rect 9548 7488 9554 7500
rect 10594 7488 10600 7500
rect 10652 7488 10658 7540
rect 10870 7488 10876 7540
rect 10928 7528 10934 7540
rect 15930 7528 15936 7540
rect 10928 7500 15936 7528
rect 10928 7488 10934 7500
rect 15930 7488 15936 7500
rect 15988 7488 15994 7540
rect 16574 7488 16580 7540
rect 16632 7528 16638 7540
rect 16879 7531 16937 7537
rect 16879 7528 16891 7531
rect 16632 7500 16891 7528
rect 16632 7488 16638 7500
rect 16879 7497 16891 7500
rect 16925 7528 16937 7531
rect 17862 7528 17868 7540
rect 16925 7500 17868 7528
rect 16925 7497 16937 7500
rect 16879 7491 16937 7497
rect 17862 7488 17868 7500
rect 17920 7488 17926 7540
rect 18506 7488 18512 7540
rect 18564 7488 18570 7540
rect 18598 7488 18604 7540
rect 18656 7528 18662 7540
rect 19610 7528 19616 7540
rect 18656 7500 19616 7528
rect 18656 7488 18662 7500
rect 19610 7488 19616 7500
rect 19668 7488 19674 7540
rect 20165 7531 20223 7537
rect 20165 7497 20177 7531
rect 20211 7528 20223 7531
rect 20211 7500 20484 7528
rect 20211 7497 20223 7500
rect 20165 7491 20223 7497
rect 4890 7460 4896 7472
rect 2332 7432 4896 7460
rect 750 7352 756 7404
rect 808 7392 814 7404
rect 2332 7401 2360 7432
rect 4890 7420 4896 7432
rect 4948 7420 4954 7472
rect 7006 7420 7012 7472
rect 7064 7460 7070 7472
rect 8205 7463 8263 7469
rect 7064 7432 7144 7460
rect 7064 7420 7070 7432
rect 1397 7395 1455 7401
rect 1397 7392 1409 7395
rect 808 7364 1409 7392
rect 808 7352 814 7364
rect 1397 7361 1409 7364
rect 1443 7361 1455 7395
rect 1397 7355 1455 7361
rect 2317 7395 2375 7401
rect 2317 7361 2329 7395
rect 2363 7361 2375 7395
rect 2869 7395 2927 7401
rect 2869 7392 2881 7395
rect 2317 7355 2375 7361
rect 2700 7364 2881 7392
rect 1578 7284 1584 7336
rect 1636 7324 1642 7336
rect 1673 7327 1731 7333
rect 1673 7324 1685 7327
rect 1636 7296 1685 7324
rect 1636 7284 1642 7296
rect 1673 7293 1685 7296
rect 1719 7293 1731 7327
rect 1673 7287 1731 7293
rect 2700 7256 2728 7364
rect 2869 7361 2881 7364
rect 2915 7361 2927 7395
rect 2869 7355 2927 7361
rect 2961 7395 3019 7401
rect 2961 7361 2973 7395
rect 3007 7361 3019 7395
rect 2961 7355 3019 7361
rect 2774 7284 2780 7336
rect 2832 7324 2838 7336
rect 2976 7324 3004 7355
rect 3142 7352 3148 7404
rect 3200 7392 3206 7404
rect 3605 7395 3663 7401
rect 3605 7392 3617 7395
rect 3200 7364 3617 7392
rect 3200 7352 3206 7364
rect 3605 7361 3617 7364
rect 3651 7392 3663 7395
rect 4062 7392 4068 7404
rect 3651 7364 4068 7392
rect 3651 7361 3663 7364
rect 3605 7355 3663 7361
rect 4062 7352 4068 7364
rect 4120 7352 4126 7404
rect 4709 7395 4767 7401
rect 4709 7361 4721 7395
rect 4755 7392 4767 7395
rect 4801 7395 4859 7401
rect 4801 7392 4813 7395
rect 4755 7364 4813 7392
rect 4755 7361 4767 7364
rect 4709 7355 4767 7361
rect 4801 7361 4813 7364
rect 4847 7361 4859 7395
rect 5902 7392 5908 7404
rect 4801 7355 4859 7361
rect 4908 7364 5908 7392
rect 2832 7296 3004 7324
rect 2832 7284 2838 7296
rect 3326 7284 3332 7336
rect 3384 7284 3390 7336
rect 3970 7284 3976 7336
rect 4028 7324 4034 7336
rect 4908 7324 4936 7364
rect 5902 7352 5908 7364
rect 5960 7352 5966 7404
rect 6638 7352 6644 7404
rect 6696 7352 6702 7404
rect 6822 7352 6828 7404
rect 6880 7352 6886 7404
rect 7116 7401 7144 7432
rect 8205 7429 8217 7463
rect 8251 7460 8263 7463
rect 8386 7460 8392 7472
rect 8251 7432 8392 7460
rect 8251 7429 8263 7432
rect 8205 7423 8263 7429
rect 8386 7420 8392 7432
rect 8444 7460 8450 7472
rect 8542 7463 8600 7469
rect 8542 7460 8554 7463
rect 8444 7432 8554 7460
rect 8444 7420 8450 7432
rect 8542 7429 8554 7432
rect 8588 7429 8600 7463
rect 8542 7423 8600 7429
rect 9674 7420 9680 7472
rect 9732 7460 9738 7472
rect 10502 7460 10508 7472
rect 9732 7432 9996 7460
rect 9732 7420 9738 7432
rect 7101 7395 7159 7401
rect 7101 7361 7113 7395
rect 7147 7361 7159 7395
rect 7101 7355 7159 7361
rect 7650 7352 7656 7404
rect 7708 7392 7714 7404
rect 7745 7395 7803 7401
rect 7745 7392 7757 7395
rect 7708 7364 7757 7392
rect 7708 7352 7714 7364
rect 7745 7361 7757 7364
rect 7791 7361 7803 7395
rect 7745 7355 7803 7361
rect 8021 7395 8079 7401
rect 8021 7361 8033 7395
rect 8067 7361 8079 7395
rect 8021 7355 8079 7361
rect 4028 7296 4936 7324
rect 6181 7327 6239 7333
rect 4028 7284 4034 7296
rect 6181 7293 6193 7327
rect 6227 7324 6239 7327
rect 6362 7324 6368 7336
rect 6227 7296 6368 7324
rect 6227 7293 6239 7296
rect 6181 7287 6239 7293
rect 6362 7284 6368 7296
rect 6420 7284 6426 7336
rect 3234 7256 3240 7268
rect 2700 7228 3240 7256
rect 3234 7216 3240 7228
rect 3292 7216 3298 7268
rect 6656 7256 6684 7352
rect 7466 7284 7472 7336
rect 7524 7324 7530 7336
rect 7837 7327 7895 7333
rect 7837 7324 7849 7327
rect 7524 7296 7849 7324
rect 7524 7284 7530 7296
rect 7837 7293 7849 7296
rect 7883 7293 7895 7327
rect 7837 7287 7895 7293
rect 7285 7259 7343 7265
rect 7285 7256 7297 7259
rect 6656 7228 7297 7256
rect 7285 7225 7297 7228
rect 7331 7225 7343 7259
rect 7285 7219 7343 7225
rect 7561 7259 7619 7265
rect 7561 7225 7573 7259
rect 7607 7256 7619 7259
rect 7926 7256 7932 7268
rect 7607 7228 7932 7256
rect 7607 7225 7619 7228
rect 7561 7219 7619 7225
rect 7926 7216 7932 7228
rect 7984 7216 7990 7268
rect 4338 7148 4344 7200
rect 4396 7148 4402 7200
rect 4709 7191 4767 7197
rect 4709 7157 4721 7191
rect 4755 7188 4767 7191
rect 7190 7188 7196 7200
rect 4755 7160 7196 7188
rect 4755 7157 4767 7160
rect 4709 7151 4767 7157
rect 7190 7148 7196 7160
rect 7248 7148 7254 7200
rect 8036 7188 8064 7355
rect 8294 7352 8300 7404
rect 8352 7352 8358 7404
rect 8846 7352 8852 7404
rect 8904 7392 8910 7404
rect 9968 7401 9996 7432
rect 10336 7432 10508 7460
rect 9953 7395 10011 7401
rect 8904 7364 9352 7392
rect 8904 7352 8910 7364
rect 9324 7324 9352 7364
rect 9953 7361 9965 7395
rect 9999 7361 10011 7395
rect 9953 7355 10011 7361
rect 10220 7395 10278 7401
rect 10220 7361 10232 7395
rect 10266 7392 10278 7395
rect 10336 7392 10364 7432
rect 10502 7420 10508 7432
rect 10560 7420 10566 7472
rect 12986 7420 12992 7472
rect 13044 7460 13050 7472
rect 13090 7463 13148 7469
rect 13090 7460 13102 7463
rect 13044 7432 13102 7460
rect 13044 7420 13050 7432
rect 13090 7429 13102 7432
rect 13136 7429 13148 7463
rect 13090 7423 13148 7429
rect 13188 7432 13492 7460
rect 10266 7364 10364 7392
rect 10266 7361 10278 7364
rect 10220 7355 10278 7361
rect 11698 7352 11704 7404
rect 11756 7352 11762 7404
rect 12710 7352 12716 7404
rect 12768 7392 12774 7404
rect 13188 7392 13216 7432
rect 13464 7401 13492 7432
rect 14642 7420 14648 7472
rect 14700 7460 14706 7472
rect 14930 7463 14988 7469
rect 14930 7460 14942 7463
rect 14700 7432 14942 7460
rect 14700 7420 14706 7432
rect 14930 7429 14942 7432
rect 14976 7429 14988 7463
rect 16206 7460 16212 7472
rect 14930 7423 14988 7429
rect 15304 7432 16212 7460
rect 15304 7404 15332 7432
rect 16206 7420 16212 7432
rect 16264 7460 16270 7472
rect 16264 7432 16620 7460
rect 16264 7420 16270 7432
rect 12768 7364 13216 7392
rect 13449 7395 13507 7401
rect 12768 7352 12774 7364
rect 13449 7361 13461 7395
rect 13495 7361 13507 7395
rect 13449 7355 13507 7361
rect 13538 7352 13544 7404
rect 13596 7392 13602 7404
rect 15197 7395 15255 7401
rect 13596 7364 15148 7392
rect 13596 7352 13602 7364
rect 9674 7324 9680 7336
rect 9324 7296 9680 7324
rect 9674 7284 9680 7296
rect 9732 7284 9738 7336
rect 11514 7284 11520 7336
rect 11572 7284 11578 7336
rect 13354 7284 13360 7336
rect 13412 7284 13418 7336
rect 15120 7324 15148 7364
rect 15197 7361 15209 7395
rect 15243 7392 15255 7395
rect 15286 7392 15292 7404
rect 15243 7364 15292 7392
rect 15243 7361 15255 7364
rect 15197 7355 15255 7361
rect 15286 7352 15292 7364
rect 15344 7352 15350 7404
rect 15378 7352 15384 7404
rect 15436 7352 15442 7404
rect 15562 7352 15568 7404
rect 15620 7392 15626 7404
rect 15657 7395 15715 7401
rect 15657 7392 15669 7395
rect 15620 7364 15669 7392
rect 15620 7352 15626 7364
rect 15657 7361 15669 7364
rect 15703 7361 15715 7395
rect 15657 7355 15715 7361
rect 15838 7352 15844 7404
rect 15896 7352 15902 7404
rect 16022 7352 16028 7404
rect 16080 7392 16086 7404
rect 16117 7395 16175 7401
rect 16117 7392 16129 7395
rect 16080 7364 16129 7392
rect 16080 7352 16086 7364
rect 16117 7361 16129 7364
rect 16163 7361 16175 7395
rect 16117 7355 16175 7361
rect 16485 7395 16543 7401
rect 16485 7361 16497 7395
rect 16531 7361 16543 7395
rect 16592 7392 16620 7432
rect 16666 7420 16672 7472
rect 16724 7460 16730 7472
rect 17034 7460 17040 7472
rect 16724 7432 17040 7460
rect 16724 7420 16730 7432
rect 17034 7420 17040 7432
rect 17092 7420 17098 7472
rect 18046 7460 18052 7472
rect 17144 7432 18052 7460
rect 17144 7401 17172 7432
rect 18046 7420 18052 7432
rect 18104 7460 18110 7472
rect 18104 7432 20300 7460
rect 18104 7420 18110 7432
rect 17129 7395 17187 7401
rect 17129 7392 17141 7395
rect 16592 7364 17141 7392
rect 16485 7355 16543 7361
rect 17129 7361 17141 7364
rect 17175 7361 17187 7395
rect 17385 7395 17443 7401
rect 17385 7392 17397 7395
rect 17129 7355 17187 7361
rect 17236 7364 17397 7392
rect 15473 7327 15531 7333
rect 15473 7324 15485 7327
rect 15120 7296 15485 7324
rect 15473 7293 15485 7296
rect 15519 7293 15531 7327
rect 15473 7287 15531 7293
rect 13633 7259 13691 7265
rect 13633 7225 13645 7259
rect 13679 7256 13691 7259
rect 15565 7259 15623 7265
rect 13679 7228 14320 7256
rect 13679 7225 13691 7228
rect 13633 7219 13691 7225
rect 14292 7200 14320 7228
rect 15565 7225 15577 7259
rect 15611 7225 15623 7259
rect 15565 7219 15623 7225
rect 8662 7188 8668 7200
rect 8036 7160 8668 7188
rect 8662 7148 8668 7160
rect 8720 7188 8726 7200
rect 9490 7188 9496 7200
rect 8720 7160 9496 7188
rect 8720 7148 8726 7160
rect 9490 7148 9496 7160
rect 9548 7148 9554 7200
rect 9677 7191 9735 7197
rect 9677 7157 9689 7191
rect 9723 7188 9735 7191
rect 9950 7188 9956 7200
rect 9723 7160 9956 7188
rect 9723 7157 9735 7160
rect 9677 7151 9735 7157
rect 9950 7148 9956 7160
rect 10008 7188 10014 7200
rect 10318 7188 10324 7200
rect 10008 7160 10324 7188
rect 10008 7148 10014 7160
rect 10318 7148 10324 7160
rect 10376 7148 10382 7200
rect 11333 7191 11391 7197
rect 11333 7157 11345 7191
rect 11379 7188 11391 7191
rect 11422 7188 11428 7200
rect 11379 7160 11428 7188
rect 11379 7157 11391 7160
rect 11333 7151 11391 7157
rect 11422 7148 11428 7160
rect 11480 7148 11486 7200
rect 11882 7148 11888 7200
rect 11940 7148 11946 7200
rect 11974 7148 11980 7200
rect 12032 7148 12038 7200
rect 13814 7148 13820 7200
rect 13872 7148 13878 7200
rect 14274 7148 14280 7200
rect 14332 7148 14338 7200
rect 14550 7148 14556 7200
rect 14608 7188 14614 7200
rect 15580 7188 15608 7219
rect 15930 7216 15936 7268
rect 15988 7256 15994 7268
rect 16301 7259 16359 7265
rect 16301 7256 16313 7259
rect 15988 7228 16313 7256
rect 15988 7216 15994 7228
rect 16301 7225 16313 7228
rect 16347 7225 16359 7259
rect 16500 7256 16528 7355
rect 17236 7324 17264 7364
rect 17385 7361 17397 7364
rect 17431 7361 17443 7395
rect 17385 7355 17443 7361
rect 17052 7296 17264 7324
rect 17052 7265 17080 7296
rect 17037 7259 17095 7265
rect 16500 7228 16988 7256
rect 16301 7219 16359 7225
rect 14608 7160 15608 7188
rect 14608 7148 14614 7160
rect 16022 7148 16028 7200
rect 16080 7188 16086 7200
rect 16666 7188 16672 7200
rect 16080 7160 16672 7188
rect 16080 7148 16086 7160
rect 16666 7148 16672 7160
rect 16724 7148 16730 7200
rect 16850 7148 16856 7200
rect 16908 7148 16914 7200
rect 16960 7188 16988 7228
rect 17037 7225 17049 7259
rect 17083 7225 17095 7259
rect 18708 7256 18736 7432
rect 18792 7395 18850 7401
rect 18792 7361 18804 7395
rect 18838 7392 18850 7395
rect 18892 7392 18920 7432
rect 19058 7401 19064 7404
rect 19052 7392 19064 7401
rect 18838 7364 18920 7392
rect 19019 7364 19064 7392
rect 18838 7361 18850 7364
rect 18792 7355 18850 7361
rect 19052 7355 19064 7364
rect 19058 7352 19064 7355
rect 19116 7352 19122 7404
rect 20272 7401 20300 7432
rect 20257 7395 20315 7401
rect 20257 7361 20269 7395
rect 20303 7392 20315 7395
rect 20346 7392 20352 7404
rect 20303 7364 20352 7392
rect 20303 7361 20315 7364
rect 20257 7355 20315 7361
rect 20346 7352 20352 7364
rect 20404 7352 20410 7404
rect 20456 7392 20484 7500
rect 21634 7488 21640 7540
rect 21692 7488 21698 7540
rect 22094 7488 22100 7540
rect 22152 7528 22158 7540
rect 22465 7531 22523 7537
rect 22465 7528 22477 7531
rect 22152 7500 22477 7528
rect 22152 7488 22158 7500
rect 22465 7497 22477 7500
rect 22511 7528 22523 7531
rect 23290 7528 23296 7540
rect 22511 7500 23296 7528
rect 22511 7497 22523 7500
rect 22465 7491 22523 7497
rect 23290 7488 23296 7500
rect 23348 7488 23354 7540
rect 23474 7488 23480 7540
rect 23532 7528 23538 7540
rect 23532 7500 24440 7528
rect 23532 7488 23538 7500
rect 20524 7463 20582 7469
rect 20524 7429 20536 7463
rect 20570 7460 20582 7463
rect 22922 7460 22928 7472
rect 20570 7432 22928 7460
rect 20570 7429 20582 7432
rect 20524 7423 20582 7429
rect 22922 7420 22928 7432
rect 22980 7420 22986 7472
rect 23198 7420 23204 7472
rect 23256 7460 23262 7472
rect 23854 7463 23912 7469
rect 23854 7460 23866 7463
rect 23256 7432 23866 7460
rect 23256 7420 23262 7432
rect 23854 7429 23866 7432
rect 23900 7429 23912 7463
rect 23854 7423 23912 7429
rect 21358 7392 21364 7404
rect 20456 7364 21364 7392
rect 21358 7352 21364 7364
rect 21416 7392 21422 7404
rect 21821 7395 21879 7401
rect 21821 7392 21833 7395
rect 21416 7364 21833 7392
rect 21416 7352 21422 7364
rect 21821 7361 21833 7364
rect 21867 7361 21879 7395
rect 21821 7355 21879 7361
rect 22646 7352 22652 7404
rect 22704 7392 22710 7404
rect 23382 7392 23388 7404
rect 22704 7364 23388 7392
rect 22704 7352 22710 7364
rect 23382 7352 23388 7364
rect 23440 7352 23446 7404
rect 24118 7352 24124 7404
rect 24176 7352 24182 7404
rect 24412 7401 24440 7500
rect 24946 7488 24952 7540
rect 25004 7488 25010 7540
rect 26510 7488 26516 7540
rect 26568 7488 26574 7540
rect 26789 7531 26847 7537
rect 26789 7497 26801 7531
rect 26835 7528 26847 7531
rect 27341 7531 27399 7537
rect 27341 7528 27353 7531
rect 26835 7500 27353 7528
rect 26835 7497 26847 7500
rect 26789 7491 26847 7497
rect 27341 7497 27353 7500
rect 27387 7497 27399 7531
rect 27341 7491 27399 7497
rect 28994 7488 29000 7540
rect 29052 7528 29058 7540
rect 29052 7500 29684 7528
rect 29052 7488 29058 7500
rect 26234 7420 26240 7472
rect 26292 7420 26298 7472
rect 26528 7460 26556 7488
rect 27433 7463 27491 7469
rect 27433 7460 27445 7463
rect 26528 7432 27445 7460
rect 27433 7429 27445 7432
rect 27479 7429 27491 7463
rect 27433 7423 27491 7429
rect 27522 7420 27528 7472
rect 27580 7460 27586 7472
rect 28252 7463 28310 7469
rect 27580 7432 28028 7460
rect 27580 7420 27586 7432
rect 24397 7395 24455 7401
rect 24397 7361 24409 7395
rect 24443 7361 24455 7395
rect 24397 7355 24455 7361
rect 25682 7352 25688 7404
rect 25740 7392 25746 7404
rect 26513 7395 26571 7401
rect 26513 7392 26525 7395
rect 25740 7364 26525 7392
rect 25740 7352 25746 7364
rect 26513 7361 26525 7364
rect 26559 7361 26571 7395
rect 26513 7355 26571 7361
rect 26605 7395 26663 7401
rect 26605 7361 26617 7395
rect 26651 7361 26663 7395
rect 26605 7355 26663 7361
rect 26418 7284 26424 7336
rect 26476 7324 26482 7336
rect 26620 7324 26648 7355
rect 26786 7352 26792 7404
rect 26844 7392 26850 7404
rect 28000 7401 28028 7432
rect 28252 7429 28264 7463
rect 28298 7460 28310 7463
rect 29546 7460 29552 7472
rect 28298 7432 29552 7460
rect 28298 7429 28310 7432
rect 28252 7423 28310 7429
rect 29546 7420 29552 7432
rect 29604 7420 29610 7472
rect 29656 7460 29684 7500
rect 30006 7488 30012 7540
rect 30064 7488 30070 7540
rect 31478 7488 31484 7540
rect 31536 7528 31542 7540
rect 31941 7531 31999 7537
rect 31941 7528 31953 7531
rect 31536 7500 31953 7528
rect 31536 7488 31542 7500
rect 31941 7497 31953 7500
rect 31987 7497 31999 7531
rect 31941 7491 31999 7497
rect 32950 7488 32956 7540
rect 33008 7488 33014 7540
rect 33042 7488 33048 7540
rect 33100 7528 33106 7540
rect 34333 7531 34391 7537
rect 33100 7500 33456 7528
rect 33100 7488 33106 7500
rect 29822 7460 29828 7472
rect 29656 7432 29828 7460
rect 29822 7420 29828 7432
rect 29880 7460 29886 7472
rect 30193 7463 30251 7469
rect 30193 7460 30205 7463
rect 29880 7432 30205 7460
rect 29880 7420 29886 7432
rect 30193 7429 30205 7432
rect 30239 7429 30251 7463
rect 30193 7423 30251 7429
rect 30828 7463 30886 7469
rect 30828 7429 30840 7463
rect 30874 7460 30886 7463
rect 32122 7460 32128 7472
rect 30874 7432 32128 7460
rect 30874 7429 30886 7432
rect 30828 7423 30886 7429
rect 32122 7420 32128 7432
rect 32180 7420 32186 7472
rect 32214 7420 32220 7472
rect 32272 7460 32278 7472
rect 32272 7432 33180 7460
rect 32272 7420 32278 7432
rect 27985 7395 28043 7401
rect 26844 7364 27568 7392
rect 26844 7352 26850 7364
rect 27540 7333 27568 7364
rect 27985 7361 27997 7395
rect 28031 7361 28043 7395
rect 27985 7355 28043 7361
rect 28534 7352 28540 7404
rect 28592 7392 28598 7404
rect 29362 7392 29368 7404
rect 28592 7364 29368 7392
rect 28592 7352 28598 7364
rect 29362 7352 29368 7364
rect 29420 7352 29426 7404
rect 29638 7352 29644 7404
rect 29696 7352 29702 7404
rect 30098 7352 30104 7404
rect 30156 7352 30162 7404
rect 30466 7352 30472 7404
rect 30524 7392 30530 7404
rect 30561 7395 30619 7401
rect 30561 7392 30573 7395
rect 30524 7364 30573 7392
rect 30524 7352 30530 7364
rect 30561 7361 30573 7364
rect 30607 7361 30619 7395
rect 30561 7355 30619 7361
rect 31588 7364 32260 7392
rect 26476 7296 26648 7324
rect 27525 7327 27583 7333
rect 26476 7284 26482 7296
rect 27525 7293 27537 7327
rect 27571 7293 27583 7327
rect 27525 7287 27583 7293
rect 18782 7256 18788 7268
rect 18708 7228 18788 7256
rect 17037 7219 17095 7225
rect 18782 7216 18788 7228
rect 18840 7216 18846 7268
rect 22370 7216 22376 7268
rect 22428 7256 22434 7268
rect 22428 7228 22876 7256
rect 22428 7216 22434 7228
rect 18598 7188 18604 7200
rect 16960 7160 18604 7188
rect 18598 7148 18604 7160
rect 18656 7148 18662 7200
rect 20162 7148 20168 7200
rect 20220 7188 20226 7200
rect 22186 7188 22192 7200
rect 20220 7160 22192 7188
rect 20220 7148 20226 7160
rect 22186 7148 22192 7160
rect 22244 7188 22250 7200
rect 22646 7188 22652 7200
rect 22244 7160 22652 7188
rect 22244 7148 22250 7160
rect 22646 7148 22652 7160
rect 22704 7188 22710 7200
rect 22741 7191 22799 7197
rect 22741 7188 22753 7191
rect 22704 7160 22753 7188
rect 22704 7148 22710 7160
rect 22741 7157 22753 7160
rect 22787 7157 22799 7191
rect 22848 7188 22876 7228
rect 24118 7216 24124 7268
rect 24176 7256 24182 7268
rect 29365 7259 29423 7265
rect 24176 7228 27200 7256
rect 24176 7216 24182 7228
rect 24213 7191 24271 7197
rect 24213 7188 24225 7191
rect 22848 7160 24225 7188
rect 22741 7151 22799 7157
rect 24213 7157 24225 7160
rect 24259 7157 24271 7191
rect 24213 7151 24271 7157
rect 25774 7148 25780 7200
rect 25832 7188 25838 7200
rect 26329 7191 26387 7197
rect 26329 7188 26341 7191
rect 25832 7160 26341 7188
rect 25832 7148 25838 7160
rect 26329 7157 26341 7160
rect 26375 7157 26387 7191
rect 26329 7151 26387 7157
rect 26973 7191 27031 7197
rect 26973 7157 26985 7191
rect 27019 7188 27031 7191
rect 27062 7188 27068 7200
rect 27019 7160 27068 7188
rect 27019 7157 27031 7160
rect 26973 7151 27031 7157
rect 27062 7148 27068 7160
rect 27120 7148 27126 7200
rect 27172 7188 27200 7228
rect 29365 7225 29377 7259
rect 29411 7256 29423 7259
rect 29656 7256 29684 7352
rect 29730 7284 29736 7336
rect 29788 7284 29794 7336
rect 29411 7228 29684 7256
rect 29411 7225 29423 7228
rect 29365 7219 29423 7225
rect 31588 7188 31616 7364
rect 31938 7284 31944 7336
rect 31996 7324 32002 7336
rect 32125 7327 32183 7333
rect 32125 7324 32137 7327
rect 31996 7296 32137 7324
rect 31996 7284 32002 7296
rect 32125 7293 32137 7296
rect 32171 7293 32183 7327
rect 32232 7324 32260 7364
rect 32582 7352 32588 7404
rect 32640 7352 32646 7404
rect 32766 7352 32772 7404
rect 32824 7392 32830 7404
rect 33152 7401 33180 7432
rect 33428 7401 33456 7500
rect 34333 7497 34345 7531
rect 34379 7528 34391 7531
rect 34422 7528 34428 7540
rect 34379 7500 34428 7528
rect 34379 7497 34391 7500
rect 34333 7491 34391 7497
rect 34422 7488 34428 7500
rect 34480 7488 34486 7540
rect 36446 7488 36452 7540
rect 36504 7528 36510 7540
rect 37461 7531 37519 7537
rect 37461 7528 37473 7531
rect 36504 7500 37473 7528
rect 36504 7488 36510 7500
rect 37461 7497 37473 7500
rect 37507 7497 37519 7531
rect 37461 7491 37519 7497
rect 38289 7531 38347 7537
rect 38289 7497 38301 7531
rect 38335 7497 38347 7531
rect 38289 7491 38347 7497
rect 38657 7531 38715 7537
rect 38657 7497 38669 7531
rect 38703 7528 38715 7531
rect 38838 7528 38844 7540
rect 38703 7500 38844 7528
rect 38703 7497 38715 7500
rect 38657 7491 38715 7497
rect 34146 7460 34152 7472
rect 33704 7432 34152 7460
rect 33704 7401 33732 7432
rect 34146 7420 34152 7432
rect 34204 7420 34210 7472
rect 34606 7420 34612 7472
rect 34664 7460 34670 7472
rect 38304 7460 38332 7491
rect 38838 7488 38844 7500
rect 38896 7488 38902 7540
rect 39025 7531 39083 7537
rect 39025 7497 39037 7531
rect 39071 7528 39083 7531
rect 39574 7528 39580 7540
rect 39071 7500 39580 7528
rect 39071 7497 39083 7500
rect 39025 7491 39083 7497
rect 39574 7488 39580 7500
rect 39632 7488 39638 7540
rect 39758 7460 39764 7472
rect 34664 7432 38148 7460
rect 38304 7432 39764 7460
rect 34664 7420 34670 7432
rect 32861 7395 32919 7401
rect 32861 7392 32873 7395
rect 32824 7364 32873 7392
rect 32824 7352 32830 7364
rect 32861 7361 32873 7364
rect 32907 7361 32919 7395
rect 32861 7355 32919 7361
rect 33137 7395 33195 7401
rect 33137 7361 33149 7395
rect 33183 7361 33195 7395
rect 33137 7355 33195 7361
rect 33413 7395 33471 7401
rect 33413 7361 33425 7395
rect 33459 7361 33471 7395
rect 33413 7355 33471 7361
rect 33689 7395 33747 7401
rect 33689 7361 33701 7395
rect 33735 7361 33747 7395
rect 33689 7355 33747 7361
rect 33962 7352 33968 7404
rect 34020 7352 34026 7404
rect 34238 7352 34244 7404
rect 34296 7352 34302 7404
rect 34514 7352 34520 7404
rect 34572 7352 34578 7404
rect 38120 7401 38148 7432
rect 39758 7420 39764 7432
rect 39816 7420 39822 7472
rect 37645 7395 37703 7401
rect 37645 7361 37657 7395
rect 37691 7361 37703 7395
rect 37645 7355 37703 7361
rect 37737 7395 37795 7401
rect 37737 7361 37749 7395
rect 37783 7361 37795 7395
rect 37737 7355 37795 7361
rect 38105 7395 38163 7401
rect 38105 7361 38117 7395
rect 38151 7361 38163 7395
rect 38105 7355 38163 7361
rect 32232 7296 33548 7324
rect 32125 7287 32183 7293
rect 32214 7216 32220 7268
rect 32272 7216 32278 7268
rect 32324 7228 32812 7256
rect 27172 7160 31616 7188
rect 31938 7148 31944 7200
rect 31996 7188 32002 7200
rect 32324 7188 32352 7228
rect 31996 7160 32352 7188
rect 31996 7148 32002 7160
rect 32490 7148 32496 7200
rect 32548 7188 32554 7200
rect 32677 7191 32735 7197
rect 32677 7188 32689 7191
rect 32548 7160 32689 7188
rect 32548 7148 32554 7160
rect 32677 7157 32689 7160
rect 32723 7157 32735 7191
rect 32784 7188 32812 7228
rect 33226 7216 33232 7268
rect 33284 7216 33290 7268
rect 33520 7265 33548 7296
rect 33778 7284 33784 7336
rect 33836 7324 33842 7336
rect 37660 7324 37688 7355
rect 33836 7296 37688 7324
rect 33836 7284 33842 7296
rect 33505 7259 33563 7265
rect 33505 7225 33517 7259
rect 33551 7225 33563 7259
rect 37752 7256 37780 7355
rect 38286 7352 38292 7404
rect 38344 7392 38350 7404
rect 38473 7395 38531 7401
rect 38473 7392 38485 7395
rect 38344 7364 38485 7392
rect 38344 7352 38350 7364
rect 38473 7361 38485 7364
rect 38519 7361 38531 7395
rect 38473 7355 38531 7361
rect 38841 7395 38899 7401
rect 38841 7361 38853 7395
rect 38887 7361 38899 7395
rect 38841 7355 38899 7361
rect 33505 7219 33563 7225
rect 33612 7228 37780 7256
rect 37921 7259 37979 7265
rect 33612 7188 33640 7228
rect 37921 7225 37933 7259
rect 37967 7256 37979 7259
rect 38562 7256 38568 7268
rect 37967 7228 38568 7256
rect 37967 7225 37979 7228
rect 37921 7219 37979 7225
rect 38562 7216 38568 7228
rect 38620 7216 38626 7268
rect 32784 7160 33640 7188
rect 32677 7151 32735 7157
rect 33778 7148 33784 7200
rect 33836 7148 33842 7200
rect 34057 7191 34115 7197
rect 34057 7157 34069 7191
rect 34103 7188 34115 7191
rect 34790 7188 34796 7200
rect 34103 7160 34796 7188
rect 34103 7157 34115 7160
rect 34057 7151 34115 7157
rect 34790 7148 34796 7160
rect 34848 7148 34854 7200
rect 35986 7148 35992 7200
rect 36044 7188 36050 7200
rect 38856 7188 38884 7355
rect 39206 7352 39212 7404
rect 39264 7352 39270 7404
rect 36044 7160 38884 7188
rect 36044 7148 36050 7160
rect 39390 7148 39396 7200
rect 39448 7148 39454 7200
rect 1104 7098 39836 7120
rect 1104 7046 1950 7098
rect 2002 7046 2014 7098
rect 2066 7046 2078 7098
rect 2130 7046 2142 7098
rect 2194 7046 2206 7098
rect 2258 7046 7950 7098
rect 8002 7046 8014 7098
rect 8066 7046 8078 7098
rect 8130 7046 8142 7098
rect 8194 7046 8206 7098
rect 8258 7046 13950 7098
rect 14002 7046 14014 7098
rect 14066 7046 14078 7098
rect 14130 7046 14142 7098
rect 14194 7046 14206 7098
rect 14258 7046 19950 7098
rect 20002 7046 20014 7098
rect 20066 7046 20078 7098
rect 20130 7046 20142 7098
rect 20194 7046 20206 7098
rect 20258 7046 25950 7098
rect 26002 7046 26014 7098
rect 26066 7046 26078 7098
rect 26130 7046 26142 7098
rect 26194 7046 26206 7098
rect 26258 7046 31950 7098
rect 32002 7046 32014 7098
rect 32066 7046 32078 7098
rect 32130 7046 32142 7098
rect 32194 7046 32206 7098
rect 32258 7046 37950 7098
rect 38002 7046 38014 7098
rect 38066 7046 38078 7098
rect 38130 7046 38142 7098
rect 38194 7046 38206 7098
rect 38258 7046 39836 7098
rect 1104 7024 39836 7046
rect 2777 6987 2835 6993
rect 2777 6953 2789 6987
rect 2823 6984 2835 6987
rect 3602 6984 3608 6996
rect 2823 6956 3608 6984
rect 2823 6953 2835 6956
rect 2777 6947 2835 6953
rect 3602 6944 3608 6956
rect 3660 6944 3666 6996
rect 3878 6944 3884 6996
rect 3936 6984 3942 6996
rect 5442 6984 5448 6996
rect 3936 6956 5448 6984
rect 3936 6944 3942 6956
rect 5442 6944 5448 6956
rect 5500 6944 5506 6996
rect 7377 6987 7435 6993
rect 7377 6984 7389 6987
rect 5552 6956 7389 6984
rect 2409 6919 2467 6925
rect 2409 6916 2421 6919
rect 1780 6888 2421 6916
rect 1394 6808 1400 6860
rect 1452 6848 1458 6860
rect 1780 6848 1808 6888
rect 2409 6885 2421 6888
rect 2455 6885 2467 6919
rect 2409 6879 2467 6885
rect 3234 6876 3240 6928
rect 3292 6916 3298 6928
rect 3292 6888 3372 6916
rect 3292 6876 3298 6888
rect 3142 6848 3148 6860
rect 1452 6820 1808 6848
rect 1872 6820 3148 6848
rect 1452 6808 1458 6820
rect 1670 6672 1676 6724
rect 1728 6712 1734 6724
rect 1872 6712 1900 6820
rect 3142 6808 3148 6820
rect 3200 6808 3206 6860
rect 1949 6783 2007 6789
rect 1949 6749 1961 6783
rect 1995 6780 2007 6783
rect 2501 6783 2559 6789
rect 1995 6752 2360 6780
rect 1995 6749 2007 6752
rect 1949 6743 2007 6749
rect 2133 6715 2191 6721
rect 2133 6712 2145 6715
rect 1728 6684 2145 6712
rect 1728 6672 1734 6684
rect 2133 6681 2145 6684
rect 2179 6681 2191 6715
rect 2332 6712 2360 6752
rect 2501 6749 2513 6783
rect 2547 6780 2559 6783
rect 2593 6783 2651 6789
rect 2593 6780 2605 6783
rect 2547 6752 2605 6780
rect 2547 6749 2559 6752
rect 2501 6743 2559 6749
rect 2593 6749 2605 6752
rect 2639 6749 2651 6783
rect 2593 6743 2651 6749
rect 3234 6740 3240 6792
rect 3292 6740 3298 6792
rect 3344 6780 3372 6888
rect 4062 6876 4068 6928
rect 4120 6916 4126 6928
rect 4246 6916 4252 6928
rect 4120 6888 4252 6916
rect 4120 6876 4126 6888
rect 4246 6876 4252 6888
rect 4304 6876 4310 6928
rect 4338 6876 4344 6928
rect 4396 6916 4402 6928
rect 5552 6916 5580 6956
rect 7377 6953 7389 6956
rect 7423 6953 7435 6987
rect 7377 6947 7435 6953
rect 7742 6944 7748 6996
rect 7800 6984 7806 6996
rect 7800 6956 11008 6984
rect 7800 6944 7806 6956
rect 4396 6888 4476 6916
rect 4396 6876 4402 6888
rect 3510 6808 3516 6860
rect 3568 6848 3574 6860
rect 4448 6857 4476 6888
rect 5092 6888 5580 6916
rect 6457 6919 6515 6925
rect 4433 6851 4491 6857
rect 3568 6820 4384 6848
rect 3568 6808 3574 6820
rect 3605 6783 3663 6789
rect 3605 6780 3617 6783
rect 3344 6752 3617 6780
rect 3605 6749 3617 6752
rect 3651 6749 3663 6783
rect 3605 6743 3663 6749
rect 4246 6740 4252 6792
rect 4304 6740 4310 6792
rect 4356 6789 4384 6820
rect 4433 6817 4445 6851
rect 4479 6817 4491 6851
rect 5092 6848 5120 6888
rect 6457 6885 6469 6919
rect 6503 6916 6515 6919
rect 6503 6888 7144 6916
rect 6503 6885 6515 6888
rect 6457 6879 6515 6885
rect 4433 6811 4491 6817
rect 4908 6820 5120 6848
rect 4341 6783 4399 6789
rect 4341 6749 4353 6783
rect 4387 6780 4399 6783
rect 4908 6780 4936 6820
rect 5166 6808 5172 6860
rect 5224 6808 5230 6860
rect 6546 6808 6552 6860
rect 6604 6848 6610 6860
rect 7116 6857 7144 6888
rect 8846 6876 8852 6928
rect 8904 6876 8910 6928
rect 10870 6916 10876 6928
rect 9968 6888 10876 6916
rect 7009 6851 7067 6857
rect 7009 6848 7021 6851
rect 6604 6820 7021 6848
rect 6604 6808 6610 6820
rect 7009 6817 7021 6820
rect 7055 6817 7067 6851
rect 7009 6811 7067 6817
rect 7101 6851 7159 6857
rect 7101 6817 7113 6851
rect 7147 6817 7159 6851
rect 8864 6848 8892 6876
rect 7101 6811 7159 6817
rect 8671 6820 8892 6848
rect 4387 6752 4936 6780
rect 4387 6749 4399 6752
rect 4341 6743 4399 6749
rect 4982 6740 4988 6792
rect 5040 6740 5046 6792
rect 5184 6780 5212 6808
rect 5353 6783 5411 6789
rect 5353 6780 5365 6783
rect 5184 6752 5365 6780
rect 5353 6749 5365 6752
rect 5399 6749 5411 6783
rect 5353 6743 5411 6749
rect 5442 6740 5448 6792
rect 5500 6740 5506 6792
rect 5721 6783 5779 6789
rect 5721 6749 5733 6783
rect 5767 6780 5779 6783
rect 5810 6780 5816 6792
rect 5767 6752 5816 6780
rect 5767 6749 5779 6752
rect 5721 6743 5779 6749
rect 5810 6740 5816 6752
rect 5868 6740 5874 6792
rect 6914 6740 6920 6792
rect 6972 6740 6978 6792
rect 8671 6780 8699 6820
rect 7300 6752 8699 6780
rect 8757 6783 8815 6789
rect 6822 6712 6828 6724
rect 2332 6684 4200 6712
rect 2133 6675 2191 6681
rect 1762 6604 1768 6656
rect 1820 6604 1826 6656
rect 2222 6604 2228 6656
rect 2280 6604 2286 6656
rect 3053 6647 3111 6653
rect 3053 6613 3065 6647
rect 3099 6644 3111 6647
rect 3326 6644 3332 6656
rect 3099 6616 3332 6644
rect 3099 6613 3111 6616
rect 3053 6607 3111 6613
rect 3326 6604 3332 6616
rect 3384 6604 3390 6656
rect 3421 6647 3479 6653
rect 3421 6613 3433 6647
rect 3467 6644 3479 6647
rect 3786 6644 3792 6656
rect 3467 6616 3792 6644
rect 3467 6613 3479 6616
rect 3421 6607 3479 6613
rect 3786 6604 3792 6616
rect 3844 6604 3850 6656
rect 3878 6604 3884 6656
rect 3936 6604 3942 6656
rect 4172 6644 4200 6684
rect 4264 6684 6828 6712
rect 4264 6644 4292 6684
rect 6822 6672 6828 6684
rect 6880 6672 6886 6724
rect 4172 6616 4292 6644
rect 4706 6604 4712 6656
rect 4764 6644 4770 6656
rect 4801 6647 4859 6653
rect 4801 6644 4813 6647
rect 4764 6616 4813 6644
rect 4764 6604 4770 6616
rect 4801 6613 4813 6616
rect 4847 6613 4859 6647
rect 4801 6607 4859 6613
rect 5166 6604 5172 6656
rect 5224 6604 5230 6656
rect 5258 6604 5264 6656
rect 5316 6644 5322 6656
rect 6549 6647 6607 6653
rect 6549 6644 6561 6647
rect 5316 6616 6561 6644
rect 5316 6604 5322 6616
rect 6549 6613 6561 6616
rect 6595 6613 6607 6647
rect 6549 6607 6607 6613
rect 6914 6604 6920 6656
rect 6972 6644 6978 6656
rect 7300 6644 7328 6752
rect 8757 6749 8769 6783
rect 8803 6780 8815 6783
rect 8846 6780 8852 6792
rect 8803 6752 8852 6780
rect 8803 6749 8815 6752
rect 8757 6743 8815 6749
rect 8846 6740 8852 6752
rect 8904 6780 8910 6792
rect 8941 6783 8999 6789
rect 8941 6780 8953 6783
rect 8904 6752 8953 6780
rect 8904 6740 8910 6752
rect 8941 6749 8953 6752
rect 8987 6780 8999 6783
rect 9582 6780 9588 6792
rect 8987 6752 9588 6780
rect 8987 6749 8999 6752
rect 8941 6743 8999 6749
rect 9582 6740 9588 6752
rect 9640 6740 9646 6792
rect 9674 6740 9680 6792
rect 9732 6780 9738 6792
rect 9968 6780 9996 6888
rect 10870 6876 10876 6888
rect 10928 6876 10934 6928
rect 10980 6916 11008 6956
rect 11054 6944 11060 6996
rect 11112 6944 11118 6996
rect 11149 6987 11207 6993
rect 11149 6953 11161 6987
rect 11195 6984 11207 6987
rect 11698 6984 11704 6996
rect 11195 6956 11704 6984
rect 11195 6953 11207 6956
rect 11149 6947 11207 6953
rect 11698 6944 11704 6956
rect 11756 6944 11762 6996
rect 12345 6987 12403 6993
rect 12345 6953 12357 6987
rect 12391 6984 12403 6987
rect 12434 6984 12440 6996
rect 12391 6956 12440 6984
rect 12391 6953 12403 6956
rect 12345 6947 12403 6953
rect 12434 6944 12440 6956
rect 12492 6984 12498 6996
rect 13354 6984 13360 6996
rect 12492 6956 13360 6984
rect 12492 6944 12498 6956
rect 13354 6944 13360 6956
rect 13412 6984 13418 6996
rect 13412 6956 15608 6984
rect 13412 6944 13418 6956
rect 10980 6888 12112 6916
rect 10428 6820 11284 6848
rect 10428 6789 10456 6820
rect 9732 6752 9996 6780
rect 10413 6783 10471 6789
rect 9732 6740 9738 6752
rect 10413 6749 10425 6783
rect 10459 6749 10471 6783
rect 10413 6743 10471 6749
rect 7742 6712 7748 6724
rect 7392 6684 7748 6712
rect 7392 6653 7420 6684
rect 7742 6672 7748 6684
rect 7800 6672 7806 6724
rect 8110 6672 8116 6724
rect 8168 6712 8174 6724
rect 8490 6715 8548 6721
rect 8490 6712 8502 6715
rect 8168 6684 8502 6712
rect 8168 6672 8174 6684
rect 8490 6681 8502 6684
rect 8536 6681 8548 6715
rect 8490 6675 8548 6681
rect 8662 6672 8668 6724
rect 8720 6712 8726 6724
rect 9186 6715 9244 6721
rect 9186 6712 9198 6715
rect 8720 6684 9198 6712
rect 8720 6672 8726 6684
rect 9186 6681 9198 6684
rect 9232 6681 9244 6715
rect 10428 6712 10456 6743
rect 10594 6740 10600 6792
rect 10652 6740 10658 6792
rect 10686 6740 10692 6792
rect 10744 6740 10750 6792
rect 10781 6783 10839 6789
rect 10781 6749 10793 6783
rect 10827 6780 10839 6783
rect 11146 6780 11152 6792
rect 10827 6752 11152 6780
rect 10827 6749 10839 6752
rect 10781 6743 10839 6749
rect 11146 6740 11152 6752
rect 11204 6740 11210 6792
rect 11256 6780 11284 6820
rect 11330 6808 11336 6860
rect 11388 6848 11394 6860
rect 11793 6851 11851 6857
rect 11793 6848 11805 6851
rect 11388 6820 11805 6848
rect 11388 6808 11394 6820
rect 11793 6817 11805 6820
rect 11839 6848 11851 6851
rect 11974 6848 11980 6860
rect 11839 6820 11980 6848
rect 11839 6817 11851 6820
rect 11793 6811 11851 6817
rect 11974 6808 11980 6820
rect 12032 6808 12038 6860
rect 12084 6848 12112 6888
rect 12802 6876 12808 6928
rect 12860 6876 12866 6928
rect 13630 6876 13636 6928
rect 13688 6916 13694 6928
rect 13725 6919 13783 6925
rect 13725 6916 13737 6919
rect 13688 6888 13737 6916
rect 13688 6876 13694 6888
rect 13725 6885 13737 6888
rect 13771 6885 13783 6919
rect 13725 6879 13783 6885
rect 12820 6848 12848 6876
rect 14550 6848 14556 6860
rect 12084 6820 12848 6848
rect 13740 6820 14556 6848
rect 12342 6780 12348 6792
rect 11256 6752 12348 6780
rect 12342 6740 12348 6752
rect 12400 6740 12406 6792
rect 12802 6740 12808 6792
rect 12860 6780 12866 6792
rect 13740 6789 13768 6820
rect 14550 6808 14556 6820
rect 14608 6808 14614 6860
rect 15580 6857 15608 6956
rect 18230 6944 18236 6996
rect 18288 6984 18294 6996
rect 18601 6987 18659 6993
rect 18601 6984 18613 6987
rect 18288 6956 18613 6984
rect 18288 6944 18294 6956
rect 18601 6953 18613 6956
rect 18647 6953 18659 6987
rect 18877 6987 18935 6993
rect 18877 6984 18889 6987
rect 18601 6947 18659 6953
rect 18708 6956 18889 6984
rect 18049 6919 18107 6925
rect 18049 6916 18061 6919
rect 17236 6888 17540 6916
rect 15565 6851 15623 6857
rect 15565 6817 15577 6851
rect 15611 6817 15623 6851
rect 15565 6811 15623 6817
rect 15654 6808 15660 6860
rect 15712 6808 15718 6860
rect 16577 6851 16635 6857
rect 16577 6817 16589 6851
rect 16623 6848 16635 6851
rect 17236 6848 17264 6888
rect 16623 6820 17264 6848
rect 16623 6817 16635 6820
rect 16577 6811 16635 6817
rect 17310 6808 17316 6860
rect 17368 6848 17374 6860
rect 17405 6851 17463 6857
rect 17405 6848 17417 6851
rect 17368 6820 17417 6848
rect 17368 6808 17374 6820
rect 17405 6817 17417 6820
rect 17451 6817 17463 6851
rect 17512 6848 17540 6888
rect 17696 6888 18061 6916
rect 17586 6848 17592 6860
rect 17512 6820 17592 6848
rect 17405 6811 17463 6817
rect 17586 6808 17592 6820
rect 17644 6808 17650 6860
rect 13725 6783 13783 6789
rect 13725 6780 13737 6783
rect 12860 6752 13737 6780
rect 12860 6740 12866 6752
rect 13725 6749 13737 6752
rect 13771 6749 13783 6783
rect 13725 6743 13783 6749
rect 13906 6740 13912 6792
rect 13964 6740 13970 6792
rect 15120 6752 15608 6780
rect 9186 6675 9244 6681
rect 9324 6684 10456 6712
rect 6972 6616 7328 6644
rect 7377 6647 7435 6653
rect 6972 6604 6978 6616
rect 7377 6613 7389 6647
rect 7423 6613 7435 6647
rect 7377 6607 7435 6613
rect 7650 6604 7656 6656
rect 7708 6644 7714 6656
rect 9324 6644 9352 6684
rect 10870 6672 10876 6724
rect 10928 6712 10934 6724
rect 12158 6712 12164 6724
rect 10928 6684 12164 6712
rect 10928 6672 10934 6684
rect 12158 6672 12164 6684
rect 12216 6672 12222 6724
rect 13630 6672 13636 6724
rect 13688 6712 13694 6724
rect 15120 6712 15148 6752
rect 13688 6684 15148 6712
rect 15320 6715 15378 6721
rect 13688 6672 13694 6684
rect 15320 6681 15332 6715
rect 15366 6712 15378 6715
rect 15470 6712 15476 6724
rect 15366 6684 15476 6712
rect 15366 6681 15378 6684
rect 15320 6675 15378 6681
rect 15470 6672 15476 6684
rect 15528 6672 15534 6724
rect 15580 6712 15608 6752
rect 16666 6740 16672 6792
rect 16724 6740 16730 6792
rect 17218 6740 17224 6792
rect 17276 6740 17282 6792
rect 17494 6740 17500 6792
rect 17552 6780 17558 6792
rect 17696 6780 17724 6888
rect 18049 6885 18061 6888
rect 18095 6885 18107 6919
rect 18049 6879 18107 6885
rect 18138 6876 18144 6928
rect 18196 6876 18202 6928
rect 18506 6876 18512 6928
rect 18564 6916 18570 6928
rect 18708 6916 18736 6956
rect 18877 6953 18889 6956
rect 18923 6953 18935 6987
rect 18877 6947 18935 6953
rect 22278 6944 22284 6996
rect 22336 6984 22342 6996
rect 23566 6984 23572 6996
rect 22336 6956 23572 6984
rect 22336 6944 22342 6956
rect 23566 6944 23572 6956
rect 23624 6944 23630 6996
rect 23661 6987 23719 6993
rect 23661 6953 23673 6987
rect 23707 6984 23719 6987
rect 25406 6984 25412 6996
rect 23707 6956 25412 6984
rect 23707 6953 23719 6956
rect 23661 6947 23719 6953
rect 25406 6944 25412 6956
rect 25464 6944 25470 6996
rect 26694 6944 26700 6996
rect 26752 6984 26758 6996
rect 29089 6987 29147 6993
rect 26752 6956 29040 6984
rect 26752 6944 26758 6956
rect 19058 6916 19064 6928
rect 18564 6888 18736 6916
rect 18800 6888 19064 6916
rect 18564 6876 18570 6888
rect 18230 6808 18236 6860
rect 18288 6808 18294 6860
rect 18417 6851 18475 6857
rect 18417 6817 18429 6851
rect 18463 6848 18475 6851
rect 18598 6848 18604 6860
rect 18463 6820 18604 6848
rect 18463 6817 18475 6820
rect 18417 6811 18475 6817
rect 18598 6808 18604 6820
rect 18656 6808 18662 6860
rect 18800 6805 18828 6888
rect 19058 6876 19064 6888
rect 19116 6876 19122 6928
rect 22002 6876 22008 6928
rect 22060 6916 22066 6928
rect 22060 6888 22508 6916
rect 22060 6876 22066 6888
rect 19337 6851 19395 6857
rect 19337 6848 19349 6851
rect 18984 6820 19349 6848
rect 18785 6799 18843 6805
rect 17552 6752 17724 6780
rect 17552 6740 17558 6752
rect 17954 6740 17960 6792
rect 18012 6780 18018 6792
rect 18130 6783 18188 6789
rect 18130 6780 18142 6783
rect 18012 6752 18142 6780
rect 18012 6740 18018 6752
rect 18130 6749 18142 6752
rect 18176 6749 18188 6783
rect 18785 6765 18797 6799
rect 18831 6765 18843 6799
rect 18785 6759 18843 6765
rect 18130 6743 18188 6749
rect 15580 6684 17816 6712
rect 7708 6616 9352 6644
rect 7708 6604 7714 6616
rect 10134 6604 10140 6656
rect 10192 6644 10198 6656
rect 10321 6647 10379 6653
rect 10321 6644 10333 6647
rect 10192 6616 10333 6644
rect 10192 6604 10198 6616
rect 10321 6613 10333 6616
rect 10367 6613 10379 6647
rect 10321 6607 10379 6613
rect 10594 6604 10600 6656
rect 10652 6644 10658 6656
rect 11149 6647 11207 6653
rect 11149 6644 11161 6647
rect 10652 6616 11161 6644
rect 10652 6604 10658 6616
rect 11149 6613 11161 6616
rect 11195 6613 11207 6647
rect 11149 6607 11207 6613
rect 11238 6604 11244 6656
rect 11296 6644 11302 6656
rect 13538 6644 13544 6656
rect 11296 6616 13544 6644
rect 11296 6604 11302 6616
rect 13538 6604 13544 6616
rect 13596 6604 13602 6656
rect 14182 6604 14188 6656
rect 14240 6604 14246 6656
rect 14274 6604 14280 6656
rect 14332 6644 14338 6656
rect 15654 6644 15660 6656
rect 14332 6616 15660 6644
rect 14332 6604 14338 6616
rect 15654 6604 15660 6616
rect 15712 6604 15718 6656
rect 16022 6604 16028 6656
rect 16080 6644 16086 6656
rect 16301 6647 16359 6653
rect 16301 6644 16313 6647
rect 16080 6616 16313 6644
rect 16080 6604 16086 6616
rect 16301 6613 16313 6616
rect 16347 6613 16359 6647
rect 16301 6607 16359 6613
rect 16758 6604 16764 6656
rect 16816 6644 16822 6656
rect 16853 6647 16911 6653
rect 16853 6644 16865 6647
rect 16816 6616 16865 6644
rect 16816 6604 16822 6616
rect 16853 6613 16865 6616
rect 16899 6613 16911 6647
rect 16853 6607 16911 6613
rect 17037 6647 17095 6653
rect 17037 6613 17049 6647
rect 17083 6644 17095 6647
rect 17126 6644 17132 6656
rect 17083 6616 17132 6644
rect 17083 6613 17095 6616
rect 17037 6607 17095 6613
rect 17126 6604 17132 6616
rect 17184 6604 17190 6656
rect 17218 6604 17224 6656
rect 17276 6644 17282 6656
rect 17589 6647 17647 6653
rect 17589 6644 17601 6647
rect 17276 6616 17601 6644
rect 17276 6604 17282 6616
rect 17589 6613 17601 6616
rect 17635 6613 17647 6647
rect 17589 6607 17647 6613
rect 17678 6604 17684 6656
rect 17736 6604 17742 6656
rect 17788 6644 17816 6684
rect 17862 6672 17868 6724
rect 17920 6712 17926 6724
rect 18984 6712 19012 6820
rect 19337 6817 19349 6820
rect 19383 6817 19395 6851
rect 19337 6811 19395 6817
rect 19052 6783 19110 6789
rect 19052 6749 19064 6783
rect 19098 6777 19110 6783
rect 19150 6777 19156 6792
rect 19098 6749 19156 6777
rect 19052 6743 19110 6749
rect 19150 6740 19156 6749
rect 19208 6740 19214 6792
rect 19352 6780 19380 6811
rect 20346 6808 20352 6860
rect 20404 6848 20410 6860
rect 20441 6851 20499 6857
rect 20441 6848 20453 6851
rect 20404 6820 20453 6848
rect 20404 6808 20410 6820
rect 20441 6817 20453 6820
rect 20487 6817 20499 6851
rect 20441 6811 20499 6817
rect 22278 6808 22284 6860
rect 22336 6848 22342 6860
rect 22373 6851 22431 6857
rect 22373 6848 22385 6851
rect 22336 6820 22385 6848
rect 22336 6808 22342 6820
rect 22373 6817 22385 6820
rect 22419 6817 22431 6851
rect 22480 6848 22508 6888
rect 23842 6876 23848 6928
rect 23900 6916 23906 6928
rect 24029 6919 24087 6925
rect 24029 6916 24041 6919
rect 23900 6888 24041 6916
rect 23900 6876 23906 6888
rect 24029 6885 24041 6888
rect 24075 6885 24087 6919
rect 24029 6879 24087 6885
rect 25777 6919 25835 6925
rect 25777 6885 25789 6919
rect 25823 6885 25835 6919
rect 25777 6879 25835 6885
rect 25792 6848 25820 6879
rect 26878 6876 26884 6928
rect 26936 6876 26942 6928
rect 22480 6820 24256 6848
rect 22373 6811 22431 6817
rect 19352 6752 19564 6780
rect 19426 6712 19432 6724
rect 17920 6684 19012 6712
rect 19260 6684 19432 6712
rect 17920 6672 17926 6684
rect 19260 6644 19288 6684
rect 19426 6672 19432 6684
rect 19484 6672 19490 6724
rect 19536 6712 19564 6752
rect 19610 6740 19616 6792
rect 19668 6740 19674 6792
rect 21358 6740 21364 6792
rect 21416 6780 21422 6792
rect 22189 6783 22247 6789
rect 22189 6780 22201 6783
rect 21416 6752 22201 6780
rect 21416 6740 21422 6752
rect 22189 6749 22201 6752
rect 22235 6780 22247 6783
rect 22388 6780 22508 6782
rect 22738 6780 22744 6792
rect 22235 6754 22744 6780
rect 22235 6752 22416 6754
rect 22480 6752 22744 6754
rect 22235 6749 22247 6752
rect 22189 6743 22247 6749
rect 22738 6740 22744 6752
rect 22796 6740 22802 6792
rect 22922 6740 22928 6792
rect 22980 6780 22986 6792
rect 23293 6783 23351 6789
rect 23293 6780 23305 6783
rect 22980 6752 23305 6780
rect 22980 6740 22986 6752
rect 23293 6749 23305 6752
rect 23339 6749 23351 6783
rect 23293 6743 23351 6749
rect 23474 6740 23480 6792
rect 23532 6740 23538 6792
rect 23566 6740 23572 6792
rect 23624 6780 23630 6792
rect 24228 6789 24256 6820
rect 24964 6820 25820 6848
rect 23753 6783 23811 6789
rect 23753 6780 23765 6783
rect 23624 6752 23765 6780
rect 23624 6740 23630 6752
rect 23753 6749 23765 6752
rect 23799 6749 23811 6783
rect 23753 6743 23811 6749
rect 24213 6783 24271 6789
rect 24213 6749 24225 6783
rect 24259 6749 24271 6783
rect 24213 6743 24271 6749
rect 24397 6783 24455 6789
rect 24397 6749 24409 6783
rect 24443 6749 24455 6783
rect 24397 6743 24455 6749
rect 20254 6712 20260 6724
rect 19536 6684 20260 6712
rect 20254 6672 20260 6684
rect 20312 6672 20318 6724
rect 22278 6672 22284 6724
rect 22336 6712 22342 6724
rect 22336 6684 24056 6712
rect 22336 6672 22342 6684
rect 17788 6616 19288 6644
rect 20349 6647 20407 6653
rect 20349 6613 20361 6647
rect 20395 6644 20407 6647
rect 21726 6644 21732 6656
rect 20395 6616 21732 6644
rect 20395 6613 20407 6616
rect 20349 6607 20407 6613
rect 21726 6604 21732 6616
rect 21784 6604 21790 6656
rect 22002 6604 22008 6656
rect 22060 6644 22066 6656
rect 22557 6647 22615 6653
rect 22557 6644 22569 6647
rect 22060 6616 22569 6644
rect 22060 6604 22066 6616
rect 22557 6613 22569 6616
rect 22603 6613 22615 6647
rect 22557 6607 22615 6613
rect 22646 6604 22652 6656
rect 22704 6604 22710 6656
rect 22922 6604 22928 6656
rect 22980 6644 22986 6656
rect 23017 6647 23075 6653
rect 23017 6644 23029 6647
rect 22980 6616 23029 6644
rect 22980 6604 22986 6616
rect 23017 6613 23029 6616
rect 23063 6613 23075 6647
rect 23017 6607 23075 6613
rect 23106 6604 23112 6656
rect 23164 6604 23170 6656
rect 23934 6604 23940 6656
rect 23992 6604 23998 6656
rect 24028 6644 24056 6684
rect 24118 6672 24124 6724
rect 24176 6712 24182 6724
rect 24412 6712 24440 6743
rect 24670 6740 24676 6792
rect 24728 6740 24734 6792
rect 24762 6740 24768 6792
rect 24820 6780 24826 6792
rect 24964 6780 24992 6820
rect 27522 6808 27528 6860
rect 27580 6848 27586 6860
rect 27709 6851 27767 6857
rect 27709 6848 27721 6851
rect 27580 6820 27721 6848
rect 27580 6808 27586 6820
rect 27709 6817 27721 6820
rect 27755 6817 27767 6851
rect 27709 6811 27767 6817
rect 24820 6752 24992 6780
rect 24820 6740 24826 6752
rect 25130 6740 25136 6792
rect 25188 6780 25194 6792
rect 25685 6783 25743 6789
rect 25685 6780 25697 6783
rect 25188 6752 25697 6780
rect 25188 6740 25194 6752
rect 25685 6749 25697 6752
rect 25731 6749 25743 6783
rect 25685 6743 25743 6749
rect 26234 6740 26240 6792
rect 26292 6780 26298 6792
rect 26513 6783 26571 6789
rect 26513 6780 26525 6783
rect 26292 6752 26525 6780
rect 26292 6740 26298 6752
rect 26513 6749 26525 6752
rect 26559 6749 26571 6783
rect 26513 6743 26571 6749
rect 26789 6783 26847 6789
rect 26789 6749 26801 6783
rect 26835 6749 26847 6783
rect 26789 6743 26847 6749
rect 24176 6684 25912 6712
rect 24176 6672 24182 6684
rect 24762 6644 24768 6656
rect 24028 6616 24768 6644
rect 24762 6604 24768 6616
rect 24820 6604 24826 6656
rect 24854 6604 24860 6656
rect 24912 6644 24918 6656
rect 25409 6647 25467 6653
rect 25409 6644 25421 6647
rect 24912 6616 25421 6644
rect 24912 6604 24918 6616
rect 25409 6613 25421 6616
rect 25455 6613 25467 6647
rect 25409 6607 25467 6613
rect 25498 6604 25504 6656
rect 25556 6604 25562 6656
rect 25884 6644 25912 6684
rect 25958 6672 25964 6724
rect 26016 6712 26022 6724
rect 26694 6712 26700 6724
rect 26016 6684 26700 6712
rect 26016 6672 26022 6684
rect 26694 6672 26700 6684
rect 26752 6672 26758 6724
rect 26804 6712 26832 6743
rect 27062 6740 27068 6792
rect 27120 6740 27126 6792
rect 27338 6740 27344 6792
rect 27396 6740 27402 6792
rect 27614 6740 27620 6792
rect 27672 6740 27678 6792
rect 27976 6783 28034 6789
rect 27976 6749 27988 6783
rect 28022 6780 28034 6783
rect 28258 6780 28264 6792
rect 28022 6752 28264 6780
rect 28022 6749 28034 6752
rect 27976 6743 28034 6749
rect 28258 6740 28264 6752
rect 28316 6740 28322 6792
rect 29012 6780 29040 6956
rect 29089 6953 29101 6987
rect 29135 6984 29147 6987
rect 30098 6984 30104 6996
rect 29135 6956 30104 6984
rect 29135 6953 29147 6956
rect 29089 6947 29147 6953
rect 30098 6944 30104 6956
rect 30156 6944 30162 6996
rect 31110 6944 31116 6996
rect 31168 6984 31174 6996
rect 32306 6984 32312 6996
rect 31168 6956 32312 6984
rect 31168 6944 31174 6956
rect 32306 6944 32312 6956
rect 32364 6944 32370 6996
rect 34514 6944 34520 6996
rect 34572 6944 34578 6996
rect 35802 6944 35808 6996
rect 35860 6984 35866 6996
rect 39206 6984 39212 6996
rect 35860 6956 39212 6984
rect 35860 6944 35866 6956
rect 39206 6944 39212 6956
rect 39264 6944 39270 6996
rect 29365 6919 29423 6925
rect 29365 6885 29377 6919
rect 29411 6916 29423 6919
rect 29411 6888 30052 6916
rect 29411 6885 29423 6888
rect 29365 6879 29423 6885
rect 29086 6808 29092 6860
rect 29144 6848 29150 6860
rect 29917 6851 29975 6857
rect 29917 6848 29929 6851
rect 29144 6820 29929 6848
rect 29144 6808 29150 6820
rect 29917 6817 29929 6820
rect 29963 6817 29975 6851
rect 30024 6848 30052 6888
rect 31018 6876 31024 6928
rect 31076 6876 31082 6928
rect 33689 6919 33747 6925
rect 33689 6885 33701 6919
rect 33735 6885 33747 6919
rect 33689 6879 33747 6885
rect 30466 6848 30472 6860
rect 30024 6820 30472 6848
rect 29917 6811 29975 6817
rect 30466 6808 30472 6820
rect 30524 6808 30530 6860
rect 30745 6851 30803 6857
rect 30745 6817 30757 6851
rect 30791 6848 30803 6851
rect 31202 6848 31208 6860
rect 30791 6820 31208 6848
rect 30791 6817 30803 6820
rect 30745 6811 30803 6817
rect 31202 6808 31208 6820
rect 31260 6808 31266 6860
rect 31386 6808 31392 6860
rect 31444 6808 31450 6860
rect 31662 6808 31668 6860
rect 31720 6848 31726 6860
rect 33704 6848 33732 6879
rect 35710 6876 35716 6928
rect 35768 6916 35774 6928
rect 37274 6916 37280 6928
rect 35768 6888 37280 6916
rect 35768 6876 35774 6888
rect 37274 6876 37280 6888
rect 37332 6876 37338 6928
rect 38197 6919 38255 6925
rect 38197 6885 38209 6919
rect 38243 6885 38255 6919
rect 38197 6879 38255 6885
rect 33873 6851 33931 6857
rect 33873 6848 33885 6851
rect 31720 6820 31984 6848
rect 33704 6820 33885 6848
rect 31720 6808 31726 6820
rect 29181 6783 29239 6789
rect 29181 6780 29193 6783
rect 29012 6752 29193 6780
rect 29181 6749 29193 6752
rect 29227 6749 29239 6783
rect 29181 6743 29239 6749
rect 29454 6740 29460 6792
rect 29512 6780 29518 6792
rect 29549 6783 29607 6789
rect 29549 6780 29561 6783
rect 29512 6752 29561 6780
rect 29512 6740 29518 6752
rect 29549 6749 29561 6752
rect 29595 6749 29607 6783
rect 29549 6743 29607 6749
rect 29822 6740 29828 6792
rect 29880 6740 29886 6792
rect 30009 6783 30067 6789
rect 30009 6749 30021 6783
rect 30055 6780 30067 6783
rect 30190 6780 30196 6792
rect 30055 6752 30196 6780
rect 30055 6749 30067 6752
rect 30009 6743 30067 6749
rect 30190 6740 30196 6752
rect 30248 6740 30254 6792
rect 30285 6783 30343 6789
rect 30285 6749 30297 6783
rect 30331 6749 30343 6783
rect 30285 6743 30343 6749
rect 27706 6712 27712 6724
rect 26804 6684 27712 6712
rect 26804 6644 26832 6684
rect 27706 6672 27712 6684
rect 27764 6672 27770 6724
rect 28626 6672 28632 6724
rect 28684 6712 28690 6724
rect 30300 6712 30328 6743
rect 30558 6740 30564 6792
rect 30616 6780 30622 6792
rect 30653 6783 30711 6789
rect 30653 6780 30665 6783
rect 30616 6752 30665 6780
rect 30616 6740 30622 6752
rect 30653 6749 30665 6752
rect 30699 6749 30711 6783
rect 30653 6743 30711 6749
rect 31478 6740 31484 6792
rect 31536 6740 31542 6792
rect 31956 6789 31984 6820
rect 33873 6817 33885 6820
rect 33919 6817 33931 6851
rect 33873 6811 33931 6817
rect 35894 6808 35900 6860
rect 35952 6848 35958 6860
rect 38212 6848 38240 6879
rect 35952 6820 38240 6848
rect 35952 6808 35958 6820
rect 31941 6783 31999 6789
rect 31941 6749 31953 6783
rect 31987 6749 31999 6783
rect 31941 6743 31999 6749
rect 32030 6740 32036 6792
rect 32088 6780 32094 6792
rect 32217 6783 32275 6789
rect 32217 6780 32229 6783
rect 32088 6752 32229 6780
rect 32088 6740 32094 6752
rect 32217 6749 32229 6752
rect 32263 6749 32275 6783
rect 32217 6743 32275 6749
rect 32398 6740 32404 6792
rect 32456 6780 32462 6792
rect 32493 6783 32551 6789
rect 32493 6780 32505 6783
rect 32456 6752 32505 6780
rect 32456 6740 32462 6752
rect 32493 6749 32505 6752
rect 32539 6749 32551 6783
rect 32493 6743 32551 6749
rect 32677 6783 32735 6789
rect 32677 6749 32689 6783
rect 32723 6749 32735 6783
rect 32677 6743 32735 6749
rect 28684 6684 30328 6712
rect 28684 6672 28690 6684
rect 30834 6672 30840 6724
rect 30892 6712 30898 6724
rect 31662 6712 31668 6724
rect 30892 6684 31668 6712
rect 30892 6672 30898 6684
rect 31662 6672 31668 6684
rect 31720 6672 31726 6724
rect 32692 6712 32720 6743
rect 32950 6740 32956 6792
rect 33008 6740 33014 6792
rect 35345 6783 35403 6789
rect 35345 6749 35357 6783
rect 35391 6780 35403 6783
rect 35434 6780 35440 6792
rect 35391 6752 35440 6780
rect 35391 6749 35403 6752
rect 35345 6743 35403 6749
rect 35434 6740 35440 6752
rect 35492 6740 35498 6792
rect 35989 6783 36047 6789
rect 35989 6749 36001 6783
rect 36035 6780 36047 6783
rect 36078 6780 36084 6792
rect 36035 6752 36084 6780
rect 36035 6749 36047 6752
rect 35989 6743 36047 6749
rect 36078 6740 36084 6752
rect 36136 6740 36142 6792
rect 36170 6740 36176 6792
rect 36228 6780 36234 6792
rect 37921 6783 37979 6789
rect 37921 6780 37933 6783
rect 36228 6752 37933 6780
rect 36228 6740 36234 6752
rect 37921 6749 37933 6752
rect 37967 6749 37979 6783
rect 37921 6743 37979 6749
rect 38105 6783 38163 6789
rect 38105 6749 38117 6783
rect 38151 6780 38163 6783
rect 38381 6783 38439 6789
rect 38381 6780 38393 6783
rect 38151 6752 38393 6780
rect 38151 6749 38163 6752
rect 38105 6743 38163 6749
rect 38381 6749 38393 6752
rect 38427 6749 38439 6783
rect 38381 6743 38439 6749
rect 38470 6740 38476 6792
rect 38528 6740 38534 6792
rect 38838 6740 38844 6792
rect 38896 6740 38902 6792
rect 39209 6783 39267 6789
rect 39209 6749 39221 6783
rect 39255 6749 39267 6783
rect 39209 6743 39267 6749
rect 32766 6712 32772 6724
rect 32692 6684 32772 6712
rect 32766 6672 32772 6684
rect 32824 6712 32830 6724
rect 34790 6712 34796 6724
rect 32824 6684 34796 6712
rect 32824 6672 32830 6684
rect 34790 6672 34796 6684
rect 34848 6672 34854 6724
rect 39224 6712 39252 6743
rect 39666 6712 39672 6724
rect 35544 6684 39252 6712
rect 39316 6684 39672 6712
rect 25884 6616 26832 6644
rect 26878 6604 26884 6656
rect 26936 6644 26942 6656
rect 27157 6647 27215 6653
rect 27157 6644 27169 6647
rect 26936 6616 27169 6644
rect 26936 6604 26942 6616
rect 27157 6613 27169 6616
rect 27203 6613 27215 6647
rect 27157 6607 27215 6613
rect 27338 6604 27344 6656
rect 27396 6644 27402 6656
rect 27433 6647 27491 6653
rect 27433 6644 27445 6647
rect 27396 6616 27445 6644
rect 27396 6604 27402 6616
rect 27433 6613 27445 6616
rect 27479 6613 27491 6647
rect 27433 6607 27491 6613
rect 28994 6604 29000 6656
rect 29052 6644 29058 6656
rect 29089 6647 29147 6653
rect 29089 6644 29101 6647
rect 29052 6616 29101 6644
rect 29052 6604 29058 6616
rect 29089 6613 29101 6616
rect 29135 6613 29147 6647
rect 29089 6607 29147 6613
rect 29638 6604 29644 6656
rect 29696 6644 29702 6656
rect 29733 6647 29791 6653
rect 29733 6644 29745 6647
rect 29696 6616 29745 6644
rect 29696 6604 29702 6616
rect 29733 6613 29745 6616
rect 29779 6613 29791 6647
rect 29733 6607 29791 6613
rect 29914 6604 29920 6656
rect 29972 6644 29978 6656
rect 30101 6647 30159 6653
rect 30101 6644 30113 6647
rect 29972 6616 30113 6644
rect 29972 6604 29978 6616
rect 30101 6613 30113 6616
rect 30147 6613 30159 6647
rect 30101 6607 30159 6613
rect 30650 6604 30656 6656
rect 30708 6644 30714 6656
rect 31113 6647 31171 6653
rect 31113 6644 31125 6647
rect 30708 6616 31125 6644
rect 30708 6604 30714 6616
rect 31113 6613 31125 6616
rect 31159 6613 31171 6647
rect 31113 6607 31171 6613
rect 31757 6647 31815 6653
rect 31757 6613 31769 6647
rect 31803 6644 31815 6647
rect 31846 6644 31852 6656
rect 31803 6616 31852 6644
rect 31803 6613 31815 6616
rect 31757 6607 31815 6613
rect 31846 6604 31852 6616
rect 31904 6604 31910 6656
rect 32030 6604 32036 6656
rect 32088 6604 32094 6656
rect 32306 6604 32312 6656
rect 32364 6604 32370 6656
rect 34054 6604 34060 6656
rect 34112 6604 34118 6656
rect 34146 6604 34152 6656
rect 34204 6604 34210 6656
rect 35544 6653 35572 6684
rect 35529 6647 35587 6653
rect 35529 6613 35541 6647
rect 35575 6613 35587 6647
rect 35529 6607 35587 6613
rect 35618 6604 35624 6656
rect 35676 6644 35682 6656
rect 35805 6647 35863 6653
rect 35805 6644 35817 6647
rect 35676 6616 35817 6644
rect 35676 6604 35682 6616
rect 35805 6613 35817 6616
rect 35851 6613 35863 6647
rect 35805 6607 35863 6613
rect 36722 6604 36728 6656
rect 36780 6644 36786 6656
rect 37737 6647 37795 6653
rect 37737 6644 37749 6647
rect 36780 6616 37749 6644
rect 36780 6604 36786 6616
rect 37737 6613 37749 6616
rect 37783 6613 37795 6647
rect 37737 6607 37795 6613
rect 38010 6604 38016 6656
rect 38068 6604 38074 6656
rect 38654 6604 38660 6656
rect 38712 6604 38718 6656
rect 39025 6647 39083 6653
rect 39025 6613 39037 6647
rect 39071 6644 39083 6647
rect 39316 6644 39344 6684
rect 39666 6672 39672 6684
rect 39724 6672 39730 6724
rect 39071 6616 39344 6644
rect 39393 6647 39451 6653
rect 39071 6613 39083 6616
rect 39025 6607 39083 6613
rect 39393 6613 39405 6647
rect 39439 6644 39451 6647
rect 39482 6644 39488 6656
rect 39439 6616 39488 6644
rect 39439 6613 39451 6616
rect 39393 6607 39451 6613
rect 39482 6604 39488 6616
rect 39540 6604 39546 6656
rect 1104 6554 39836 6576
rect 1104 6502 3010 6554
rect 3062 6502 3074 6554
rect 3126 6502 3138 6554
rect 3190 6502 3202 6554
rect 3254 6502 3266 6554
rect 3318 6502 9010 6554
rect 9062 6502 9074 6554
rect 9126 6502 9138 6554
rect 9190 6502 9202 6554
rect 9254 6502 9266 6554
rect 9318 6502 15010 6554
rect 15062 6502 15074 6554
rect 15126 6502 15138 6554
rect 15190 6502 15202 6554
rect 15254 6502 15266 6554
rect 15318 6502 21010 6554
rect 21062 6502 21074 6554
rect 21126 6502 21138 6554
rect 21190 6502 21202 6554
rect 21254 6502 21266 6554
rect 21318 6502 27010 6554
rect 27062 6502 27074 6554
rect 27126 6502 27138 6554
rect 27190 6502 27202 6554
rect 27254 6502 27266 6554
rect 27318 6502 33010 6554
rect 33062 6502 33074 6554
rect 33126 6502 33138 6554
rect 33190 6502 33202 6554
rect 33254 6502 33266 6554
rect 33318 6502 39010 6554
rect 39062 6502 39074 6554
rect 39126 6502 39138 6554
rect 39190 6502 39202 6554
rect 39254 6502 39266 6554
rect 39318 6502 39836 6554
rect 1104 6480 39836 6502
rect 1486 6400 1492 6452
rect 1544 6440 1550 6452
rect 1581 6443 1639 6449
rect 1581 6440 1593 6443
rect 1544 6412 1593 6440
rect 1544 6400 1550 6412
rect 1581 6409 1593 6412
rect 1627 6409 1639 6443
rect 1581 6403 1639 6409
rect 2317 6443 2375 6449
rect 2317 6409 2329 6443
rect 2363 6440 2375 6443
rect 2866 6440 2872 6452
rect 2363 6412 2872 6440
rect 2363 6409 2375 6412
rect 2317 6403 2375 6409
rect 2866 6400 2872 6412
rect 2924 6400 2930 6452
rect 3418 6400 3424 6452
rect 3476 6440 3482 6452
rect 5350 6440 5356 6452
rect 3476 6412 5356 6440
rect 3476 6400 3482 6412
rect 5350 6400 5356 6412
rect 5408 6400 5414 6452
rect 5997 6443 6055 6449
rect 5997 6409 6009 6443
rect 6043 6440 6055 6443
rect 6178 6440 6184 6452
rect 6043 6412 6184 6440
rect 6043 6409 6055 6412
rect 5997 6403 6055 6409
rect 6178 6400 6184 6412
rect 6236 6400 6242 6452
rect 6454 6400 6460 6452
rect 6512 6400 6518 6452
rect 6825 6443 6883 6449
rect 6825 6409 6837 6443
rect 6871 6440 6883 6443
rect 7006 6440 7012 6452
rect 6871 6412 7012 6440
rect 6871 6409 6883 6412
rect 6825 6403 6883 6409
rect 7006 6400 7012 6412
rect 7064 6400 7070 6452
rect 7098 6400 7104 6452
rect 7156 6440 7162 6452
rect 7193 6443 7251 6449
rect 7193 6440 7205 6443
rect 7156 6412 7205 6440
rect 7156 6400 7162 6412
rect 7193 6409 7205 6412
rect 7239 6409 7251 6443
rect 7193 6403 7251 6409
rect 7558 6400 7564 6452
rect 7616 6400 7622 6452
rect 7742 6400 7748 6452
rect 7800 6440 7806 6452
rect 7800 6412 8616 6440
rect 7800 6400 7806 6412
rect 1302 6332 1308 6384
rect 1360 6372 1366 6384
rect 1949 6375 2007 6381
rect 1949 6372 1961 6375
rect 1360 6344 1961 6372
rect 1360 6332 1366 6344
rect 1949 6341 1961 6344
rect 1995 6341 2007 6375
rect 1949 6335 2007 6341
rect 2406 6332 2412 6384
rect 2464 6372 2470 6384
rect 3697 6375 3755 6381
rect 3697 6372 3709 6375
rect 2464 6344 3709 6372
rect 2464 6332 2470 6344
rect 3697 6341 3709 6344
rect 3743 6372 3755 6375
rect 3970 6372 3976 6384
rect 3743 6344 3976 6372
rect 3743 6341 3755 6344
rect 3697 6335 3755 6341
rect 3970 6332 3976 6344
rect 4028 6332 4034 6384
rect 4338 6372 4344 6384
rect 4172 6344 4344 6372
rect 1765 6307 1823 6313
rect 1765 6273 1777 6307
rect 1811 6273 1823 6307
rect 1765 6267 1823 6273
rect 1780 6168 1808 6267
rect 1854 6264 1860 6316
rect 1912 6304 1918 6316
rect 2501 6307 2559 6313
rect 2501 6304 2513 6307
rect 1912 6276 2513 6304
rect 1912 6264 1918 6276
rect 2501 6273 2513 6276
rect 2547 6273 2559 6307
rect 2501 6267 2559 6273
rect 3145 6307 3203 6313
rect 3145 6273 3157 6307
rect 3191 6304 3203 6307
rect 4172 6304 4200 6344
rect 4338 6332 4344 6344
rect 4396 6332 4402 6384
rect 7466 6332 7472 6384
rect 7524 6372 7530 6384
rect 7524 6344 7880 6372
rect 7524 6332 7530 6344
rect 3191 6276 4200 6304
rect 4249 6307 4307 6313
rect 3191 6273 3203 6276
rect 3145 6267 3203 6273
rect 4249 6273 4261 6307
rect 4295 6304 4307 6307
rect 4430 6304 4436 6316
rect 4295 6276 4436 6304
rect 4295 6273 4307 6276
rect 4249 6267 4307 6273
rect 4430 6264 4436 6276
rect 4488 6264 4494 6316
rect 4614 6264 4620 6316
rect 4672 6264 4678 6316
rect 4985 6307 5043 6313
rect 4985 6273 4997 6307
rect 5031 6304 5043 6307
rect 5442 6304 5448 6316
rect 5031 6276 5448 6304
rect 5031 6273 5043 6276
rect 4985 6267 5043 6273
rect 5442 6264 5448 6276
rect 5500 6304 5506 6316
rect 5902 6304 5908 6316
rect 5500 6276 5908 6304
rect 5500 6264 5506 6276
rect 5902 6264 5908 6276
rect 5960 6264 5966 6316
rect 6181 6307 6239 6313
rect 6181 6273 6193 6307
rect 6227 6273 6239 6307
rect 6181 6267 6239 6273
rect 2130 6196 2136 6248
rect 2188 6196 2194 6248
rect 3237 6239 3295 6245
rect 3237 6205 3249 6239
rect 3283 6205 3295 6239
rect 3237 6199 3295 6205
rect 3142 6168 3148 6180
rect 1780 6140 3148 6168
rect 3142 6128 3148 6140
rect 3200 6128 3206 6180
rect 2777 6103 2835 6109
rect 2777 6069 2789 6103
rect 2823 6100 2835 6103
rect 2866 6100 2872 6112
rect 2823 6072 2872 6100
rect 2823 6069 2835 6072
rect 2777 6063 2835 6069
rect 2866 6060 2872 6072
rect 2924 6060 2930 6112
rect 3252 6100 3280 6199
rect 3326 6196 3332 6248
rect 3384 6196 3390 6248
rect 4709 6239 4767 6245
rect 4709 6205 4721 6239
rect 4755 6205 4767 6239
rect 6196 6236 6224 6267
rect 6638 6264 6644 6316
rect 6696 6264 6702 6316
rect 7009 6307 7067 6313
rect 7009 6273 7021 6307
rect 7055 6304 7067 6307
rect 7098 6304 7104 6316
rect 7055 6276 7104 6304
rect 7055 6273 7067 6276
rect 7009 6267 7067 6273
rect 7098 6264 7104 6276
rect 7156 6264 7162 6316
rect 7282 6264 7288 6316
rect 7340 6304 7346 6316
rect 7377 6307 7435 6313
rect 7377 6304 7389 6307
rect 7340 6276 7389 6304
rect 7340 6264 7346 6276
rect 7377 6273 7389 6276
rect 7423 6273 7435 6307
rect 7377 6267 7435 6273
rect 7558 6264 7564 6316
rect 7616 6304 7622 6316
rect 7852 6313 7880 6344
rect 8110 6332 8116 6384
rect 8168 6372 8174 6384
rect 8297 6375 8355 6381
rect 8297 6372 8309 6375
rect 8168 6344 8309 6372
rect 8168 6332 8174 6344
rect 8297 6341 8309 6344
rect 8343 6341 8355 6375
rect 8297 6335 8355 6341
rect 8588 6372 8616 6412
rect 8754 6400 8760 6452
rect 8812 6440 8818 6452
rect 9401 6443 9459 6449
rect 8812 6412 9352 6440
rect 8812 6400 8818 6412
rect 9030 6372 9036 6384
rect 8588 6344 9036 6372
rect 8588 6313 8616 6344
rect 9030 6332 9036 6344
rect 9088 6332 9094 6384
rect 7745 6307 7803 6313
rect 7745 6304 7757 6307
rect 7616 6276 7757 6304
rect 7616 6264 7622 6276
rect 7745 6273 7757 6276
rect 7791 6273 7803 6307
rect 7745 6267 7803 6273
rect 7837 6307 7895 6313
rect 7837 6273 7849 6307
rect 7883 6273 7895 6307
rect 7837 6267 7895 6273
rect 8021 6307 8079 6313
rect 8021 6273 8033 6307
rect 8067 6273 8079 6307
rect 8021 6267 8079 6273
rect 8205 6307 8263 6313
rect 8205 6273 8217 6307
rect 8251 6273 8263 6307
rect 8205 6267 8263 6273
rect 8573 6307 8631 6313
rect 8573 6273 8585 6307
rect 8619 6273 8631 6307
rect 8573 6267 8631 6273
rect 7650 6236 7656 6248
rect 6196 6208 7656 6236
rect 4709 6199 4767 6205
rect 3881 6171 3939 6177
rect 3881 6137 3893 6171
rect 3927 6168 3939 6171
rect 3970 6168 3976 6180
rect 3927 6140 3976 6168
rect 3927 6137 3939 6140
rect 3881 6131 3939 6137
rect 3970 6128 3976 6140
rect 4028 6128 4034 6180
rect 4433 6171 4491 6177
rect 4433 6137 4445 6171
rect 4479 6168 4491 6171
rect 4522 6168 4528 6180
rect 4479 6140 4528 6168
rect 4479 6137 4491 6140
rect 4433 6131 4491 6137
rect 4522 6128 4528 6140
rect 4580 6128 4586 6180
rect 4614 6128 4620 6180
rect 4672 6168 4678 6180
rect 4724 6168 4752 6199
rect 7650 6196 7656 6208
rect 7708 6196 7714 6248
rect 8036 6236 8064 6267
rect 8110 6236 8116 6248
rect 8036 6208 8116 6236
rect 8110 6196 8116 6208
rect 8168 6196 8174 6248
rect 8220 6236 8248 6267
rect 8662 6264 8668 6316
rect 8720 6264 8726 6316
rect 8754 6264 8760 6316
rect 8812 6264 8818 6316
rect 8941 6307 8999 6313
rect 8941 6273 8953 6307
rect 8987 6304 8999 6307
rect 9122 6304 9128 6316
rect 8987 6276 9128 6304
rect 8987 6273 8999 6276
rect 8941 6267 8999 6273
rect 8680 6236 8708 6264
rect 8220 6208 8708 6236
rect 4672 6140 4752 6168
rect 5368 6140 5856 6168
rect 4672 6128 4678 6140
rect 3602 6100 3608 6112
rect 3252 6072 3608 6100
rect 3602 6060 3608 6072
rect 3660 6060 3666 6112
rect 3694 6060 3700 6112
rect 3752 6100 3758 6112
rect 4065 6103 4123 6109
rect 4065 6100 4077 6103
rect 3752 6072 4077 6100
rect 3752 6060 3758 6072
rect 4065 6069 4077 6072
rect 4111 6069 4123 6103
rect 4065 6063 4123 6069
rect 4706 6060 4712 6112
rect 4764 6100 4770 6112
rect 5368 6100 5396 6140
rect 4764 6072 5396 6100
rect 4764 6060 4770 6072
rect 5534 6060 5540 6112
rect 5592 6100 5598 6112
rect 5721 6103 5779 6109
rect 5721 6100 5733 6103
rect 5592 6072 5733 6100
rect 5592 6060 5598 6072
rect 5721 6069 5733 6072
rect 5767 6069 5779 6103
rect 5828 6100 5856 6140
rect 6454 6128 6460 6180
rect 6512 6168 6518 6180
rect 7742 6168 7748 6180
rect 6512 6140 7748 6168
rect 6512 6128 6518 6140
rect 7742 6128 7748 6140
rect 7800 6128 7806 6180
rect 8018 6128 8024 6180
rect 8076 6168 8082 6180
rect 8956 6168 8984 6267
rect 9122 6264 9128 6276
rect 9180 6264 9186 6316
rect 9217 6307 9275 6313
rect 9217 6273 9229 6307
rect 9263 6273 9275 6307
rect 9324 6304 9352 6412
rect 9401 6409 9413 6443
rect 9447 6440 9459 6443
rect 10502 6440 10508 6452
rect 9447 6412 10508 6440
rect 9447 6409 9459 6412
rect 9401 6403 9459 6409
rect 10502 6400 10508 6412
rect 10560 6440 10566 6452
rect 10686 6440 10692 6452
rect 10560 6412 10692 6440
rect 10560 6400 10566 6412
rect 10686 6400 10692 6412
rect 10744 6400 10750 6452
rect 10781 6443 10839 6449
rect 10781 6409 10793 6443
rect 10827 6440 10839 6443
rect 10870 6440 10876 6452
rect 10827 6412 10876 6440
rect 10827 6409 10839 6412
rect 10781 6403 10839 6409
rect 10870 6400 10876 6412
rect 10928 6400 10934 6452
rect 11072 6412 12112 6440
rect 9490 6332 9496 6384
rect 9548 6332 9554 6384
rect 10321 6375 10379 6381
rect 10321 6341 10333 6375
rect 10367 6372 10379 6375
rect 10410 6372 10416 6384
rect 10367 6344 10416 6372
rect 10367 6341 10379 6344
rect 10321 6335 10379 6341
rect 10410 6332 10416 6344
rect 10468 6332 10474 6384
rect 9582 6304 9588 6316
rect 9324 6276 9588 6304
rect 9217 6267 9275 6273
rect 9033 6239 9091 6245
rect 9033 6205 9045 6239
rect 9079 6205 9091 6239
rect 9232 6236 9260 6267
rect 9582 6264 9588 6276
rect 9640 6264 9646 6316
rect 10134 6264 10140 6316
rect 10192 6304 10198 6316
rect 11072 6313 11100 6412
rect 11333 6375 11391 6381
rect 11333 6341 11345 6375
rect 11379 6372 11391 6375
rect 12084 6372 12112 6412
rect 12158 6400 12164 6452
rect 12216 6440 12222 6452
rect 18230 6440 18236 6452
rect 12216 6412 18236 6440
rect 12216 6400 12222 6412
rect 18230 6400 18236 6412
rect 18288 6400 18294 6452
rect 18322 6400 18328 6452
rect 18380 6440 18386 6452
rect 25958 6440 25964 6452
rect 18380 6412 25964 6440
rect 18380 6400 18386 6412
rect 25958 6400 25964 6412
rect 26016 6400 26022 6452
rect 26418 6400 26424 6452
rect 26476 6440 26482 6452
rect 26513 6443 26571 6449
rect 26513 6440 26525 6443
rect 26476 6412 26525 6440
rect 26476 6400 26482 6412
rect 26513 6409 26525 6412
rect 26559 6409 26571 6443
rect 26513 6403 26571 6409
rect 26786 6400 26792 6452
rect 26844 6400 26850 6452
rect 26970 6400 26976 6452
rect 27028 6440 27034 6452
rect 27433 6443 27491 6449
rect 27433 6440 27445 6443
rect 27028 6412 27445 6440
rect 27028 6400 27034 6412
rect 27433 6409 27445 6412
rect 27479 6409 27491 6443
rect 27433 6403 27491 6409
rect 27522 6400 27528 6452
rect 27580 6440 27586 6452
rect 27580 6412 28994 6440
rect 27580 6400 27586 6412
rect 12710 6372 12716 6384
rect 11379 6344 12020 6372
rect 12084 6344 12716 6372
rect 11379 6341 11391 6344
rect 11333 6335 11391 6341
rect 10505 6307 10563 6313
rect 10505 6304 10517 6307
rect 10192 6276 10517 6304
rect 10192 6264 10198 6276
rect 10505 6273 10517 6276
rect 10551 6273 10563 6307
rect 10505 6267 10563 6273
rect 10597 6307 10655 6313
rect 10597 6273 10609 6307
rect 10643 6273 10655 6307
rect 10597 6267 10655 6273
rect 11057 6307 11115 6313
rect 11057 6273 11069 6307
rect 11103 6273 11115 6307
rect 11057 6267 11115 6273
rect 11149 6307 11207 6313
rect 11149 6273 11161 6307
rect 11195 6304 11207 6307
rect 11238 6304 11244 6316
rect 11195 6276 11244 6304
rect 11195 6273 11207 6276
rect 11149 6267 11207 6273
rect 9398 6236 9404 6248
rect 9232 6208 9404 6236
rect 9033 6199 9091 6205
rect 8076 6140 8984 6168
rect 9048 6168 9076 6199
rect 9398 6196 9404 6208
rect 9456 6196 9462 6248
rect 10612 6236 10640 6267
rect 11238 6264 11244 6276
rect 11296 6264 11302 6316
rect 11882 6313 11888 6316
rect 11876 6304 11888 6313
rect 11843 6276 11888 6304
rect 11876 6267 11888 6276
rect 11882 6264 11888 6267
rect 11940 6264 11946 6316
rect 11992 6304 12020 6344
rect 12710 6332 12716 6344
rect 12768 6372 12774 6384
rect 12768 6344 13032 6372
rect 12768 6332 12774 6344
rect 13004 6304 13032 6344
rect 13538 6332 13544 6384
rect 13596 6372 13602 6384
rect 13814 6372 13820 6384
rect 13596 6344 13820 6372
rect 13596 6332 13602 6344
rect 13814 6332 13820 6344
rect 13872 6332 13878 6384
rect 13906 6332 13912 6384
rect 13964 6372 13970 6384
rect 15470 6372 15476 6384
rect 13964 6344 15476 6372
rect 13964 6332 13970 6344
rect 15470 6332 15476 6344
rect 15528 6372 15534 6384
rect 15528 6344 16344 6372
rect 15528 6332 15534 6344
rect 13633 6307 13691 6313
rect 13633 6304 13645 6307
rect 11992 6276 12940 6304
rect 13004 6276 13645 6304
rect 11422 6236 11428 6248
rect 10612 6208 11428 6236
rect 11422 6196 11428 6208
rect 11480 6196 11486 6248
rect 11609 6239 11667 6245
rect 11609 6205 11621 6239
rect 11655 6205 11667 6239
rect 12912 6236 12940 6276
rect 13633 6273 13645 6276
rect 13679 6273 13691 6307
rect 13633 6267 13691 6273
rect 14458 6264 14464 6316
rect 14516 6304 14522 6316
rect 15102 6304 15108 6316
rect 14516 6276 15108 6304
rect 14516 6264 14522 6276
rect 15102 6264 15108 6276
rect 15160 6264 15166 6316
rect 15562 6264 15568 6316
rect 15620 6304 15626 6316
rect 16316 6313 16344 6344
rect 16390 6332 16396 6384
rect 16448 6332 16454 6384
rect 17218 6332 17224 6384
rect 17276 6372 17282 6384
rect 17402 6372 17408 6384
rect 17276 6344 17408 6372
rect 17276 6332 17282 6344
rect 17402 6332 17408 6344
rect 17460 6332 17466 6384
rect 17862 6332 17868 6384
rect 17920 6372 17926 6384
rect 19521 6375 19579 6381
rect 19521 6372 19533 6375
rect 17920 6344 19533 6372
rect 17920 6332 17926 6344
rect 19521 6341 19533 6344
rect 19567 6341 19579 6375
rect 19521 6335 19579 6341
rect 21269 6375 21327 6381
rect 21269 6341 21281 6375
rect 21315 6372 21327 6375
rect 21358 6372 21364 6384
rect 21315 6344 21364 6372
rect 21315 6341 21327 6344
rect 21269 6335 21327 6341
rect 21358 6332 21364 6344
rect 21416 6332 21422 6384
rect 22186 6332 22192 6384
rect 22244 6332 22250 6384
rect 22419 6341 22477 6347
rect 22419 6338 22431 6341
rect 15942 6307 16000 6313
rect 15942 6304 15954 6307
rect 15620 6276 15954 6304
rect 15620 6264 15626 6276
rect 15942 6273 15954 6276
rect 15988 6273 16000 6307
rect 15942 6267 16000 6273
rect 16301 6307 16359 6313
rect 16301 6273 16313 6307
rect 16347 6273 16359 6307
rect 16301 6267 16359 6273
rect 16479 6307 16537 6313
rect 16479 6273 16491 6307
rect 16525 6294 16537 6307
rect 16574 6294 16580 6316
rect 16525 6273 16580 6294
rect 16479 6267 16580 6273
rect 14182 6236 14188 6248
rect 12912 6208 14188 6236
rect 11609 6199 11667 6205
rect 10686 6168 10692 6180
rect 9048 6140 10692 6168
rect 8076 6128 8082 6140
rect 10686 6128 10692 6140
rect 10744 6128 10750 6180
rect 10226 6100 10232 6112
rect 5828 6072 10232 6100
rect 5721 6063 5779 6069
rect 10226 6060 10232 6072
rect 10284 6060 10290 6112
rect 10318 6060 10324 6112
rect 10376 6060 10382 6112
rect 10870 6060 10876 6112
rect 10928 6060 10934 6112
rect 11330 6060 11336 6112
rect 11388 6060 11394 6112
rect 11624 6100 11652 6199
rect 14182 6196 14188 6208
rect 14240 6236 14246 6248
rect 14553 6239 14611 6245
rect 14553 6236 14565 6239
rect 14240 6208 14565 6236
rect 14240 6196 14246 6208
rect 14553 6205 14565 6208
rect 14599 6205 14611 6239
rect 14553 6199 14611 6205
rect 16209 6239 16267 6245
rect 16209 6205 16221 6239
rect 16255 6205 16267 6239
rect 16209 6199 16267 6205
rect 13814 6128 13820 6180
rect 13872 6168 13878 6180
rect 14918 6168 14924 6180
rect 13872 6140 14924 6168
rect 13872 6128 13878 6140
rect 14918 6128 14924 6140
rect 14976 6128 14982 6180
rect 11974 6100 11980 6112
rect 11624 6072 11980 6100
rect 11974 6060 11980 6072
rect 12032 6060 12038 6112
rect 12710 6060 12716 6112
rect 12768 6100 12774 6112
rect 12989 6103 13047 6109
rect 12989 6100 13001 6103
rect 12768 6072 13001 6100
rect 12768 6060 12774 6072
rect 12989 6069 13001 6072
rect 13035 6069 13047 6103
rect 12989 6063 13047 6069
rect 13078 6060 13084 6112
rect 13136 6060 13142 6112
rect 13538 6060 13544 6112
rect 13596 6100 13602 6112
rect 14001 6103 14059 6109
rect 14001 6100 14013 6103
rect 13596 6072 14013 6100
rect 13596 6060 13602 6072
rect 14001 6069 14013 6072
rect 14047 6069 14059 6103
rect 14001 6063 14059 6069
rect 14550 6060 14556 6112
rect 14608 6100 14614 6112
rect 14829 6103 14887 6109
rect 14829 6100 14841 6103
rect 14608 6072 14841 6100
rect 14608 6060 14614 6072
rect 14829 6069 14841 6072
rect 14875 6069 14887 6103
rect 16224 6100 16252 6199
rect 16316 6168 16344 6267
rect 16500 6266 16580 6267
rect 16574 6264 16580 6266
rect 16632 6264 16638 6316
rect 16850 6264 16856 6316
rect 16908 6264 16914 6316
rect 16942 6264 16948 6316
rect 17000 6304 17006 6316
rect 17129 6308 17187 6313
rect 17052 6307 17187 6308
rect 17052 6304 17141 6307
rect 17000 6280 17141 6304
rect 17000 6276 17080 6280
rect 17000 6264 17006 6276
rect 17129 6273 17141 6280
rect 17175 6273 17187 6307
rect 17129 6267 17187 6273
rect 17681 6307 17739 6313
rect 17681 6273 17693 6307
rect 17727 6304 17739 6307
rect 17727 6276 18184 6304
rect 17727 6273 17739 6276
rect 17681 6267 17739 6273
rect 18156 6248 18184 6276
rect 18598 6264 18604 6316
rect 18656 6264 18662 6316
rect 18785 6307 18843 6313
rect 18785 6273 18797 6307
rect 18831 6273 18843 6307
rect 18785 6267 18843 6273
rect 19061 6307 19119 6313
rect 19061 6273 19073 6307
rect 19107 6304 19119 6307
rect 19242 6304 19248 6316
rect 19107 6276 19248 6304
rect 19107 6273 19119 6276
rect 19061 6267 19119 6273
rect 16390 6196 16396 6248
rect 16448 6236 16454 6248
rect 16669 6239 16727 6245
rect 16669 6236 16681 6239
rect 16448 6208 16681 6236
rect 16448 6196 16454 6208
rect 16669 6205 16681 6208
rect 16715 6205 16727 6239
rect 16669 6199 16727 6205
rect 17034 6196 17040 6248
rect 17092 6196 17098 6248
rect 17402 6196 17408 6248
rect 17460 6196 17466 6248
rect 18138 6196 18144 6248
rect 18196 6196 18202 6248
rect 18414 6196 18420 6248
rect 18472 6236 18478 6248
rect 18800 6236 18828 6267
rect 19242 6264 19248 6276
rect 19300 6264 19306 6316
rect 19429 6307 19487 6313
rect 19429 6273 19441 6307
rect 19475 6304 19487 6307
rect 20622 6304 20628 6316
rect 19475 6276 20628 6304
rect 19475 6273 19487 6276
rect 19429 6267 19487 6273
rect 20622 6264 20628 6276
rect 20680 6264 20686 6316
rect 21542 6264 21548 6316
rect 21600 6264 21606 6316
rect 22005 6307 22063 6313
rect 22005 6273 22017 6307
rect 22051 6304 22063 6307
rect 22094 6304 22100 6316
rect 22051 6276 22100 6304
rect 22051 6273 22063 6276
rect 22005 6267 22063 6273
rect 22094 6264 22100 6276
rect 22152 6264 22158 6316
rect 22404 6307 22431 6338
rect 22465 6316 22477 6341
rect 22646 6332 22652 6384
rect 22704 6372 22710 6384
rect 25498 6372 25504 6384
rect 22704 6344 25504 6372
rect 22704 6332 22710 6344
rect 25498 6332 25504 6344
rect 25556 6332 25562 6384
rect 25774 6332 25780 6384
rect 25832 6372 25838 6384
rect 25832 6344 27016 6372
rect 25832 6332 25838 6344
rect 22465 6307 22468 6316
rect 22404 6276 22468 6307
rect 22462 6264 22468 6276
rect 22520 6264 22526 6316
rect 22741 6307 22799 6313
rect 22741 6273 22753 6307
rect 22787 6273 22799 6307
rect 22741 6267 22799 6273
rect 22925 6307 22983 6313
rect 22925 6273 22937 6307
rect 22971 6304 22983 6307
rect 23106 6304 23112 6316
rect 22971 6276 23112 6304
rect 22971 6273 22983 6276
rect 22925 6267 22983 6273
rect 21913 6239 21971 6245
rect 21913 6236 21925 6239
rect 18472 6208 18828 6236
rect 19076 6208 21925 6236
rect 18472 6196 18478 6208
rect 19076 6180 19104 6208
rect 21913 6205 21925 6208
rect 21959 6205 21971 6239
rect 22756 6236 22784 6267
rect 23106 6264 23112 6276
rect 23164 6264 23170 6316
rect 23474 6264 23480 6316
rect 23532 6304 23538 6316
rect 24121 6307 24179 6313
rect 24121 6304 24133 6307
rect 23532 6276 24133 6304
rect 23532 6264 23538 6276
rect 24121 6273 24133 6276
rect 24167 6304 24179 6307
rect 24670 6304 24676 6316
rect 24167 6276 24676 6304
rect 24167 6273 24179 6276
rect 24121 6267 24179 6273
rect 24670 6264 24676 6276
rect 24728 6264 24734 6316
rect 25222 6264 25228 6316
rect 25280 6264 25286 6316
rect 25682 6264 25688 6316
rect 25740 6264 25746 6316
rect 25866 6264 25872 6316
rect 25924 6304 25930 6316
rect 25961 6307 26019 6313
rect 25961 6304 25973 6307
rect 25924 6276 25973 6304
rect 25924 6264 25930 6276
rect 25961 6273 25973 6276
rect 26007 6273 26019 6307
rect 25961 6267 26019 6273
rect 26234 6264 26240 6316
rect 26292 6304 26298 6316
rect 26329 6307 26387 6313
rect 26329 6304 26341 6307
rect 26292 6276 26341 6304
rect 26292 6264 26298 6276
rect 26329 6273 26341 6276
rect 26375 6273 26387 6307
rect 26329 6267 26387 6273
rect 26602 6264 26608 6316
rect 26660 6264 26666 6316
rect 26988 6313 27016 6344
rect 27080 6344 28019 6372
rect 26973 6307 27031 6313
rect 26973 6273 26985 6307
rect 27019 6273 27031 6307
rect 26973 6267 27031 6273
rect 23382 6236 23388 6248
rect 22756 6208 23388 6236
rect 21913 6199 21971 6205
rect 23382 6196 23388 6208
rect 23440 6196 23446 6248
rect 23566 6196 23572 6248
rect 23624 6236 23630 6248
rect 23845 6239 23903 6245
rect 23845 6236 23857 6239
rect 23624 6208 23857 6236
rect 23624 6196 23630 6208
rect 23845 6205 23857 6208
rect 23891 6205 23903 6239
rect 26620 6236 26648 6264
rect 27080 6236 27108 6344
rect 27614 6264 27620 6316
rect 27672 6264 27678 6316
rect 27991 6313 28019 6344
rect 27985 6307 28043 6313
rect 27985 6273 27997 6307
rect 28031 6273 28043 6307
rect 27985 6267 28043 6273
rect 26620 6208 27108 6236
rect 23845 6199 23903 6205
rect 27522 6196 27528 6248
rect 27580 6236 27586 6248
rect 27709 6239 27767 6245
rect 27709 6236 27721 6239
rect 27580 6208 27721 6236
rect 27580 6196 27586 6208
rect 27709 6205 27721 6208
rect 27755 6205 27767 6239
rect 28644 6236 28672 6412
rect 28966 6372 28994 6412
rect 29730 6400 29736 6452
rect 29788 6440 29794 6452
rect 29825 6443 29883 6449
rect 29825 6440 29837 6443
rect 29788 6412 29837 6440
rect 29788 6400 29794 6412
rect 29825 6409 29837 6412
rect 29871 6409 29883 6443
rect 29825 6403 29883 6409
rect 31386 6400 31392 6452
rect 31444 6400 31450 6452
rect 31570 6400 31576 6452
rect 31628 6440 31634 6452
rect 31665 6443 31723 6449
rect 31665 6440 31677 6443
rect 31628 6412 31677 6440
rect 31628 6400 31634 6412
rect 31665 6409 31677 6412
rect 31711 6409 31723 6443
rect 31665 6403 31723 6409
rect 31938 6400 31944 6452
rect 31996 6440 32002 6452
rect 33781 6443 33839 6449
rect 33781 6440 33793 6443
rect 31996 6412 33793 6440
rect 31996 6400 32002 6412
rect 33781 6409 33793 6412
rect 33827 6409 33839 6443
rect 33781 6403 33839 6409
rect 33873 6443 33931 6449
rect 33873 6409 33885 6443
rect 33919 6440 33931 6443
rect 34054 6440 34060 6452
rect 33919 6412 34060 6440
rect 33919 6409 33931 6412
rect 33873 6403 33931 6409
rect 34054 6400 34060 6412
rect 34112 6400 34118 6452
rect 34882 6400 34888 6452
rect 34940 6440 34946 6452
rect 35526 6440 35532 6452
rect 34940 6412 35532 6440
rect 34940 6400 34946 6412
rect 35526 6400 35532 6412
rect 35584 6400 35590 6452
rect 36078 6400 36084 6452
rect 36136 6400 36142 6452
rect 36906 6400 36912 6452
rect 36964 6440 36970 6452
rect 38470 6440 38476 6452
rect 36964 6412 38476 6440
rect 36964 6400 36970 6412
rect 38470 6400 38476 6412
rect 38528 6400 38534 6452
rect 39390 6400 39396 6452
rect 39448 6400 39454 6452
rect 28966 6344 29592 6372
rect 28718 6264 28724 6316
rect 28776 6304 28782 6316
rect 29089 6307 29147 6313
rect 29089 6304 29101 6307
rect 28776 6276 29101 6304
rect 28776 6264 28782 6276
rect 29089 6273 29101 6276
rect 29135 6273 29147 6307
rect 29564 6304 29592 6344
rect 31110 6332 31116 6384
rect 31168 6372 31174 6384
rect 36449 6375 36507 6381
rect 36449 6372 36461 6375
rect 31168 6344 36461 6372
rect 31168 6332 31174 6344
rect 36449 6341 36461 6344
rect 36495 6341 36507 6375
rect 36449 6335 36507 6341
rect 36630 6332 36636 6384
rect 36688 6372 36694 6384
rect 38838 6372 38844 6384
rect 36688 6344 38844 6372
rect 36688 6332 36694 6344
rect 38838 6332 38844 6344
rect 38896 6332 38902 6384
rect 30098 6304 30104 6316
rect 29564 6276 30104 6304
rect 29089 6267 29147 6273
rect 30098 6264 30104 6276
rect 30156 6264 30162 6316
rect 30282 6264 30288 6316
rect 30340 6264 30346 6316
rect 30650 6264 30656 6316
rect 30708 6304 30714 6316
rect 30708 6276 30972 6304
rect 30708 6264 30714 6276
rect 28813 6239 28871 6245
rect 28813 6236 28825 6239
rect 28644 6208 28825 6236
rect 27709 6199 27767 6205
rect 28813 6205 28825 6208
rect 28859 6205 28871 6239
rect 28813 6199 28871 6205
rect 30006 6196 30012 6248
rect 30064 6236 30070 6248
rect 30377 6239 30435 6245
rect 30377 6236 30389 6239
rect 30064 6208 30389 6236
rect 30064 6196 30070 6208
rect 30377 6205 30389 6208
rect 30423 6205 30435 6239
rect 30944 6236 30972 6276
rect 31018 6264 31024 6316
rect 31076 6304 31082 6316
rect 31481 6307 31539 6313
rect 31481 6304 31493 6307
rect 31076 6276 31493 6304
rect 31076 6264 31082 6276
rect 31481 6273 31493 6276
rect 31527 6273 31539 6307
rect 31481 6267 31539 6273
rect 31754 6264 31760 6316
rect 31812 6304 31818 6316
rect 31941 6307 31999 6313
rect 31941 6304 31953 6307
rect 31812 6276 31953 6304
rect 31812 6264 31818 6276
rect 31941 6273 31953 6276
rect 31987 6273 31999 6307
rect 32585 6307 32643 6313
rect 32585 6304 32597 6307
rect 31941 6267 31999 6273
rect 32048 6276 32597 6304
rect 32048 6236 32076 6276
rect 32585 6273 32597 6276
rect 32631 6273 32643 6307
rect 32585 6267 32643 6273
rect 34514 6264 34520 6316
rect 34572 6304 34578 6316
rect 35253 6307 35311 6313
rect 35253 6304 35265 6307
rect 34572 6276 35265 6304
rect 34572 6264 34578 6276
rect 35253 6273 35265 6276
rect 35299 6304 35311 6307
rect 35342 6304 35348 6316
rect 35299 6276 35348 6304
rect 35299 6273 35311 6276
rect 35253 6267 35311 6273
rect 35342 6264 35348 6276
rect 35400 6264 35406 6316
rect 35618 6264 35624 6316
rect 35676 6304 35682 6316
rect 36170 6304 36176 6316
rect 35676 6276 36176 6304
rect 35676 6264 35682 6276
rect 36170 6264 36176 6276
rect 36228 6264 36234 6316
rect 37090 6264 37096 6316
rect 37148 6304 37154 6316
rect 38565 6307 38623 6313
rect 38565 6304 38577 6307
rect 37148 6276 38577 6304
rect 37148 6264 37154 6276
rect 38565 6273 38577 6276
rect 38611 6273 38623 6307
rect 38565 6267 38623 6273
rect 38657 6307 38715 6313
rect 38657 6273 38669 6307
rect 38703 6273 38715 6307
rect 38657 6267 38715 6273
rect 39117 6307 39175 6313
rect 39117 6273 39129 6307
rect 39163 6304 39175 6307
rect 39209 6307 39267 6313
rect 39209 6304 39221 6307
rect 39163 6276 39221 6304
rect 39163 6273 39175 6276
rect 39117 6267 39175 6273
rect 39209 6273 39221 6276
rect 39255 6273 39267 6307
rect 39209 6267 39267 6273
rect 30944 6208 32076 6236
rect 30377 6199 30435 6205
rect 32306 6196 32312 6248
rect 32364 6196 32370 6248
rect 33873 6239 33931 6245
rect 33873 6236 33885 6239
rect 33244 6208 33885 6236
rect 16942 6168 16948 6180
rect 16316 6140 16948 6168
rect 16942 6128 16948 6140
rect 17000 6128 17006 6180
rect 18064 6140 18920 6168
rect 16298 6100 16304 6112
rect 16224 6072 16304 6100
rect 14829 6063 14887 6069
rect 16298 6060 16304 6072
rect 16356 6060 16362 6112
rect 17313 6103 17371 6109
rect 17313 6069 17325 6103
rect 17359 6100 17371 6103
rect 17494 6100 17500 6112
rect 17359 6072 17500 6100
rect 17359 6069 17371 6072
rect 17313 6063 17371 6069
rect 17494 6060 17500 6072
rect 17552 6060 17558 6112
rect 17678 6060 17684 6112
rect 17736 6100 17742 6112
rect 18064 6100 18092 6140
rect 17736 6072 18092 6100
rect 17736 6060 17742 6072
rect 18414 6060 18420 6112
rect 18472 6060 18478 6112
rect 18506 6060 18512 6112
rect 18564 6100 18570 6112
rect 18892 6109 18920 6140
rect 19058 6128 19064 6180
rect 19116 6128 19122 6180
rect 22278 6168 22284 6180
rect 19168 6140 22284 6168
rect 18601 6103 18659 6109
rect 18601 6100 18613 6103
rect 18564 6072 18613 6100
rect 18564 6060 18570 6072
rect 18601 6069 18613 6072
rect 18647 6069 18659 6103
rect 18601 6063 18659 6069
rect 18877 6103 18935 6109
rect 18877 6069 18889 6103
rect 18923 6100 18935 6103
rect 19168 6100 19196 6140
rect 22278 6128 22284 6140
rect 22336 6128 22342 6180
rect 22554 6128 22560 6180
rect 22612 6128 22618 6180
rect 23474 6168 23480 6180
rect 22848 6140 23480 6168
rect 18923 6072 19196 6100
rect 18923 6069 18935 6072
rect 18877 6063 18935 6069
rect 19242 6060 19248 6112
rect 19300 6060 19306 6112
rect 19426 6060 19432 6112
rect 19484 6100 19490 6112
rect 20809 6103 20867 6109
rect 20809 6100 20821 6103
rect 19484 6072 20821 6100
rect 19484 6060 19490 6072
rect 20809 6069 20821 6072
rect 20855 6069 20867 6103
rect 20809 6063 20867 6069
rect 21361 6103 21419 6109
rect 21361 6069 21373 6103
rect 21407 6100 21419 6103
rect 21450 6100 21456 6112
rect 21407 6072 21456 6100
rect 21407 6069 21419 6072
rect 21361 6063 21419 6069
rect 21450 6060 21456 6072
rect 21508 6060 21514 6112
rect 22373 6103 22431 6109
rect 22373 6069 22385 6103
rect 22419 6100 22431 6103
rect 22848 6100 22876 6140
rect 23474 6128 23480 6140
rect 23532 6168 23538 6180
rect 23750 6168 23756 6180
rect 23532 6140 23756 6168
rect 23532 6128 23538 6140
rect 23750 6128 23756 6140
rect 23808 6128 23814 6180
rect 24504 6140 27568 6168
rect 22419 6072 22876 6100
rect 22419 6069 22431 6072
rect 22373 6063 22431 6069
rect 22922 6060 22928 6112
rect 22980 6060 22986 6112
rect 23014 6060 23020 6112
rect 23072 6100 23078 6112
rect 24504 6100 24532 6140
rect 23072 6072 24532 6100
rect 24857 6103 24915 6109
rect 23072 6060 23078 6072
rect 24857 6069 24869 6103
rect 24903 6100 24915 6103
rect 24946 6100 24952 6112
rect 24903 6072 24952 6100
rect 24903 6069 24915 6072
rect 24857 6063 24915 6069
rect 24946 6060 24952 6072
rect 25004 6060 25010 6112
rect 25038 6060 25044 6112
rect 25096 6060 25102 6112
rect 25498 6060 25504 6112
rect 25556 6060 25562 6112
rect 25682 6060 25688 6112
rect 25740 6100 25746 6112
rect 25777 6103 25835 6109
rect 25777 6100 25789 6103
rect 25740 6072 25789 6100
rect 25740 6060 25746 6072
rect 25777 6069 25789 6072
rect 25823 6069 25835 6103
rect 25777 6063 25835 6069
rect 25866 6060 25872 6112
rect 25924 6100 25930 6112
rect 26970 6100 26976 6112
rect 25924 6072 26976 6100
rect 25924 6060 25930 6072
rect 26970 6060 26976 6072
rect 27028 6060 27034 6112
rect 27154 6060 27160 6112
rect 27212 6060 27218 6112
rect 27540 6100 27568 6140
rect 28368 6140 28856 6168
rect 28368 6100 28396 6140
rect 27540 6072 28396 6100
rect 28626 6060 28632 6112
rect 28684 6100 28690 6112
rect 28721 6103 28779 6109
rect 28721 6100 28733 6103
rect 28684 6072 28733 6100
rect 28684 6060 28690 6072
rect 28721 6069 28733 6072
rect 28767 6069 28779 6103
rect 28828 6100 28856 6140
rect 29472 6140 30236 6168
rect 29472 6100 29500 6140
rect 28828 6072 29500 6100
rect 28721 6063 28779 6069
rect 29546 6060 29552 6112
rect 29604 6100 29610 6112
rect 30101 6103 30159 6109
rect 30101 6100 30113 6103
rect 29604 6072 30113 6100
rect 29604 6060 29610 6072
rect 30101 6069 30113 6072
rect 30147 6069 30159 6103
rect 30208 6100 30236 6140
rect 31036 6140 32444 6168
rect 31036 6100 31064 6140
rect 30208 6072 31064 6100
rect 30101 6063 30159 6069
rect 31294 6060 31300 6112
rect 31352 6100 31358 6112
rect 31757 6103 31815 6109
rect 31757 6100 31769 6103
rect 31352 6072 31769 6100
rect 31352 6060 31358 6072
rect 31757 6069 31769 6072
rect 31803 6069 31815 6103
rect 31757 6063 31815 6069
rect 32030 6060 32036 6112
rect 32088 6100 32094 6112
rect 32306 6100 32312 6112
rect 32088 6072 32312 6100
rect 32088 6060 32094 6072
rect 32306 6060 32312 6072
rect 32364 6060 32370 6112
rect 32416 6100 32444 6140
rect 33244 6100 33272 6208
rect 33873 6205 33885 6208
rect 33919 6205 33931 6239
rect 33873 6199 33931 6205
rect 33965 6239 34023 6245
rect 33965 6205 33977 6239
rect 34011 6205 34023 6239
rect 33965 6199 34023 6205
rect 33321 6171 33379 6177
rect 33321 6137 33333 6171
rect 33367 6168 33379 6171
rect 33980 6168 34008 6199
rect 34882 6196 34888 6248
rect 34940 6236 34946 6248
rect 34977 6239 35035 6245
rect 34977 6236 34989 6239
rect 34940 6208 34989 6236
rect 34940 6196 34946 6208
rect 34977 6205 34989 6208
rect 35023 6205 35035 6239
rect 34977 6199 35035 6205
rect 36262 6196 36268 6248
rect 36320 6236 36326 6248
rect 36541 6239 36599 6245
rect 36541 6236 36553 6239
rect 36320 6208 36553 6236
rect 36320 6196 36326 6208
rect 36541 6205 36553 6208
rect 36587 6205 36599 6239
rect 36541 6199 36599 6205
rect 36633 6239 36691 6245
rect 36633 6205 36645 6239
rect 36679 6205 36691 6239
rect 36633 6199 36691 6205
rect 33367 6140 34008 6168
rect 35989 6171 36047 6177
rect 33367 6137 33379 6140
rect 33321 6131 33379 6137
rect 35989 6137 36001 6171
rect 36035 6168 36047 6171
rect 36648 6168 36676 6199
rect 38470 6196 38476 6248
rect 38528 6236 38534 6248
rect 38672 6236 38700 6267
rect 38528 6208 38700 6236
rect 38528 6196 38534 6208
rect 36035 6140 36676 6168
rect 36035 6137 36047 6140
rect 35989 6131 36047 6137
rect 37550 6128 37556 6180
rect 37608 6168 37614 6180
rect 38381 6171 38439 6177
rect 38381 6168 38393 6171
rect 37608 6140 38393 6168
rect 37608 6128 37614 6140
rect 38381 6137 38393 6140
rect 38427 6137 38439 6171
rect 39025 6171 39083 6177
rect 39025 6168 39037 6171
rect 38381 6131 38439 6137
rect 38488 6140 39037 6168
rect 32416 6072 33272 6100
rect 33410 6060 33416 6112
rect 33468 6060 33474 6112
rect 35250 6060 35256 6112
rect 35308 6100 35314 6112
rect 38488 6100 38516 6140
rect 39025 6137 39037 6140
rect 39071 6137 39083 6171
rect 39025 6131 39083 6137
rect 35308 6072 38516 6100
rect 35308 6060 35314 6072
rect 38838 6060 38844 6112
rect 38896 6060 38902 6112
rect 1104 6010 39836 6032
rect 1104 5958 1950 6010
rect 2002 5958 2014 6010
rect 2066 5958 2078 6010
rect 2130 5958 2142 6010
rect 2194 5958 2206 6010
rect 2258 5958 7950 6010
rect 8002 5958 8014 6010
rect 8066 5958 8078 6010
rect 8130 5958 8142 6010
rect 8194 5958 8206 6010
rect 8258 5958 13950 6010
rect 14002 5958 14014 6010
rect 14066 5958 14078 6010
rect 14130 5958 14142 6010
rect 14194 5958 14206 6010
rect 14258 5958 19950 6010
rect 20002 5958 20014 6010
rect 20066 5958 20078 6010
rect 20130 5958 20142 6010
rect 20194 5958 20206 6010
rect 20258 5958 25950 6010
rect 26002 5958 26014 6010
rect 26066 5958 26078 6010
rect 26130 5958 26142 6010
rect 26194 5958 26206 6010
rect 26258 5958 31950 6010
rect 32002 5958 32014 6010
rect 32066 5958 32078 6010
rect 32130 5958 32142 6010
rect 32194 5958 32206 6010
rect 32258 5958 37950 6010
rect 38002 5958 38014 6010
rect 38066 5958 38078 6010
rect 38130 5958 38142 6010
rect 38194 5958 38206 6010
rect 38258 5958 39836 6010
rect 1104 5936 39836 5958
rect 2041 5899 2099 5905
rect 2041 5865 2053 5899
rect 2087 5896 2099 5899
rect 2498 5896 2504 5908
rect 2087 5868 2504 5896
rect 2087 5865 2099 5868
rect 2041 5859 2099 5865
rect 2498 5856 2504 5868
rect 2556 5856 2562 5908
rect 2593 5899 2651 5905
rect 2593 5865 2605 5899
rect 2639 5896 2651 5899
rect 3326 5896 3332 5908
rect 2639 5868 3332 5896
rect 2639 5865 2651 5868
rect 2593 5859 2651 5865
rect 3326 5856 3332 5868
rect 3384 5856 3390 5908
rect 4154 5856 4160 5908
rect 4212 5896 4218 5908
rect 4249 5899 4307 5905
rect 4249 5896 4261 5899
rect 4212 5868 4261 5896
rect 4212 5856 4218 5868
rect 4249 5865 4261 5868
rect 4295 5865 4307 5899
rect 4249 5859 4307 5865
rect 4614 5856 4620 5908
rect 4672 5896 4678 5908
rect 4672 5868 6408 5896
rect 4672 5856 4678 5868
rect 1765 5831 1823 5837
rect 1765 5797 1777 5831
rect 1811 5828 1823 5831
rect 2682 5828 2688 5840
rect 1811 5800 2688 5828
rect 1811 5797 1823 5800
rect 1765 5791 1823 5797
rect 2682 5788 2688 5800
rect 2740 5788 2746 5840
rect 3881 5831 3939 5837
rect 3881 5797 3893 5831
rect 3927 5828 3939 5831
rect 5074 5828 5080 5840
rect 3927 5800 5080 5828
rect 3927 5797 3939 5800
rect 3881 5791 3939 5797
rect 5074 5788 5080 5800
rect 5132 5788 5138 5840
rect 5828 5828 5856 5868
rect 5736 5800 5856 5828
rect 6380 5828 6408 5868
rect 6730 5856 6736 5908
rect 6788 5896 6794 5908
rect 7009 5899 7067 5905
rect 7009 5896 7021 5899
rect 6788 5868 7021 5896
rect 6788 5856 6794 5868
rect 7009 5865 7021 5868
rect 7055 5865 7067 5899
rect 7009 5859 7067 5865
rect 7374 5856 7380 5908
rect 7432 5896 7438 5908
rect 7561 5899 7619 5905
rect 7561 5896 7573 5899
rect 7432 5868 7573 5896
rect 7432 5856 7438 5868
rect 7561 5865 7573 5868
rect 7607 5865 7619 5899
rect 7561 5859 7619 5865
rect 7834 5856 7840 5908
rect 7892 5896 7898 5908
rect 8113 5899 8171 5905
rect 8113 5896 8125 5899
rect 7892 5868 8125 5896
rect 7892 5856 7898 5868
rect 8113 5865 8125 5868
rect 8159 5865 8171 5899
rect 8113 5859 8171 5865
rect 8386 5856 8392 5908
rect 8444 5856 8450 5908
rect 9306 5896 9312 5908
rect 8772 5868 9312 5896
rect 7190 5828 7196 5840
rect 6380 5800 7196 5828
rect 4706 5720 4712 5772
rect 4764 5760 4770 5772
rect 5442 5760 5448 5772
rect 4764 5732 5448 5760
rect 4764 5720 4770 5732
rect 5442 5720 5448 5732
rect 5500 5720 5506 5772
rect 5534 5720 5540 5772
rect 5592 5720 5598 5772
rect 5736 5769 5764 5800
rect 7190 5788 7196 5800
rect 7248 5788 7254 5840
rect 8404 5828 8432 5856
rect 7760 5800 8432 5828
rect 5721 5763 5779 5769
rect 5721 5729 5733 5763
rect 5767 5729 5779 5763
rect 5721 5723 5779 5729
rect 1026 5652 1032 5704
rect 1084 5692 1090 5704
rect 1949 5695 2007 5701
rect 1949 5692 1961 5695
rect 1084 5664 1961 5692
rect 1084 5652 1090 5664
rect 1949 5661 1961 5664
rect 1995 5661 2007 5695
rect 1949 5655 2007 5661
rect 2314 5652 2320 5704
rect 2372 5652 2378 5704
rect 2498 5652 2504 5704
rect 2556 5652 2562 5704
rect 3329 5695 3387 5701
rect 3329 5661 3341 5695
rect 3375 5661 3387 5695
rect 3329 5655 3387 5661
rect 3605 5695 3663 5701
rect 3605 5661 3617 5695
rect 3651 5661 3663 5695
rect 3605 5655 3663 5661
rect 382 5584 388 5636
rect 440 5624 446 5636
rect 1581 5627 1639 5633
rect 1581 5624 1593 5627
rect 440 5596 1593 5624
rect 440 5584 446 5596
rect 1581 5593 1593 5596
rect 1627 5593 1639 5627
rect 3344 5624 3372 5655
rect 3510 5624 3516 5636
rect 3344 5596 3516 5624
rect 1581 5587 1639 5593
rect 3510 5584 3516 5596
rect 3568 5584 3574 5636
rect 3620 5624 3648 5655
rect 3970 5652 3976 5704
rect 4028 5692 4034 5704
rect 4065 5695 4123 5701
rect 4065 5692 4077 5695
rect 4028 5664 4077 5692
rect 4028 5652 4034 5664
rect 4065 5661 4077 5664
rect 4111 5661 4123 5695
rect 4065 5655 4123 5661
rect 4433 5695 4491 5701
rect 4433 5661 4445 5695
rect 4479 5692 4491 5695
rect 4522 5692 4528 5704
rect 4479 5664 4528 5692
rect 4479 5661 4491 5664
rect 4433 5655 4491 5661
rect 4522 5652 4528 5664
rect 4580 5652 4586 5704
rect 4801 5695 4859 5701
rect 4801 5661 4813 5695
rect 4847 5692 4859 5695
rect 5261 5695 5319 5701
rect 5261 5692 5273 5695
rect 4847 5664 5273 5692
rect 4847 5661 4859 5664
rect 4801 5655 4859 5661
rect 5261 5661 5273 5664
rect 5307 5692 5319 5695
rect 5350 5692 5356 5704
rect 5307 5664 5356 5692
rect 5307 5661 5319 5664
rect 5261 5655 5319 5661
rect 5350 5652 5356 5664
rect 5408 5652 5414 5704
rect 5902 5652 5908 5704
rect 5960 5692 5966 5704
rect 5997 5695 6055 5701
rect 5997 5692 6009 5695
rect 5960 5664 6009 5692
rect 5960 5652 5966 5664
rect 5997 5661 6009 5664
rect 6043 5661 6055 5695
rect 5997 5655 6055 5661
rect 7193 5695 7251 5701
rect 7193 5661 7205 5695
rect 7239 5692 7251 5695
rect 7282 5692 7288 5704
rect 7239 5664 7288 5692
rect 7239 5661 7251 5664
rect 7193 5655 7251 5661
rect 7282 5652 7288 5664
rect 7340 5652 7346 5704
rect 7760 5701 7788 5800
rect 8389 5763 8447 5769
rect 8389 5760 8401 5763
rect 8220 5732 8401 5760
rect 7745 5695 7803 5701
rect 7745 5661 7757 5695
rect 7791 5661 7803 5695
rect 7745 5655 7803 5661
rect 4614 5624 4620 5636
rect 3620 5596 4620 5624
rect 4614 5584 4620 5596
rect 4672 5584 4678 5636
rect 5810 5624 5816 5636
rect 4816 5596 5816 5624
rect 2498 5516 2504 5568
rect 2556 5556 2562 5568
rect 4816 5556 4844 5596
rect 5810 5584 5816 5596
rect 5868 5584 5874 5636
rect 7466 5584 7472 5636
rect 7524 5624 7530 5636
rect 8220 5624 8248 5732
rect 8389 5729 8401 5732
rect 8435 5760 8447 5763
rect 8772 5760 8800 5868
rect 9306 5856 9312 5868
rect 9364 5856 9370 5908
rect 10410 5856 10416 5908
rect 10468 5856 10474 5908
rect 10686 5856 10692 5908
rect 10744 5896 10750 5908
rect 13814 5896 13820 5908
rect 10744 5868 13820 5896
rect 10744 5856 10750 5868
rect 13814 5856 13820 5868
rect 13872 5856 13878 5908
rect 14093 5899 14151 5905
rect 14093 5865 14105 5899
rect 14139 5896 14151 5899
rect 14274 5896 14280 5908
rect 14139 5868 14280 5896
rect 14139 5865 14151 5868
rect 14093 5859 14151 5865
rect 14274 5856 14280 5868
rect 14332 5856 14338 5908
rect 15102 5856 15108 5908
rect 15160 5896 15166 5908
rect 15160 5868 15516 5896
rect 15160 5856 15166 5868
rect 8435 5732 8800 5760
rect 8435 5729 8447 5732
rect 8389 5723 8447 5729
rect 8846 5720 8852 5772
rect 8904 5760 8910 5772
rect 9033 5763 9091 5769
rect 9033 5760 9045 5763
rect 8904 5732 9045 5760
rect 8904 5720 8910 5732
rect 9033 5729 9045 5732
rect 9079 5729 9091 5763
rect 10428 5760 10456 5856
rect 10870 5788 10876 5840
rect 10928 5828 10934 5840
rect 14458 5828 14464 5840
rect 10928 5800 14464 5828
rect 10928 5788 10934 5800
rect 14458 5788 14464 5800
rect 14516 5788 14522 5840
rect 15488 5828 15516 5868
rect 15562 5856 15568 5908
rect 15620 5856 15626 5908
rect 15930 5856 15936 5908
rect 15988 5896 15994 5908
rect 15988 5868 17264 5896
rect 15988 5856 15994 5868
rect 16206 5828 16212 5840
rect 15488 5800 16212 5828
rect 16206 5788 16212 5800
rect 16264 5788 16270 5840
rect 16298 5788 16304 5840
rect 16356 5788 16362 5840
rect 17236 5828 17264 5868
rect 17310 5856 17316 5908
rect 17368 5856 17374 5908
rect 17586 5856 17592 5908
rect 17644 5896 17650 5908
rect 17681 5899 17739 5905
rect 17681 5896 17693 5899
rect 17644 5868 17693 5896
rect 17644 5856 17650 5868
rect 17681 5865 17693 5868
rect 17727 5865 17739 5899
rect 17681 5859 17739 5865
rect 17788 5868 20300 5896
rect 17788 5828 17816 5868
rect 18506 5828 18512 5840
rect 17236 5800 17816 5828
rect 17880 5800 18512 5828
rect 11057 5763 11115 5769
rect 11057 5760 11069 5763
rect 10428 5732 11069 5760
rect 9033 5723 9091 5729
rect 11057 5729 11069 5732
rect 11103 5729 11115 5763
rect 13078 5760 13084 5772
rect 11057 5723 11115 5729
rect 11164 5732 13084 5760
rect 8297 5695 8355 5701
rect 8297 5661 8309 5695
rect 8343 5661 8355 5695
rect 8297 5655 8355 5661
rect 8573 5695 8631 5701
rect 8573 5661 8585 5695
rect 8619 5692 8631 5695
rect 9674 5692 9680 5704
rect 8619 5664 9680 5692
rect 8619 5661 8631 5664
rect 8573 5655 8631 5661
rect 7524 5596 8248 5624
rect 8312 5624 8340 5655
rect 9674 5652 9680 5664
rect 9732 5692 9738 5704
rect 11164 5692 11192 5732
rect 13078 5720 13084 5732
rect 13136 5720 13142 5772
rect 16316 5760 16344 5788
rect 15948 5732 16344 5760
rect 9732 5664 11192 5692
rect 9732 5652 9738 5664
rect 11422 5652 11428 5704
rect 11480 5652 11486 5704
rect 11606 5652 11612 5704
rect 11664 5652 11670 5704
rect 11701 5695 11759 5701
rect 11701 5661 11713 5695
rect 11747 5661 11759 5695
rect 11701 5655 11759 5661
rect 11793 5695 11851 5701
rect 11793 5661 11805 5695
rect 11839 5692 11851 5695
rect 12250 5692 12256 5704
rect 11839 5664 12256 5692
rect 11839 5661 11851 5664
rect 11793 5655 11851 5661
rect 8662 5624 8668 5636
rect 8312 5596 8668 5624
rect 7524 5584 7530 5596
rect 8662 5584 8668 5596
rect 8720 5584 8726 5636
rect 8757 5627 8815 5633
rect 8757 5593 8769 5627
rect 8803 5624 8815 5627
rect 9278 5627 9336 5633
rect 9278 5624 9290 5627
rect 8803 5596 9290 5624
rect 8803 5593 8815 5596
rect 8757 5587 8815 5593
rect 9278 5593 9290 5596
rect 9324 5624 9336 5627
rect 10318 5624 10324 5636
rect 9324 5596 10324 5624
rect 9324 5593 9336 5596
rect 9278 5587 9336 5593
rect 10318 5584 10324 5596
rect 10376 5584 10382 5636
rect 11330 5584 11336 5636
rect 11388 5624 11394 5636
rect 11716 5624 11744 5655
rect 12250 5652 12256 5664
rect 12308 5652 12314 5704
rect 13630 5652 13636 5704
rect 13688 5692 13694 5704
rect 13909 5695 13967 5701
rect 13909 5692 13921 5695
rect 13688 5664 13921 5692
rect 13688 5652 13694 5664
rect 13909 5661 13921 5664
rect 13955 5661 13967 5695
rect 13909 5655 13967 5661
rect 15470 5652 15476 5704
rect 15528 5652 15534 5704
rect 15654 5652 15660 5704
rect 15712 5692 15718 5704
rect 15948 5701 15976 5732
rect 15841 5695 15899 5701
rect 15841 5692 15853 5695
rect 15712 5664 15853 5692
rect 15712 5652 15718 5664
rect 15841 5661 15853 5664
rect 15887 5661 15899 5695
rect 15841 5655 15899 5661
rect 15933 5695 15991 5701
rect 15933 5661 15945 5695
rect 15979 5661 15991 5695
rect 15933 5655 15991 5661
rect 11388 5596 11744 5624
rect 11388 5584 11394 5596
rect 12066 5584 12072 5636
rect 12124 5584 12130 5636
rect 12158 5584 12164 5636
rect 12216 5584 12222 5636
rect 15102 5624 15108 5636
rect 12268 5596 15108 5624
rect 2556 5528 4844 5556
rect 4893 5559 4951 5565
rect 2556 5516 2562 5528
rect 4893 5525 4905 5559
rect 4939 5556 4951 5559
rect 5166 5556 5172 5568
rect 4939 5528 5172 5556
rect 4939 5525 4951 5528
rect 4893 5519 4951 5525
rect 5166 5516 5172 5528
rect 5224 5516 5230 5568
rect 5350 5516 5356 5568
rect 5408 5516 5414 5568
rect 6546 5516 6552 5568
rect 6604 5556 6610 5568
rect 6733 5559 6791 5565
rect 6733 5556 6745 5559
rect 6604 5528 6745 5556
rect 6604 5516 6610 5528
rect 6733 5525 6745 5528
rect 6779 5525 6791 5559
rect 6733 5519 6791 5525
rect 8294 5516 8300 5568
rect 8352 5556 8358 5568
rect 10505 5559 10563 5565
rect 10505 5556 10517 5559
rect 8352 5528 10517 5556
rect 8352 5516 8358 5528
rect 10505 5525 10517 5528
rect 10551 5525 10563 5559
rect 10505 5519 10563 5525
rect 11422 5516 11428 5568
rect 11480 5556 11486 5568
rect 12268 5556 12296 5596
rect 15102 5584 15108 5596
rect 15160 5584 15166 5636
rect 15228 5627 15286 5633
rect 15228 5593 15240 5627
rect 15274 5624 15286 5627
rect 15948 5624 15976 5655
rect 16022 5652 16028 5704
rect 16080 5652 16086 5704
rect 16206 5652 16212 5704
rect 16264 5652 16270 5704
rect 16301 5695 16359 5701
rect 16301 5661 16313 5695
rect 16347 5692 16359 5695
rect 16347 5664 16436 5692
rect 16347 5661 16359 5664
rect 16301 5655 16359 5661
rect 15274 5596 15976 5624
rect 16408 5624 16436 5664
rect 16574 5652 16580 5704
rect 16632 5652 16638 5704
rect 17497 5695 17555 5701
rect 17497 5661 17509 5695
rect 17543 5692 17555 5695
rect 17770 5692 17776 5704
rect 17543 5664 17776 5692
rect 17543 5661 17555 5664
rect 17497 5655 17555 5661
rect 17770 5652 17776 5664
rect 17828 5652 17834 5704
rect 16666 5624 16672 5636
rect 16408 5596 16672 5624
rect 15274 5593 15286 5596
rect 15228 5587 15286 5593
rect 16666 5584 16672 5596
rect 16724 5584 16730 5636
rect 17880 5624 17908 5800
rect 18506 5788 18512 5800
rect 18564 5788 18570 5840
rect 17957 5763 18015 5769
rect 17957 5729 17969 5763
rect 18003 5760 18015 5763
rect 18414 5760 18420 5772
rect 18003 5732 18420 5760
rect 18003 5729 18015 5732
rect 17957 5723 18015 5729
rect 18414 5720 18420 5732
rect 18472 5720 18478 5772
rect 18874 5720 18880 5772
rect 18932 5760 18938 5772
rect 19245 5763 19303 5769
rect 19245 5760 19257 5763
rect 18932 5732 19257 5760
rect 18932 5720 18938 5732
rect 19245 5729 19257 5732
rect 19291 5729 19303 5763
rect 20272 5760 20300 5868
rect 20714 5856 20720 5908
rect 20772 5896 20778 5908
rect 24486 5896 24492 5908
rect 20772 5868 24492 5896
rect 20772 5856 20778 5868
rect 24486 5856 24492 5868
rect 24544 5856 24550 5908
rect 26510 5856 26516 5908
rect 26568 5896 26574 5908
rect 27154 5896 27160 5908
rect 26568 5868 27160 5896
rect 26568 5856 26574 5868
rect 27154 5856 27160 5868
rect 27212 5856 27218 5908
rect 27890 5856 27896 5908
rect 27948 5896 27954 5908
rect 28169 5899 28227 5905
rect 28169 5896 28181 5899
rect 27948 5868 28181 5896
rect 27948 5856 27954 5868
rect 28169 5865 28181 5868
rect 28215 5865 28227 5899
rect 28169 5859 28227 5865
rect 28258 5856 28264 5908
rect 28316 5896 28322 5908
rect 29546 5896 29552 5908
rect 28316 5868 29552 5896
rect 28316 5856 28322 5868
rect 29546 5856 29552 5868
rect 29604 5856 29610 5908
rect 30009 5899 30067 5905
rect 30009 5865 30021 5899
rect 30055 5896 30067 5899
rect 30055 5868 31156 5896
rect 30055 5865 30067 5868
rect 30009 5859 30067 5865
rect 23106 5788 23112 5840
rect 23164 5788 23170 5840
rect 24026 5788 24032 5840
rect 24084 5788 24090 5840
rect 24210 5788 24216 5840
rect 24268 5828 24274 5840
rect 27065 5831 27123 5837
rect 24268 5800 24624 5828
rect 24268 5788 24274 5800
rect 24596 5772 24624 5800
rect 27065 5797 27077 5831
rect 27111 5828 27123 5831
rect 28074 5828 28080 5840
rect 27111 5800 28080 5828
rect 27111 5797 27123 5800
rect 27065 5791 27123 5797
rect 28074 5788 28080 5800
rect 28132 5788 28138 5840
rect 28629 5831 28687 5837
rect 28629 5797 28641 5831
rect 28675 5828 28687 5831
rect 29178 5828 29184 5840
rect 28675 5800 29184 5828
rect 28675 5797 28687 5800
rect 28629 5791 28687 5797
rect 29178 5788 29184 5800
rect 29236 5788 29242 5840
rect 29365 5831 29423 5837
rect 29365 5797 29377 5831
rect 29411 5828 29423 5831
rect 30190 5828 30196 5840
rect 29411 5800 30196 5828
rect 29411 5797 29423 5800
rect 29365 5791 29423 5797
rect 30190 5788 30196 5800
rect 30248 5788 30254 5840
rect 31128 5828 31156 5868
rect 31202 5856 31208 5908
rect 31260 5856 31266 5908
rect 32217 5899 32275 5905
rect 32217 5865 32229 5899
rect 32263 5896 32275 5899
rect 36630 5896 36636 5908
rect 32263 5868 36636 5896
rect 32263 5865 32275 5868
rect 32217 5859 32275 5865
rect 36630 5856 36636 5868
rect 36688 5856 36694 5908
rect 36814 5856 36820 5908
rect 36872 5896 36878 5908
rect 37461 5899 37519 5905
rect 37461 5896 37473 5899
rect 36872 5868 37473 5896
rect 36872 5856 36878 5868
rect 37461 5865 37473 5868
rect 37507 5865 37519 5899
rect 37461 5859 37519 5865
rect 37826 5856 37832 5908
rect 37884 5896 37890 5908
rect 37921 5899 37979 5905
rect 37921 5896 37933 5899
rect 37884 5868 37933 5896
rect 37884 5856 37890 5868
rect 37921 5865 37933 5868
rect 37967 5865 37979 5899
rect 37921 5859 37979 5865
rect 34146 5828 34152 5840
rect 31128 5800 34152 5828
rect 34146 5788 34152 5800
rect 34204 5788 34210 5840
rect 36354 5788 36360 5840
rect 36412 5828 36418 5840
rect 38565 5831 38623 5837
rect 38565 5828 38577 5831
rect 36412 5800 38577 5828
rect 36412 5788 36418 5800
rect 38565 5797 38577 5800
rect 38611 5797 38623 5831
rect 38565 5791 38623 5797
rect 39390 5788 39396 5840
rect 39448 5788 39454 5840
rect 21269 5763 21327 5769
rect 21269 5760 21281 5763
rect 20272 5732 21281 5760
rect 19245 5723 19303 5729
rect 21269 5729 21281 5732
rect 21315 5729 21327 5763
rect 21913 5763 21971 5769
rect 21913 5760 21925 5763
rect 21269 5723 21327 5729
rect 21376 5732 21925 5760
rect 18141 5695 18199 5701
rect 18141 5661 18153 5695
rect 18187 5692 18199 5695
rect 18322 5692 18328 5704
rect 18187 5664 18328 5692
rect 18187 5661 18199 5664
rect 18141 5655 18199 5661
rect 18322 5652 18328 5664
rect 18380 5652 18386 5704
rect 18782 5652 18788 5704
rect 18840 5652 18846 5704
rect 19061 5695 19119 5701
rect 19061 5661 19073 5695
rect 19107 5661 19119 5695
rect 19061 5655 19119 5661
rect 19076 5624 19104 5655
rect 19334 5652 19340 5704
rect 19392 5692 19398 5704
rect 19501 5695 19559 5701
rect 19501 5692 19513 5695
rect 19392 5664 19513 5692
rect 19392 5652 19398 5664
rect 19501 5661 19513 5664
rect 19547 5661 19559 5695
rect 19501 5655 19559 5661
rect 21084 5695 21142 5701
rect 21084 5661 21096 5695
rect 21130 5661 21142 5695
rect 21084 5655 21142 5661
rect 21177 5695 21235 5701
rect 21177 5661 21189 5695
rect 21223 5692 21235 5695
rect 21376 5692 21404 5732
rect 21913 5729 21925 5732
rect 21959 5760 21971 5763
rect 22002 5760 22008 5772
rect 21959 5732 22008 5760
rect 21959 5729 21971 5732
rect 21913 5723 21971 5729
rect 22002 5720 22008 5732
rect 22060 5720 22066 5772
rect 22278 5720 22284 5772
rect 22336 5769 22342 5772
rect 22336 5763 22364 5769
rect 22352 5729 22364 5763
rect 22646 5760 22652 5772
rect 22336 5723 22364 5729
rect 22404 5732 22652 5760
rect 22336 5720 22342 5723
rect 21223 5664 21404 5692
rect 21453 5695 21511 5701
rect 21223 5661 21235 5664
rect 21177 5655 21235 5661
rect 21453 5661 21465 5695
rect 21499 5692 21511 5695
rect 21634 5692 21640 5704
rect 21499 5664 21640 5692
rect 21499 5661 21511 5664
rect 21453 5655 21511 5661
rect 19702 5624 19708 5636
rect 16776 5596 17908 5624
rect 17972 5596 18644 5624
rect 19076 5596 19708 5624
rect 11480 5528 12296 5556
rect 11480 5516 11486 5528
rect 12342 5516 12348 5568
rect 12400 5556 12406 5568
rect 16776 5556 16804 5596
rect 12400 5528 16804 5556
rect 12400 5516 12406 5528
rect 16942 5516 16948 5568
rect 17000 5556 17006 5568
rect 17126 5556 17132 5568
rect 17000 5528 17132 5556
rect 17000 5516 17006 5528
rect 17126 5516 17132 5528
rect 17184 5516 17190 5568
rect 17770 5516 17776 5568
rect 17828 5556 17834 5568
rect 17972 5556 18000 5596
rect 17828 5528 18000 5556
rect 18049 5559 18107 5565
rect 17828 5516 17834 5528
rect 18049 5525 18061 5559
rect 18095 5556 18107 5559
rect 18322 5556 18328 5568
rect 18095 5528 18328 5556
rect 18095 5525 18107 5528
rect 18049 5519 18107 5525
rect 18322 5516 18328 5528
rect 18380 5516 18386 5568
rect 18506 5516 18512 5568
rect 18564 5516 18570 5568
rect 18616 5565 18644 5596
rect 19702 5584 19708 5596
rect 19760 5584 19766 5636
rect 21100 5624 21128 5655
rect 21634 5652 21640 5664
rect 21692 5652 21698 5704
rect 22189 5695 22247 5701
rect 22189 5661 22201 5695
rect 22235 5692 22247 5695
rect 22404 5692 22432 5732
rect 22646 5720 22652 5732
rect 22704 5720 22710 5772
rect 24578 5720 24584 5772
rect 24636 5760 24642 5772
rect 24857 5763 24915 5769
rect 24857 5760 24869 5763
rect 24636 5732 24869 5760
rect 24636 5720 24642 5732
rect 24857 5729 24869 5732
rect 24903 5729 24915 5763
rect 24857 5723 24915 5729
rect 24946 5720 24952 5772
rect 25004 5720 25010 5772
rect 27430 5720 27436 5772
rect 27488 5760 27494 5772
rect 27709 5763 27767 5769
rect 27709 5760 27721 5763
rect 27488 5732 27721 5760
rect 27488 5720 27494 5732
rect 27709 5729 27721 5732
rect 27755 5729 27767 5763
rect 28905 5763 28963 5769
rect 28905 5760 28917 5763
rect 27709 5723 27767 5729
rect 28644 5732 28917 5760
rect 28644 5704 28672 5732
rect 28905 5729 28917 5732
rect 28951 5729 28963 5763
rect 28905 5723 28963 5729
rect 29270 5720 29276 5772
rect 29328 5760 29334 5772
rect 29328 5732 29868 5760
rect 29328 5720 29334 5732
rect 22235 5664 22432 5692
rect 22235 5661 22247 5664
rect 22189 5655 22247 5661
rect 22462 5652 22468 5704
rect 22520 5652 22526 5704
rect 23106 5652 23112 5704
rect 23164 5692 23170 5704
rect 23385 5695 23443 5701
rect 23385 5692 23397 5695
rect 23164 5664 23397 5692
rect 23164 5652 23170 5664
rect 23385 5661 23397 5664
rect 23431 5661 23443 5695
rect 23385 5655 23443 5661
rect 24213 5695 24271 5701
rect 24213 5661 24225 5695
rect 24259 5692 24271 5695
rect 24394 5692 24400 5704
rect 24259 5664 24400 5692
rect 24259 5661 24271 5664
rect 24213 5655 24271 5661
rect 24394 5652 24400 5664
rect 24452 5652 24458 5704
rect 24762 5652 24768 5704
rect 24820 5692 24826 5704
rect 25866 5692 25872 5704
rect 24820 5664 25872 5692
rect 24820 5652 24826 5664
rect 25866 5652 25872 5664
rect 25924 5652 25930 5704
rect 26326 5652 26332 5704
rect 26384 5692 26390 5704
rect 28353 5695 28411 5701
rect 26384 5668 26740 5692
rect 26881 5671 26939 5677
rect 26881 5668 26893 5671
rect 26384 5664 26893 5668
rect 26384 5652 26390 5664
rect 26712 5640 26893 5664
rect 26881 5637 26893 5640
rect 26927 5637 26939 5671
rect 28353 5661 28365 5695
rect 28399 5661 28411 5695
rect 28353 5655 28411 5661
rect 28445 5695 28503 5701
rect 28445 5661 28457 5695
rect 28491 5661 28503 5695
rect 28445 5655 28503 5661
rect 21358 5624 21364 5636
rect 21100 5596 21364 5624
rect 21358 5584 21364 5596
rect 21416 5584 21422 5636
rect 23750 5624 23756 5636
rect 22940 5596 23756 5624
rect 18601 5559 18659 5565
rect 18601 5525 18613 5559
rect 18647 5525 18659 5559
rect 18601 5519 18659 5525
rect 18782 5516 18788 5568
rect 18840 5556 18846 5568
rect 18877 5559 18935 5565
rect 18877 5556 18889 5559
rect 18840 5528 18889 5556
rect 18840 5516 18846 5528
rect 18877 5525 18889 5528
rect 18923 5525 18935 5559
rect 18877 5519 18935 5525
rect 19058 5516 19064 5568
rect 19116 5556 19122 5568
rect 20625 5559 20683 5565
rect 20625 5556 20637 5559
rect 19116 5528 20637 5556
rect 19116 5516 19122 5528
rect 20625 5525 20637 5528
rect 20671 5525 20683 5559
rect 20625 5519 20683 5525
rect 20809 5559 20867 5565
rect 20809 5525 20821 5559
rect 20855 5556 20867 5559
rect 21450 5556 21456 5568
rect 20855 5528 21456 5556
rect 20855 5525 20867 5528
rect 20809 5519 20867 5525
rect 21450 5516 21456 5528
rect 21508 5516 21514 5568
rect 22002 5516 22008 5568
rect 22060 5556 22066 5568
rect 22940 5556 22968 5596
rect 23750 5584 23756 5596
rect 23808 5584 23814 5636
rect 23934 5584 23940 5636
rect 23992 5624 23998 5636
rect 26881 5631 26939 5637
rect 27525 5627 27583 5633
rect 27525 5624 27537 5627
rect 23992 5596 26648 5624
rect 23992 5584 23998 5596
rect 22060 5528 22968 5556
rect 22060 5516 22066 5528
rect 23198 5516 23204 5568
rect 23256 5516 23262 5568
rect 23566 5516 23572 5568
rect 23624 5556 23630 5568
rect 24210 5556 24216 5568
rect 23624 5528 24216 5556
rect 23624 5516 23630 5528
rect 24210 5516 24216 5528
rect 24268 5516 24274 5568
rect 24394 5516 24400 5568
rect 24452 5516 24458 5568
rect 24854 5516 24860 5568
rect 24912 5556 24918 5568
rect 26418 5556 26424 5568
rect 24912 5528 26424 5556
rect 24912 5516 24918 5528
rect 26418 5516 26424 5528
rect 26476 5516 26482 5568
rect 26620 5556 26648 5596
rect 26988 5596 27537 5624
rect 26988 5556 27016 5596
rect 27525 5593 27537 5596
rect 27571 5624 27583 5627
rect 28258 5624 28264 5636
rect 27571 5596 28264 5624
rect 27571 5593 27583 5596
rect 27525 5587 27583 5593
rect 28258 5584 28264 5596
rect 28316 5584 28322 5636
rect 26620 5528 27016 5556
rect 27157 5559 27215 5565
rect 27157 5525 27169 5559
rect 27203 5556 27215 5559
rect 27338 5556 27344 5568
rect 27203 5528 27344 5556
rect 27203 5525 27215 5528
rect 27157 5519 27215 5525
rect 27338 5516 27344 5528
rect 27396 5516 27402 5568
rect 27614 5516 27620 5568
rect 27672 5516 27678 5568
rect 28368 5556 28396 5655
rect 28460 5624 28488 5655
rect 28626 5652 28632 5704
rect 28684 5652 28690 5704
rect 28718 5652 28724 5704
rect 28776 5652 28782 5704
rect 28994 5652 29000 5704
rect 29052 5652 29058 5704
rect 29086 5652 29092 5704
rect 29144 5692 29150 5704
rect 29840 5701 29868 5732
rect 30760 5732 32076 5760
rect 30760 5704 30788 5732
rect 32048 5704 32076 5732
rect 32950 5720 32956 5772
rect 33008 5760 33014 5772
rect 34606 5760 34612 5772
rect 33008 5732 34612 5760
rect 33008 5720 33014 5732
rect 34606 5720 34612 5732
rect 34664 5720 34670 5772
rect 34790 5720 34796 5772
rect 34848 5720 34854 5772
rect 37274 5720 37280 5772
rect 37332 5760 37338 5772
rect 37332 5732 38792 5760
rect 37332 5720 37338 5732
rect 29733 5695 29791 5701
rect 29733 5692 29745 5695
rect 29144 5664 29745 5692
rect 29144 5652 29150 5664
rect 29733 5661 29745 5664
rect 29779 5661 29791 5695
rect 29733 5655 29791 5661
rect 29825 5695 29883 5701
rect 29825 5661 29837 5695
rect 29871 5661 29883 5695
rect 29825 5655 29883 5661
rect 30006 5652 30012 5704
rect 30064 5692 30070 5704
rect 30193 5695 30251 5701
rect 30193 5692 30205 5695
rect 30064 5664 30205 5692
rect 30064 5652 30070 5664
rect 30193 5661 30205 5664
rect 30239 5661 30251 5695
rect 30193 5655 30251 5661
rect 30374 5652 30380 5704
rect 30432 5692 30438 5704
rect 30469 5695 30527 5701
rect 30469 5692 30481 5695
rect 30432 5664 30481 5692
rect 30432 5652 30438 5664
rect 30469 5661 30481 5664
rect 30515 5692 30527 5695
rect 30742 5692 30748 5704
rect 30515 5664 30748 5692
rect 30515 5661 30527 5664
rect 30469 5655 30527 5661
rect 30742 5652 30748 5664
rect 30800 5652 30806 5704
rect 31765 5695 31823 5701
rect 31765 5661 31777 5695
rect 31811 5692 31823 5695
rect 31811 5664 31892 5692
rect 31811 5661 31823 5664
rect 31765 5655 31823 5661
rect 29638 5624 29644 5636
rect 28460 5596 29644 5624
rect 29638 5584 29644 5596
rect 29696 5584 29702 5636
rect 30650 5584 30656 5636
rect 30708 5624 30714 5636
rect 31864 5624 31892 5664
rect 32030 5652 32036 5704
rect 32088 5652 32094 5704
rect 32214 5652 32220 5704
rect 32272 5692 32278 5704
rect 32272 5664 33364 5692
rect 32272 5652 32278 5664
rect 30708 5596 31892 5624
rect 33336 5624 33364 5664
rect 33410 5652 33416 5704
rect 33468 5652 33474 5704
rect 34514 5652 34520 5704
rect 34572 5692 34578 5704
rect 35069 5695 35127 5701
rect 35069 5692 35081 5695
rect 34572 5688 34744 5692
rect 34808 5688 35081 5692
rect 34572 5664 35081 5688
rect 34572 5652 34578 5664
rect 34716 5660 34836 5664
rect 35069 5661 35081 5664
rect 35115 5661 35127 5695
rect 35069 5655 35127 5661
rect 35526 5652 35532 5704
rect 35584 5692 35590 5704
rect 37645 5695 37703 5701
rect 37645 5692 37657 5695
rect 35584 5664 36676 5692
rect 35584 5652 35590 5664
rect 33336 5596 35848 5624
rect 30708 5584 30714 5596
rect 28994 5556 29000 5568
rect 28368 5528 29000 5556
rect 28994 5516 29000 5528
rect 29052 5516 29058 5568
rect 29546 5516 29552 5568
rect 29604 5516 29610 5568
rect 31941 5559 31999 5565
rect 31941 5525 31953 5559
rect 31987 5556 31999 5559
rect 32950 5556 32956 5568
rect 31987 5528 32956 5556
rect 31987 5525 31999 5528
rect 31941 5519 31999 5525
rect 32950 5516 32956 5528
rect 33008 5516 33014 5568
rect 33226 5516 33232 5568
rect 33284 5516 33290 5568
rect 34790 5516 34796 5568
rect 34848 5556 34854 5568
rect 35526 5556 35532 5568
rect 34848 5528 35532 5556
rect 34848 5516 34854 5528
rect 35526 5516 35532 5528
rect 35584 5516 35590 5568
rect 35820 5565 35848 5596
rect 35805 5559 35863 5565
rect 35805 5525 35817 5559
rect 35851 5525 35863 5559
rect 36648 5556 36676 5664
rect 37292 5664 37657 5692
rect 37292 5636 37320 5664
rect 37645 5661 37657 5664
rect 37691 5661 37703 5695
rect 37645 5655 37703 5661
rect 37737 5695 37795 5701
rect 37737 5661 37749 5695
rect 37783 5661 37795 5695
rect 37737 5655 37795 5661
rect 38473 5695 38531 5701
rect 38473 5661 38485 5695
rect 38519 5692 38531 5695
rect 38562 5692 38568 5704
rect 38519 5664 38568 5692
rect 38519 5661 38531 5664
rect 38473 5655 38531 5661
rect 37274 5584 37280 5636
rect 37332 5584 37338 5636
rect 37550 5584 37556 5636
rect 37608 5624 37614 5636
rect 37752 5624 37780 5655
rect 38562 5652 38568 5664
rect 38620 5652 38626 5704
rect 38764 5701 38792 5732
rect 38749 5695 38807 5701
rect 38749 5661 38761 5695
rect 38795 5661 38807 5695
rect 38749 5655 38807 5661
rect 38841 5695 38899 5701
rect 38841 5661 38853 5695
rect 38887 5661 38899 5695
rect 38841 5655 38899 5661
rect 37608 5596 37780 5624
rect 38856 5624 38884 5655
rect 39206 5652 39212 5704
rect 39264 5652 39270 5704
rect 39758 5624 39764 5636
rect 38856 5596 39764 5624
rect 37608 5584 37614 5596
rect 39758 5584 39764 5596
rect 39816 5584 39822 5636
rect 38289 5559 38347 5565
rect 38289 5556 38301 5559
rect 36648 5528 38301 5556
rect 35805 5519 35863 5525
rect 38289 5525 38301 5528
rect 38335 5525 38347 5559
rect 38289 5519 38347 5525
rect 39025 5559 39083 5565
rect 39025 5525 39037 5559
rect 39071 5556 39083 5559
rect 39942 5556 39948 5568
rect 39071 5528 39948 5556
rect 39071 5525 39083 5528
rect 39025 5519 39083 5525
rect 39942 5516 39948 5528
rect 40000 5516 40006 5568
rect 1104 5466 39836 5488
rect 1104 5414 3010 5466
rect 3062 5414 3074 5466
rect 3126 5414 3138 5466
rect 3190 5414 3202 5466
rect 3254 5414 3266 5466
rect 3318 5414 9010 5466
rect 9062 5414 9074 5466
rect 9126 5414 9138 5466
rect 9190 5414 9202 5466
rect 9254 5414 9266 5466
rect 9318 5414 15010 5466
rect 15062 5414 15074 5466
rect 15126 5414 15138 5466
rect 15190 5414 15202 5466
rect 15254 5414 15266 5466
rect 15318 5414 21010 5466
rect 21062 5414 21074 5466
rect 21126 5414 21138 5466
rect 21190 5414 21202 5466
rect 21254 5414 21266 5466
rect 21318 5414 27010 5466
rect 27062 5414 27074 5466
rect 27126 5414 27138 5466
rect 27190 5414 27202 5466
rect 27254 5414 27266 5466
rect 27318 5414 33010 5466
rect 33062 5414 33074 5466
rect 33126 5414 33138 5466
rect 33190 5414 33202 5466
rect 33254 5414 33266 5466
rect 33318 5414 39010 5466
rect 39062 5414 39074 5466
rect 39126 5414 39138 5466
rect 39190 5414 39202 5466
rect 39254 5414 39266 5466
rect 39318 5414 39836 5466
rect 1104 5392 39836 5414
rect 1486 5312 1492 5364
rect 1544 5352 1550 5364
rect 1762 5352 1768 5364
rect 1544 5324 1768 5352
rect 1544 5312 1550 5324
rect 1762 5312 1768 5324
rect 1820 5312 1826 5364
rect 2041 5355 2099 5361
rect 2041 5321 2053 5355
rect 2087 5321 2099 5355
rect 2041 5315 2099 5321
rect 1210 5244 1216 5296
rect 1268 5284 1274 5296
rect 2056 5284 2084 5315
rect 2774 5312 2780 5364
rect 2832 5352 2838 5364
rect 3053 5355 3111 5361
rect 3053 5352 3065 5355
rect 2832 5324 3065 5352
rect 2832 5312 2838 5324
rect 3053 5321 3065 5324
rect 3099 5321 3111 5355
rect 5902 5352 5908 5364
rect 3053 5315 3111 5321
rect 3160 5324 5908 5352
rect 3160 5284 3188 5324
rect 5902 5312 5908 5324
rect 5960 5312 5966 5364
rect 5997 5355 6055 5361
rect 5997 5321 6009 5355
rect 6043 5352 6055 5355
rect 6270 5352 6276 5364
rect 6043 5324 6276 5352
rect 6043 5321 6055 5324
rect 5997 5315 6055 5321
rect 6270 5312 6276 5324
rect 6328 5312 6334 5364
rect 6822 5352 6828 5364
rect 6472 5324 6828 5352
rect 3878 5284 3884 5296
rect 1268 5256 1992 5284
rect 2056 5256 3188 5284
rect 3252 5256 3884 5284
rect 1268 5244 1274 5256
rect 842 5176 848 5228
rect 900 5216 906 5228
rect 1581 5219 1639 5225
rect 1581 5216 1593 5219
rect 900 5188 1593 5216
rect 900 5176 906 5188
rect 1581 5185 1593 5188
rect 1627 5185 1639 5219
rect 1581 5179 1639 5185
rect 1857 5219 1915 5225
rect 1857 5185 1869 5219
rect 1903 5185 1915 5219
rect 1964 5216 1992 5256
rect 3252 5225 3280 5256
rect 3878 5244 3884 5256
rect 3936 5244 3942 5296
rect 5169 5287 5227 5293
rect 5169 5253 5181 5287
rect 5215 5284 5227 5287
rect 5350 5284 5356 5296
rect 5215 5256 5356 5284
rect 5215 5253 5227 5256
rect 5169 5247 5227 5253
rect 5350 5244 5356 5256
rect 5408 5244 5414 5296
rect 5920 5284 5948 5312
rect 6472 5293 6500 5324
rect 6822 5312 6828 5324
rect 6880 5312 6886 5364
rect 6917 5355 6975 5361
rect 6917 5321 6929 5355
rect 6963 5352 6975 5355
rect 7006 5352 7012 5364
rect 6963 5324 7012 5352
rect 6963 5321 6975 5324
rect 6917 5315 6975 5321
rect 7006 5312 7012 5324
rect 7064 5312 7070 5364
rect 8938 5352 8944 5364
rect 7116 5324 8944 5352
rect 6457 5287 6515 5293
rect 6457 5284 6469 5287
rect 5920 5256 6469 5284
rect 6457 5253 6469 5256
rect 6503 5253 6515 5287
rect 7116 5284 7144 5324
rect 8938 5312 8944 5324
rect 8996 5312 9002 5364
rect 9674 5312 9680 5364
rect 9732 5352 9738 5364
rect 9732 5324 16160 5352
rect 9732 5312 9738 5324
rect 10686 5284 10692 5296
rect 6457 5247 6515 5253
rect 6564 5256 7144 5284
rect 7392 5256 10180 5284
rect 2225 5219 2283 5225
rect 2225 5216 2237 5219
rect 1964 5188 2237 5216
rect 1857 5179 1915 5185
rect 2225 5185 2237 5188
rect 2271 5185 2283 5219
rect 2225 5179 2283 5185
rect 2593 5219 2651 5225
rect 2593 5185 2605 5219
rect 2639 5185 2651 5219
rect 2593 5179 2651 5185
rect 3237 5219 3295 5225
rect 3237 5185 3249 5219
rect 3283 5185 3295 5219
rect 3237 5179 3295 5185
rect 3329 5219 3387 5225
rect 3329 5185 3341 5219
rect 3375 5216 3387 5219
rect 3510 5216 3516 5228
rect 3375 5188 3516 5216
rect 3375 5185 3387 5188
rect 3329 5179 3387 5185
rect 934 5108 940 5160
rect 992 5148 998 5160
rect 1872 5148 1900 5179
rect 992 5120 1900 5148
rect 992 5108 998 5120
rect 1762 5040 1768 5092
rect 1820 5040 1826 5092
rect 2608 5080 2636 5179
rect 3510 5176 3516 5188
rect 3568 5176 3574 5228
rect 3602 5176 3608 5228
rect 3660 5216 3666 5228
rect 4525 5219 4583 5225
rect 4525 5216 4537 5219
rect 3660 5188 4537 5216
rect 3660 5176 3666 5188
rect 4525 5185 4537 5188
rect 4571 5185 4583 5219
rect 4525 5179 4583 5185
rect 5261 5219 5319 5225
rect 5261 5185 5273 5219
rect 5307 5185 5319 5219
rect 5261 5179 5319 5185
rect 4985 5151 5043 5157
rect 4985 5117 4997 5151
rect 5031 5117 5043 5151
rect 5276 5148 5304 5179
rect 6178 5176 6184 5228
rect 6236 5176 6242 5228
rect 6270 5176 6276 5228
rect 6328 5216 6334 5228
rect 6564 5216 6592 5256
rect 6328 5188 6592 5216
rect 6733 5219 6791 5225
rect 6328 5176 6334 5188
rect 6733 5185 6745 5219
rect 6779 5216 6791 5219
rect 7006 5216 7012 5228
rect 6779 5188 7012 5216
rect 6779 5185 6791 5188
rect 6733 5179 6791 5185
rect 7006 5176 7012 5188
rect 7064 5176 7070 5228
rect 7392 5148 7420 5256
rect 7834 5176 7840 5228
rect 7892 5216 7898 5228
rect 8122 5219 8180 5225
rect 8122 5216 8134 5219
rect 7892 5188 8134 5216
rect 7892 5176 7898 5188
rect 8122 5185 8134 5188
rect 8168 5185 8180 5219
rect 8122 5179 8180 5185
rect 8748 5219 8806 5225
rect 8748 5185 8760 5219
rect 8794 5216 8806 5219
rect 9030 5216 9036 5228
rect 8794 5188 9036 5216
rect 8794 5185 8806 5188
rect 8748 5179 8806 5185
rect 9030 5176 9036 5188
rect 9088 5176 9094 5228
rect 9122 5176 9128 5228
rect 9180 5216 9186 5228
rect 9858 5216 9864 5228
rect 9180 5188 9864 5216
rect 9180 5176 9186 5188
rect 9858 5176 9864 5188
rect 9916 5176 9922 5228
rect 5276 5120 7420 5148
rect 8389 5151 8447 5157
rect 4985 5111 5043 5117
rect 8389 5117 8401 5151
rect 8435 5148 8447 5151
rect 8478 5148 8484 5160
rect 8435 5120 8484 5148
rect 8435 5117 8447 5120
rect 8389 5111 8447 5117
rect 1872 5052 2636 5080
rect 106 4972 112 5024
rect 164 5012 170 5024
rect 1872 5012 1900 5052
rect 2774 5040 2780 5092
rect 2832 5040 2838 5092
rect 4341 5083 4399 5089
rect 4341 5049 4353 5083
rect 4387 5080 4399 5083
rect 5000 5080 5028 5111
rect 8478 5108 8484 5120
rect 8536 5108 8542 5160
rect 10152 5148 10180 5256
rect 10244 5256 10692 5284
rect 10244 5225 10272 5256
rect 10686 5244 10692 5256
rect 10744 5244 10750 5296
rect 11238 5244 11244 5296
rect 11296 5284 11302 5296
rect 13354 5284 13360 5296
rect 11296 5256 11744 5284
rect 11296 5244 11302 5256
rect 10229 5219 10287 5225
rect 10229 5185 10241 5219
rect 10275 5185 10287 5219
rect 10229 5179 10287 5185
rect 10318 5176 10324 5228
rect 10376 5176 10382 5228
rect 10410 5176 10416 5228
rect 10468 5176 10474 5228
rect 10597 5219 10655 5225
rect 10597 5185 10609 5219
rect 10643 5216 10655 5219
rect 11422 5216 11428 5228
rect 10643 5188 11428 5216
rect 10643 5185 10655 5188
rect 10597 5179 10655 5185
rect 11422 5176 11428 5188
rect 11480 5216 11486 5228
rect 11716 5225 11744 5256
rect 11900 5256 13360 5284
rect 11517 5219 11575 5225
rect 11517 5216 11529 5219
rect 11480 5188 11529 5216
rect 11480 5176 11486 5188
rect 11517 5185 11529 5188
rect 11563 5185 11575 5219
rect 11517 5179 11575 5185
rect 11701 5219 11759 5225
rect 11701 5185 11713 5219
rect 11747 5185 11759 5219
rect 11701 5179 11759 5185
rect 11790 5176 11796 5228
rect 11848 5176 11854 5228
rect 11900 5225 11928 5256
rect 13354 5244 13360 5256
rect 13412 5244 13418 5296
rect 14752 5256 15240 5284
rect 14752 5228 14780 5256
rect 11885 5219 11943 5225
rect 11885 5185 11897 5219
rect 11931 5185 11943 5219
rect 11885 5179 11943 5185
rect 11974 5176 11980 5228
rect 12032 5216 12038 5228
rect 12437 5219 12495 5225
rect 12437 5216 12449 5219
rect 12032 5188 12449 5216
rect 12032 5176 12038 5188
rect 12437 5185 12449 5188
rect 12483 5216 12495 5219
rect 14734 5216 14740 5228
rect 12483 5188 14740 5216
rect 12483 5185 12495 5188
rect 12437 5179 12495 5185
rect 14734 5176 14740 5188
rect 14792 5176 14798 5228
rect 15212 5216 15240 5256
rect 15470 5244 15476 5296
rect 15528 5244 15534 5296
rect 15654 5244 15660 5296
rect 15712 5293 15718 5296
rect 15712 5284 15724 5293
rect 15712 5256 15757 5284
rect 15712 5247 15724 5256
rect 15712 5244 15718 5247
rect 15488 5216 15516 5244
rect 15933 5219 15991 5225
rect 15933 5216 15945 5219
rect 15212 5215 15700 5216
rect 15764 5215 15945 5216
rect 15212 5188 15945 5215
rect 15672 5187 15792 5188
rect 15933 5185 15945 5188
rect 15979 5185 15991 5219
rect 15933 5179 15991 5185
rect 16025 5219 16083 5225
rect 16025 5185 16037 5219
rect 16071 5185 16083 5219
rect 16132 5216 16160 5324
rect 16206 5312 16212 5364
rect 16264 5312 16270 5364
rect 18322 5352 18328 5364
rect 18064 5324 18328 5352
rect 17402 5284 17408 5296
rect 16684 5256 17408 5284
rect 16684 5225 16712 5256
rect 17402 5244 17408 5256
rect 17460 5244 17466 5296
rect 17586 5244 17592 5296
rect 17644 5284 17650 5296
rect 18064 5293 18092 5324
rect 18322 5312 18328 5324
rect 18380 5312 18386 5364
rect 18690 5312 18696 5364
rect 18748 5361 18754 5364
rect 18748 5355 18797 5361
rect 18748 5321 18751 5355
rect 18785 5321 18797 5355
rect 18748 5315 18797 5321
rect 18748 5312 18754 5315
rect 19426 5312 19432 5364
rect 19484 5352 19490 5364
rect 19484 5324 21312 5352
rect 19484 5312 19490 5324
rect 18049 5287 18107 5293
rect 18049 5284 18061 5287
rect 17644 5256 18061 5284
rect 17644 5244 17650 5256
rect 18049 5253 18061 5256
rect 18095 5253 18107 5287
rect 18049 5247 18107 5253
rect 18141 5287 18199 5293
rect 18141 5253 18153 5287
rect 18187 5284 18199 5287
rect 21174 5284 21180 5296
rect 18187 5256 21180 5284
rect 18187 5253 18199 5256
rect 18141 5247 18199 5253
rect 21174 5244 21180 5256
rect 21232 5244 21238 5296
rect 16669 5219 16727 5225
rect 16669 5216 16681 5219
rect 16132 5188 16681 5216
rect 16025 5179 16083 5185
rect 16669 5185 16681 5188
rect 16715 5185 16727 5219
rect 16669 5179 16727 5185
rect 11333 5151 11391 5157
rect 10152 5120 11192 5148
rect 4387 5052 5028 5080
rect 4387 5049 4399 5052
rect 4341 5043 4399 5049
rect 5350 5040 5356 5092
rect 5408 5080 5414 5092
rect 6362 5080 6368 5092
rect 5408 5052 6368 5080
rect 5408 5040 5414 5052
rect 6362 5040 6368 5052
rect 6420 5080 6426 5092
rect 6641 5083 6699 5089
rect 6420 5052 6592 5080
rect 6420 5040 6426 5052
rect 164 4984 1900 5012
rect 2317 5015 2375 5021
rect 164 4972 170 4984
rect 2317 4981 2329 5015
rect 2363 5012 2375 5015
rect 3418 5012 3424 5024
rect 2363 4984 3424 5012
rect 2363 4981 2375 4984
rect 2317 4975 2375 4981
rect 3418 4972 3424 4984
rect 3476 4972 3482 5024
rect 4614 4972 4620 5024
rect 4672 4972 4678 5024
rect 5534 4972 5540 5024
rect 5592 5012 5598 5024
rect 5629 5015 5687 5021
rect 5629 5012 5641 5015
rect 5592 4984 5641 5012
rect 5592 4972 5598 4984
rect 5629 4981 5641 4984
rect 5675 4981 5687 5015
rect 5629 4975 5687 4981
rect 5810 4972 5816 5024
rect 5868 5012 5874 5024
rect 6086 5012 6092 5024
rect 5868 4984 6092 5012
rect 5868 4972 5874 4984
rect 6086 4972 6092 4984
rect 6144 4972 6150 5024
rect 6564 5012 6592 5052
rect 6641 5049 6653 5083
rect 6687 5080 6699 5083
rect 6730 5080 6736 5092
rect 6687 5052 6736 5080
rect 6687 5049 6699 5052
rect 6641 5043 6699 5049
rect 6730 5040 6736 5052
rect 6788 5040 6794 5092
rect 10226 5080 10232 5092
rect 9416 5052 10232 5080
rect 7009 5015 7067 5021
rect 7009 5012 7021 5015
rect 6564 4984 7021 5012
rect 7009 4981 7021 4984
rect 7055 4981 7067 5015
rect 7009 4975 7067 4981
rect 7466 4972 7472 5024
rect 7524 5012 7530 5024
rect 9416 5012 9444 5052
rect 10226 5040 10232 5052
rect 10284 5040 10290 5092
rect 7524 4984 9444 5012
rect 7524 4972 7530 4984
rect 9858 4972 9864 5024
rect 9916 4972 9922 5024
rect 9950 4972 9956 5024
rect 10008 4972 10014 5024
rect 10689 5015 10747 5021
rect 10689 4981 10701 5015
rect 10735 5012 10747 5015
rect 11054 5012 11060 5024
rect 10735 4984 11060 5012
rect 10735 4981 10747 4984
rect 10689 4975 10747 4981
rect 11054 4972 11060 4984
rect 11112 4972 11118 5024
rect 11164 5012 11192 5120
rect 11333 5117 11345 5151
rect 11379 5148 11391 5151
rect 12894 5148 12900 5160
rect 11379 5120 12900 5148
rect 11379 5117 11391 5120
rect 11333 5111 11391 5117
rect 12894 5108 12900 5120
rect 12952 5108 12958 5160
rect 14182 5108 14188 5160
rect 14240 5148 14246 5160
rect 14826 5148 14832 5160
rect 14240 5120 14832 5148
rect 14240 5108 14246 5120
rect 14826 5108 14832 5120
rect 14884 5108 14890 5160
rect 12158 5040 12164 5092
rect 12216 5040 12222 5092
rect 12618 5040 12624 5092
rect 12676 5080 12682 5092
rect 12676 5052 14688 5080
rect 12676 5040 12682 5052
rect 14182 5012 14188 5024
rect 11164 4984 14188 5012
rect 14182 4972 14188 4984
rect 14240 4972 14246 5024
rect 14458 4972 14464 5024
rect 14516 5012 14522 5024
rect 14553 5015 14611 5021
rect 14553 5012 14565 5015
rect 14516 4984 14565 5012
rect 14516 4972 14522 4984
rect 14553 4981 14565 4984
rect 14599 4981 14611 5015
rect 14660 5012 14688 5052
rect 16040 5012 16068 5179
rect 16942 5176 16948 5228
rect 17000 5176 17006 5228
rect 17420 5216 17448 5244
rect 18842 5219 18900 5225
rect 17420 5188 18000 5216
rect 17865 5151 17923 5157
rect 17865 5117 17877 5151
rect 17911 5117 17923 5151
rect 17972 5148 18000 5188
rect 18842 5185 18854 5219
rect 18888 5216 18900 5219
rect 18966 5216 18972 5228
rect 18888 5188 18972 5216
rect 18888 5185 18900 5188
rect 18842 5179 18900 5185
rect 18966 5176 18972 5188
rect 19024 5176 19030 5228
rect 19150 5216 19156 5228
rect 19111 5188 19156 5216
rect 19150 5176 19156 5188
rect 19208 5216 19214 5228
rect 19610 5216 19616 5228
rect 19208 5188 19616 5216
rect 19208 5176 19214 5188
rect 19610 5176 19616 5188
rect 19668 5216 19674 5228
rect 19705 5219 19763 5225
rect 19705 5216 19717 5219
rect 19668 5188 19717 5216
rect 19668 5176 19674 5188
rect 19705 5185 19717 5188
rect 19751 5185 19763 5219
rect 19705 5179 19763 5185
rect 20438 5176 20444 5228
rect 20496 5216 20502 5228
rect 20809 5219 20867 5225
rect 20809 5216 20821 5219
rect 20496 5188 20821 5216
rect 20496 5176 20502 5188
rect 20809 5185 20821 5188
rect 20855 5185 20867 5219
rect 20809 5179 20867 5185
rect 19426 5148 19432 5160
rect 17972 5120 19432 5148
rect 17865 5111 17923 5117
rect 17681 5083 17739 5089
rect 17681 5049 17693 5083
rect 17727 5080 17739 5083
rect 17880 5080 17908 5111
rect 19426 5108 19432 5120
rect 19484 5108 19490 5160
rect 20346 5108 20352 5160
rect 20404 5148 20410 5160
rect 20533 5151 20591 5157
rect 20533 5148 20545 5151
rect 20404 5120 20545 5148
rect 20404 5108 20410 5120
rect 20533 5117 20545 5120
rect 20579 5117 20591 5151
rect 21284 5148 21312 5324
rect 21542 5312 21548 5364
rect 21600 5352 21606 5364
rect 21821 5355 21879 5361
rect 21821 5352 21833 5355
rect 21600 5324 21833 5352
rect 21600 5312 21606 5324
rect 21821 5321 21833 5324
rect 21867 5321 21879 5355
rect 21821 5315 21879 5321
rect 23474 5312 23480 5364
rect 23532 5312 23538 5364
rect 25133 5355 25191 5361
rect 25133 5321 25145 5355
rect 25179 5352 25191 5355
rect 25314 5352 25320 5364
rect 25179 5324 25320 5352
rect 25179 5321 25191 5324
rect 25133 5315 25191 5321
rect 25314 5312 25320 5324
rect 25372 5312 25378 5364
rect 26694 5312 26700 5364
rect 26752 5352 26758 5364
rect 26973 5355 27031 5361
rect 26973 5352 26985 5355
rect 26752 5324 26985 5352
rect 26752 5312 26758 5324
rect 26973 5321 26985 5324
rect 27019 5321 27031 5355
rect 26973 5315 27031 5321
rect 27154 5312 27160 5364
rect 27212 5352 27218 5364
rect 27430 5352 27436 5364
rect 27212 5324 27436 5352
rect 27212 5312 27218 5324
rect 27430 5312 27436 5324
rect 27488 5312 27494 5364
rect 29086 5312 29092 5364
rect 29144 5312 29150 5364
rect 29178 5312 29184 5364
rect 29236 5312 29242 5364
rect 29638 5312 29644 5364
rect 29696 5352 29702 5364
rect 29825 5355 29883 5361
rect 29825 5352 29837 5355
rect 29696 5324 29837 5352
rect 29696 5312 29702 5324
rect 29825 5321 29837 5324
rect 29871 5352 29883 5355
rect 30193 5355 30251 5361
rect 30193 5352 30205 5355
rect 29871 5324 30205 5352
rect 29871 5321 29883 5324
rect 29825 5315 29883 5321
rect 30193 5321 30205 5324
rect 30239 5321 30251 5355
rect 30193 5315 30251 5321
rect 30282 5312 30288 5364
rect 30340 5352 30346 5364
rect 31757 5355 31815 5361
rect 31757 5352 31769 5355
rect 30340 5324 31769 5352
rect 30340 5312 30346 5324
rect 31757 5321 31769 5324
rect 31803 5352 31815 5355
rect 32398 5352 32404 5364
rect 31803 5324 32404 5352
rect 31803 5321 31815 5324
rect 31757 5315 31815 5321
rect 32398 5312 32404 5324
rect 32456 5312 32462 5364
rect 36538 5312 36544 5364
rect 36596 5352 36602 5364
rect 37277 5355 37335 5361
rect 37277 5352 37289 5355
rect 36596 5324 37289 5352
rect 36596 5312 36602 5324
rect 37277 5321 37289 5324
rect 37323 5321 37335 5355
rect 37277 5315 37335 5321
rect 38289 5355 38347 5361
rect 38289 5321 38301 5355
rect 38335 5352 38347 5355
rect 38378 5352 38384 5364
rect 38335 5324 38384 5352
rect 38335 5321 38347 5324
rect 38289 5315 38347 5321
rect 38378 5312 38384 5324
rect 38436 5312 38442 5364
rect 38565 5355 38623 5361
rect 38565 5321 38577 5355
rect 38611 5352 38623 5355
rect 38746 5352 38752 5364
rect 38611 5324 38752 5352
rect 38611 5321 38623 5324
rect 38565 5315 38623 5321
rect 38746 5312 38752 5324
rect 38804 5312 38810 5364
rect 39390 5312 39396 5364
rect 39448 5312 39454 5364
rect 21450 5244 21456 5296
rect 21508 5284 21514 5296
rect 21508 5256 22968 5284
rect 21508 5244 21514 5256
rect 22189 5219 22247 5225
rect 22189 5185 22201 5219
rect 22235 5216 22247 5219
rect 22235 5188 22876 5216
rect 22235 5185 22247 5188
rect 22189 5179 22247 5185
rect 22094 5148 22100 5160
rect 21284 5120 22100 5148
rect 20533 5111 20591 5117
rect 19150 5080 19156 5092
rect 17727 5052 17908 5080
rect 18432 5052 19156 5080
rect 17727 5049 17739 5052
rect 17681 5043 17739 5049
rect 14660 4984 16068 5012
rect 14553 4975 14611 4981
rect 16206 4972 16212 5024
rect 16264 5012 16270 5024
rect 18432 5012 18460 5052
rect 19150 5040 19156 5052
rect 19208 5040 19214 5092
rect 19334 5040 19340 5092
rect 19392 5040 19398 5092
rect 21652 5024 21680 5120
rect 22094 5108 22100 5120
rect 22152 5148 22158 5160
rect 22281 5151 22339 5157
rect 22281 5148 22293 5151
rect 22152 5120 22293 5148
rect 22152 5108 22158 5120
rect 22281 5117 22293 5120
rect 22327 5117 22339 5151
rect 22281 5111 22339 5117
rect 22370 5108 22376 5160
rect 22428 5108 22434 5160
rect 22848 5080 22876 5188
rect 22940 5148 22968 5256
rect 23198 5244 23204 5296
rect 23256 5284 23262 5296
rect 25498 5284 25504 5296
rect 23256 5256 25504 5284
rect 23256 5244 23262 5256
rect 25498 5244 25504 5256
rect 25556 5244 25562 5296
rect 26326 5284 26332 5296
rect 25792 5256 26332 5284
rect 23014 5176 23020 5228
rect 23072 5176 23078 5228
rect 23109 5219 23167 5225
rect 23109 5185 23121 5219
rect 23155 5216 23167 5219
rect 23382 5216 23388 5228
rect 23155 5188 23388 5216
rect 23155 5185 23167 5188
rect 23109 5179 23167 5185
rect 23382 5176 23388 5188
rect 23440 5176 23446 5228
rect 23566 5176 23572 5228
rect 23624 5176 23630 5228
rect 23750 5176 23756 5228
rect 23808 5176 23814 5228
rect 25590 5216 25596 5228
rect 24964 5188 25596 5216
rect 24964 5157 24992 5188
rect 25590 5176 25596 5188
rect 25648 5176 25654 5228
rect 25792 5225 25820 5256
rect 26326 5244 26332 5256
rect 26384 5244 26390 5296
rect 26418 5244 26424 5296
rect 26476 5284 26482 5296
rect 26476 5256 27476 5284
rect 26476 5244 26482 5256
rect 25777 5219 25835 5225
rect 25777 5185 25789 5219
rect 25823 5185 25835 5219
rect 25777 5179 25835 5185
rect 25958 5176 25964 5228
rect 26016 5216 26022 5228
rect 26053 5219 26111 5225
rect 26053 5216 26065 5219
rect 26016 5188 26065 5216
rect 26016 5176 26022 5188
rect 26053 5185 26065 5188
rect 26099 5185 26111 5219
rect 26053 5179 26111 5185
rect 27157 5219 27215 5225
rect 27157 5185 27169 5219
rect 27203 5216 27215 5219
rect 27338 5216 27344 5228
rect 27203 5188 27344 5216
rect 27203 5185 27215 5188
rect 27157 5179 27215 5185
rect 27338 5176 27344 5188
rect 27396 5176 27402 5228
rect 27448 5216 27476 5256
rect 29454 5244 29460 5296
rect 29512 5284 29518 5296
rect 29512 5256 31064 5284
rect 29512 5244 29518 5256
rect 27614 5216 27620 5228
rect 27448 5188 27620 5216
rect 27614 5176 27620 5188
rect 27672 5176 27678 5228
rect 28350 5225 28356 5228
rect 28307 5219 28356 5225
rect 28307 5185 28319 5219
rect 28353 5185 28356 5219
rect 28307 5179 28356 5185
rect 28350 5176 28356 5179
rect 28408 5176 28414 5228
rect 30650 5176 30656 5228
rect 30708 5216 30714 5228
rect 30929 5219 30987 5225
rect 30929 5216 30941 5219
rect 30708 5188 30941 5216
rect 30708 5176 30714 5188
rect 30929 5185 30941 5188
rect 30975 5185 30987 5219
rect 31036 5216 31064 5256
rect 32030 5244 32036 5296
rect 32088 5284 32094 5296
rect 32088 5256 32444 5284
rect 32088 5244 32094 5256
rect 32416 5225 32444 5256
rect 31941 5219 31999 5225
rect 31941 5216 31953 5219
rect 31036 5188 31953 5216
rect 30929 5179 30987 5185
rect 31941 5185 31953 5188
rect 31987 5216 31999 5219
rect 32125 5219 32183 5225
rect 32125 5216 32137 5219
rect 31987 5188 32137 5216
rect 31987 5185 31999 5188
rect 31941 5179 31999 5185
rect 32125 5185 32137 5188
rect 32171 5185 32183 5219
rect 32125 5179 32183 5185
rect 32401 5219 32459 5225
rect 32401 5185 32413 5219
rect 32447 5185 32459 5219
rect 32401 5179 32459 5185
rect 37461 5219 37519 5225
rect 37461 5185 37473 5219
rect 37507 5216 37519 5219
rect 37734 5216 37740 5228
rect 37507 5188 37740 5216
rect 37507 5185 37519 5188
rect 37461 5179 37519 5185
rect 37734 5176 37740 5188
rect 37792 5176 37798 5228
rect 38194 5176 38200 5228
rect 38252 5216 38258 5228
rect 38473 5219 38531 5225
rect 38473 5216 38485 5219
rect 38252 5188 38485 5216
rect 38252 5176 38258 5188
rect 38473 5185 38485 5188
rect 38519 5185 38531 5219
rect 38473 5179 38531 5185
rect 38654 5176 38660 5228
rect 38712 5216 38718 5228
rect 38749 5219 38807 5225
rect 38749 5216 38761 5219
rect 38712 5188 38761 5216
rect 38712 5176 38718 5188
rect 38749 5185 38761 5188
rect 38795 5185 38807 5219
rect 38749 5179 38807 5185
rect 38841 5219 38899 5225
rect 38841 5185 38853 5219
rect 38887 5185 38899 5219
rect 38841 5179 38899 5185
rect 39209 5219 39267 5225
rect 39209 5185 39221 5219
rect 39255 5185 39267 5219
rect 39209 5179 39267 5185
rect 23201 5151 23259 5157
rect 23201 5148 23213 5151
rect 22940 5120 23213 5148
rect 23201 5117 23213 5120
rect 23247 5117 23259 5151
rect 23201 5111 23259 5117
rect 23293 5151 23351 5157
rect 23293 5117 23305 5151
rect 23339 5148 23351 5151
rect 23661 5151 23719 5157
rect 23661 5148 23673 5151
rect 23339 5120 23673 5148
rect 23339 5117 23351 5120
rect 23293 5111 23351 5117
rect 23661 5117 23673 5120
rect 23707 5117 23719 5151
rect 23661 5111 23719 5117
rect 24949 5151 25007 5157
rect 24949 5117 24961 5151
rect 24995 5117 25007 5151
rect 24949 5111 25007 5117
rect 25041 5151 25099 5157
rect 25041 5117 25053 5151
rect 25087 5148 25099 5151
rect 25682 5148 25688 5160
rect 25087 5120 25688 5148
rect 25087 5117 25099 5120
rect 25041 5111 25099 5117
rect 25056 5080 25084 5111
rect 25682 5108 25688 5120
rect 25740 5108 25746 5160
rect 26786 5108 26792 5160
rect 26844 5108 26850 5160
rect 27062 5108 27068 5160
rect 27120 5148 27126 5160
rect 27249 5151 27307 5157
rect 27249 5148 27261 5151
rect 27120 5120 27261 5148
rect 27120 5108 27126 5120
rect 27249 5117 27261 5120
rect 27295 5117 27307 5151
rect 27249 5111 27307 5117
rect 27433 5151 27491 5157
rect 27433 5117 27445 5151
rect 27479 5117 27491 5151
rect 27632 5148 27660 5176
rect 28169 5151 28227 5157
rect 28169 5148 28181 5151
rect 27632 5120 28181 5148
rect 27433 5111 27491 5117
rect 28169 5117 28181 5120
rect 28215 5117 28227 5151
rect 28169 5111 28227 5117
rect 22848 5052 25084 5080
rect 26804 5080 26832 5108
rect 27448 5080 27476 5111
rect 28442 5108 28448 5160
rect 28500 5108 28506 5160
rect 29365 5151 29423 5157
rect 29365 5148 29377 5151
rect 28828 5120 29377 5148
rect 26804 5052 27476 5080
rect 27448 5024 27476 5052
rect 27890 5040 27896 5092
rect 27948 5040 27954 5092
rect 16264 4984 18460 5012
rect 18509 5015 18567 5021
rect 16264 4972 16270 4984
rect 18509 4981 18521 5015
rect 18555 5012 18567 5015
rect 19058 5012 19064 5024
rect 18555 4984 19064 5012
rect 18555 4981 18567 4984
rect 18509 4975 18567 4981
rect 19058 4972 19064 4984
rect 19116 4972 19122 5024
rect 20441 5015 20499 5021
rect 20441 4981 20453 5015
rect 20487 5012 20499 5015
rect 21266 5012 21272 5024
rect 20487 4984 21272 5012
rect 20487 4981 20499 4984
rect 20441 4975 20499 4981
rect 21266 4972 21272 4984
rect 21324 4972 21330 5024
rect 21542 4972 21548 5024
rect 21600 4972 21606 5024
rect 21634 4972 21640 5024
rect 21692 4972 21698 5024
rect 21726 4972 21732 5024
rect 21784 5012 21790 5024
rect 22278 5012 22284 5024
rect 21784 4984 22284 5012
rect 21784 4972 21790 4984
rect 22278 4972 22284 4984
rect 22336 4972 22342 5024
rect 23290 4972 23296 5024
rect 23348 5012 23354 5024
rect 25222 5012 25228 5024
rect 23348 4984 25228 5012
rect 23348 4972 23354 4984
rect 25222 4972 25228 4984
rect 25280 4972 25286 5024
rect 25501 5015 25559 5021
rect 25501 4981 25513 5015
rect 25547 5012 25559 5015
rect 26694 5012 26700 5024
rect 25547 4984 26700 5012
rect 25547 4981 25559 4984
rect 25501 4975 25559 4981
rect 26694 4972 26700 4984
rect 26752 4972 26758 5024
rect 26786 4972 26792 5024
rect 26844 4972 26850 5024
rect 27430 4972 27436 5024
rect 27488 4972 27494 5024
rect 27522 4972 27528 5024
rect 27580 5012 27586 5024
rect 28828 5012 28856 5120
rect 29365 5117 29377 5120
rect 29411 5117 29423 5151
rect 29365 5111 29423 5117
rect 29457 5151 29515 5157
rect 29457 5117 29469 5151
rect 29503 5117 29515 5151
rect 29457 5111 29515 5117
rect 28902 5040 28908 5092
rect 28960 5080 28966 5092
rect 29472 5080 29500 5111
rect 31202 5108 31208 5160
rect 31260 5108 31266 5160
rect 33870 5108 33876 5160
rect 33928 5148 33934 5160
rect 38856 5148 38884 5179
rect 33928 5120 38884 5148
rect 33928 5108 33934 5120
rect 39224 5080 39252 5179
rect 28960 5052 29500 5080
rect 31726 5052 31892 5080
rect 28960 5040 28966 5052
rect 27580 4984 28856 5012
rect 27580 4972 27586 4984
rect 29822 4972 29828 5024
rect 29880 5012 29886 5024
rect 31726 5012 31754 5052
rect 29880 4984 31754 5012
rect 31864 5012 31892 5052
rect 33060 5052 39252 5080
rect 33060 5012 33088 5052
rect 31864 4984 33088 5012
rect 33137 5015 33195 5021
rect 29880 4972 29886 4984
rect 33137 4981 33149 5015
rect 33183 5012 33195 5015
rect 33502 5012 33508 5024
rect 33183 4984 33508 5012
rect 33183 4981 33195 4984
rect 33137 4975 33195 4981
rect 33502 4972 33508 4984
rect 33560 4972 33566 5024
rect 38194 4972 38200 5024
rect 38252 5012 38258 5024
rect 38470 5012 38476 5024
rect 38252 4984 38476 5012
rect 38252 4972 38258 4984
rect 38470 4972 38476 4984
rect 38528 4972 38534 5024
rect 39022 4972 39028 5024
rect 39080 4972 39086 5024
rect 1104 4922 39836 4944
rect 1104 4870 1950 4922
rect 2002 4870 2014 4922
rect 2066 4870 2078 4922
rect 2130 4870 2142 4922
rect 2194 4870 2206 4922
rect 2258 4870 7950 4922
rect 8002 4870 8014 4922
rect 8066 4870 8078 4922
rect 8130 4870 8142 4922
rect 8194 4870 8206 4922
rect 8258 4870 13950 4922
rect 14002 4870 14014 4922
rect 14066 4870 14078 4922
rect 14130 4870 14142 4922
rect 14194 4870 14206 4922
rect 14258 4870 19950 4922
rect 20002 4870 20014 4922
rect 20066 4870 20078 4922
rect 20130 4870 20142 4922
rect 20194 4870 20206 4922
rect 20258 4870 25950 4922
rect 26002 4870 26014 4922
rect 26066 4870 26078 4922
rect 26130 4870 26142 4922
rect 26194 4870 26206 4922
rect 26258 4870 31950 4922
rect 32002 4870 32014 4922
rect 32066 4870 32078 4922
rect 32130 4870 32142 4922
rect 32194 4870 32206 4922
rect 32258 4870 37950 4922
rect 38002 4870 38014 4922
rect 38066 4870 38078 4922
rect 38130 4870 38142 4922
rect 38194 4870 38206 4922
rect 38258 4870 39836 4922
rect 1104 4848 39836 4870
rect 1486 4768 1492 4820
rect 1544 4808 1550 4820
rect 1581 4811 1639 4817
rect 1581 4808 1593 4811
rect 1544 4780 1593 4808
rect 1544 4768 1550 4780
rect 1581 4777 1593 4780
rect 1627 4777 1639 4811
rect 1581 4771 1639 4777
rect 2406 4768 2412 4820
rect 2464 4768 2470 4820
rect 3421 4811 3479 4817
rect 3421 4777 3433 4811
rect 3467 4808 3479 4811
rect 4798 4808 4804 4820
rect 3467 4780 4804 4808
rect 3467 4777 3479 4780
rect 3421 4771 3479 4777
rect 4798 4768 4804 4780
rect 4856 4768 4862 4820
rect 5092 4780 6592 4808
rect 1118 4700 1124 4752
rect 1176 4740 1182 4752
rect 3789 4743 3847 4749
rect 1176 4712 2268 4740
rect 1176 4700 1182 4712
rect 750 4632 756 4684
rect 808 4672 814 4684
rect 808 4644 1532 4672
rect 808 4632 814 4644
rect 1504 4613 1532 4644
rect 2240 4613 2268 4712
rect 3789 4709 3801 4743
rect 3835 4709 3847 4743
rect 3789 4703 3847 4709
rect 4709 4743 4767 4749
rect 4709 4709 4721 4743
rect 4755 4740 4767 4743
rect 5092 4740 5120 4780
rect 6454 4740 6460 4752
rect 4755 4712 5120 4740
rect 5920 4712 6460 4740
rect 4755 4709 4767 4712
rect 4709 4703 4767 4709
rect 1489 4607 1547 4613
rect 1489 4573 1501 4607
rect 1535 4573 1547 4607
rect 1489 4567 1547 4573
rect 2225 4607 2283 4613
rect 2225 4573 2237 4607
rect 2271 4573 2283 4607
rect 2225 4567 2283 4573
rect 2501 4607 2559 4613
rect 2501 4573 2513 4607
rect 2547 4604 2559 4607
rect 2590 4604 2596 4616
rect 2547 4576 2596 4604
rect 2547 4573 2559 4576
rect 2501 4567 2559 4573
rect 2590 4564 2596 4576
rect 2648 4564 2654 4616
rect 2866 4564 2872 4616
rect 2924 4564 2930 4616
rect 3237 4607 3295 4613
rect 3237 4573 3249 4607
rect 3283 4604 3295 4607
rect 3804 4604 3832 4703
rect 3878 4632 3884 4684
rect 3936 4672 3942 4684
rect 4341 4675 4399 4681
rect 4341 4672 4353 4675
rect 3936 4644 4353 4672
rect 3936 4632 3942 4644
rect 4341 4641 4353 4644
rect 4387 4641 4399 4675
rect 5604 4675 5662 4681
rect 5604 4672 5616 4675
rect 4341 4635 4399 4641
rect 4908 4644 5616 4672
rect 3283 4576 3832 4604
rect 4157 4607 4215 4613
rect 3283 4573 3295 4576
rect 3237 4567 3295 4573
rect 4157 4573 4169 4607
rect 4203 4604 4215 4607
rect 4617 4607 4675 4613
rect 4617 4604 4629 4607
rect 4203 4576 4629 4604
rect 4203 4573 4215 4576
rect 4157 4567 4215 4573
rect 4617 4573 4629 4576
rect 4663 4573 4675 4607
rect 4617 4567 4675 4573
rect 1857 4539 1915 4545
rect 1857 4536 1869 4539
rect 1504 4508 1869 4536
rect 198 4428 204 4480
rect 256 4468 262 4480
rect 1504 4468 1532 4508
rect 1857 4505 1869 4508
rect 1903 4505 1915 4539
rect 1857 4499 1915 4505
rect 2038 4496 2044 4548
rect 2096 4496 2102 4548
rect 4249 4539 4307 4545
rect 4249 4505 4261 4539
rect 4295 4536 4307 4539
rect 4908 4536 4936 4644
rect 5604 4641 5616 4644
rect 5650 4672 5662 4675
rect 5920 4672 5948 4712
rect 6454 4700 6460 4712
rect 6512 4700 6518 4752
rect 6564 4740 6592 4780
rect 6840 4780 7420 4808
rect 6840 4740 6868 4780
rect 6564 4712 6868 4740
rect 5650 4644 5948 4672
rect 5997 4675 6055 4681
rect 5650 4641 5662 4644
rect 5604 4635 5662 4641
rect 5997 4641 6009 4675
rect 6043 4672 6055 4675
rect 6086 4672 6092 4684
rect 6043 4644 6092 4672
rect 6043 4641 6055 4644
rect 5997 4635 6055 4641
rect 6086 4632 6092 4644
rect 6144 4632 6150 4684
rect 6362 4632 6368 4684
rect 6420 4672 6426 4684
rect 6641 4675 6699 4681
rect 6641 4672 6653 4675
rect 6420 4644 6653 4672
rect 6420 4632 6426 4644
rect 6641 4641 6653 4644
rect 6687 4641 6699 4675
rect 7392 4672 7420 4780
rect 7834 4768 7840 4820
rect 7892 4808 7898 4820
rect 8113 4811 8171 4817
rect 8113 4808 8125 4811
rect 7892 4780 8125 4808
rect 7892 4768 7898 4780
rect 8113 4777 8125 4780
rect 8159 4777 8171 4811
rect 8113 4771 8171 4777
rect 9398 4768 9404 4820
rect 9456 4768 9462 4820
rect 9490 4768 9496 4820
rect 9548 4808 9554 4820
rect 11882 4808 11888 4820
rect 9548 4780 11888 4808
rect 9548 4768 9554 4780
rect 11882 4768 11888 4780
rect 11940 4768 11946 4820
rect 13078 4768 13084 4820
rect 13136 4808 13142 4820
rect 14093 4811 14151 4817
rect 14093 4808 14105 4811
rect 13136 4780 14105 4808
rect 13136 4768 13142 4780
rect 14093 4777 14105 4780
rect 14139 4777 14151 4811
rect 14918 4808 14924 4820
rect 14093 4771 14151 4777
rect 14568 4780 14924 4808
rect 7742 4700 7748 4752
rect 7800 4700 7806 4752
rect 8386 4740 8392 4752
rect 7852 4712 8392 4740
rect 7852 4672 7880 4712
rect 8386 4700 8392 4712
rect 8444 4700 8450 4752
rect 9416 4740 9444 4768
rect 9140 4712 9444 4740
rect 10704 4712 11284 4740
rect 9030 4672 9036 4684
rect 7392 4644 7880 4672
rect 8496 4644 9036 4672
rect 6641 4635 6699 4641
rect 5442 4564 5448 4616
rect 5500 4564 5506 4616
rect 5718 4564 5724 4616
rect 5776 4564 5782 4616
rect 6270 4564 6276 4616
rect 6328 4604 6334 4616
rect 6457 4607 6515 4613
rect 6457 4604 6469 4607
rect 6328 4576 6469 4604
rect 6328 4564 6334 4576
rect 6457 4573 6469 4576
rect 6503 4573 6515 4607
rect 6733 4607 6791 4613
rect 6733 4604 6745 4607
rect 6457 4567 6515 4573
rect 6656 4576 6745 4604
rect 6656 4548 6684 4576
rect 6733 4573 6745 4576
rect 6779 4573 6791 4607
rect 6733 4567 6791 4573
rect 7009 4607 7067 4613
rect 7009 4573 7021 4607
rect 7055 4573 7067 4607
rect 7009 4567 7067 4573
rect 4295 4508 4936 4536
rect 4295 4505 4307 4508
rect 4249 4499 4307 4505
rect 6638 4496 6644 4548
rect 6696 4496 6702 4548
rect 256 4440 1532 4468
rect 256 4428 262 4440
rect 2682 4428 2688 4480
rect 2740 4428 2746 4480
rect 3053 4471 3111 4477
rect 3053 4437 3065 4471
rect 3099 4468 3111 4471
rect 4062 4468 4068 4480
rect 3099 4440 4068 4468
rect 3099 4437 3111 4440
rect 3053 4431 3111 4437
rect 4062 4428 4068 4440
rect 4120 4428 4126 4480
rect 4801 4471 4859 4477
rect 4801 4437 4813 4471
rect 4847 4468 4859 4471
rect 5350 4468 5356 4480
rect 4847 4440 5356 4468
rect 4847 4437 4859 4440
rect 4801 4431 4859 4437
rect 5350 4428 5356 4440
rect 5408 4428 5414 4480
rect 6822 4428 6828 4480
rect 6880 4468 6886 4480
rect 7024 4468 7052 4567
rect 8110 4564 8116 4616
rect 8168 4604 8174 4616
rect 8496 4613 8524 4644
rect 9030 4632 9036 4644
rect 9088 4632 9094 4684
rect 8389 4607 8447 4613
rect 8389 4604 8401 4607
rect 8168 4576 8401 4604
rect 8168 4564 8174 4576
rect 8389 4573 8401 4576
rect 8435 4573 8447 4607
rect 8389 4567 8447 4573
rect 8481 4607 8539 4613
rect 8757 4607 8815 4613
rect 8481 4573 8493 4607
rect 8527 4573 8539 4607
rect 8481 4567 8539 4573
rect 8573 4601 8631 4607
rect 8573 4567 8585 4601
rect 8619 4567 8631 4601
rect 8757 4573 8769 4607
rect 8803 4604 8815 4607
rect 9140 4604 9168 4712
rect 9306 4632 9312 4684
rect 9364 4672 9370 4684
rect 9401 4675 9459 4681
rect 9401 4672 9413 4675
rect 9364 4644 9413 4672
rect 9364 4632 9370 4644
rect 9401 4641 9413 4644
rect 9447 4641 9459 4675
rect 9401 4635 9459 4641
rect 8803 4576 9168 4604
rect 9217 4607 9275 4613
rect 8803 4573 8815 4576
rect 8757 4567 8815 4573
rect 9217 4573 9229 4607
rect 9263 4604 9275 4607
rect 9416 4604 9444 4635
rect 9490 4632 9496 4684
rect 9548 4632 9554 4684
rect 10704 4604 10732 4712
rect 10778 4632 10784 4684
rect 10836 4672 10842 4684
rect 11256 4672 11284 4712
rect 11330 4700 11336 4752
rect 11388 4700 11394 4752
rect 11514 4700 11520 4752
rect 11572 4700 11578 4752
rect 12618 4700 12624 4752
rect 12676 4740 12682 4752
rect 12989 4743 13047 4749
rect 12989 4740 13001 4743
rect 12676 4712 13001 4740
rect 12676 4700 12682 4712
rect 12989 4709 13001 4712
rect 13035 4740 13047 4743
rect 13354 4740 13360 4752
rect 13035 4712 13360 4740
rect 13035 4709 13047 4712
rect 12989 4703 13047 4709
rect 13354 4700 13360 4712
rect 13412 4740 13418 4752
rect 14458 4740 14464 4752
rect 13412 4712 13860 4740
rect 13412 4700 13418 4712
rect 11532 4672 11560 4700
rect 10836 4644 11192 4672
rect 11256 4644 11560 4672
rect 10836 4632 10842 4644
rect 11164 4613 11192 4644
rect 13262 4632 13268 4684
rect 13320 4632 13326 4684
rect 10965 4607 11023 4613
rect 10965 4604 10977 4607
rect 9263 4576 9352 4604
rect 9416 4576 10977 4604
rect 9263 4573 9275 4576
rect 9217 4567 9275 4573
rect 8573 4561 8631 4567
rect 8579 4480 8607 4561
rect 6880 4440 7052 4468
rect 6880 4428 6886 4440
rect 8570 4428 8576 4480
rect 8628 4428 8634 4480
rect 9324 4468 9352 4576
rect 10965 4573 10977 4576
rect 11011 4573 11023 4607
rect 10965 4567 11023 4573
rect 11149 4607 11207 4613
rect 11149 4573 11161 4607
rect 11195 4573 11207 4607
rect 11149 4567 11207 4573
rect 11514 4564 11520 4616
rect 11572 4604 11578 4616
rect 11609 4607 11667 4613
rect 11609 4604 11621 4607
rect 11572 4576 11621 4604
rect 11572 4564 11578 4576
rect 11609 4573 11621 4576
rect 11655 4604 11667 4607
rect 12434 4604 12440 4616
rect 11655 4576 12440 4604
rect 11655 4573 11667 4576
rect 11609 4567 11667 4573
rect 12434 4564 12440 4576
rect 12492 4564 12498 4616
rect 13832 4604 13860 4712
rect 13924 4712 14464 4740
rect 13924 4681 13952 4712
rect 14458 4700 14464 4712
rect 14516 4700 14522 4752
rect 13909 4675 13967 4681
rect 13909 4641 13921 4675
rect 13955 4641 13967 4675
rect 14568 4672 14596 4780
rect 14918 4768 14924 4780
rect 14976 4768 14982 4820
rect 15470 4768 15476 4820
rect 15528 4808 15534 4820
rect 16666 4808 16672 4820
rect 15528 4780 16672 4808
rect 15528 4768 15534 4780
rect 16666 4768 16672 4780
rect 16724 4768 16730 4820
rect 17126 4768 17132 4820
rect 17184 4768 17190 4820
rect 18969 4811 19027 4817
rect 17328 4780 18920 4808
rect 16117 4743 16175 4749
rect 16117 4709 16129 4743
rect 16163 4740 16175 4743
rect 16163 4712 16712 4740
rect 16163 4709 16175 4712
rect 16117 4703 16175 4709
rect 13909 4635 13967 4641
rect 14476 4644 14596 4672
rect 14182 4604 14188 4616
rect 13832 4576 14188 4604
rect 14182 4564 14188 4576
rect 14240 4564 14246 4616
rect 14277 4607 14335 4613
rect 14277 4573 14289 4607
rect 14323 4604 14335 4607
rect 14366 4604 14372 4616
rect 14323 4576 14372 4604
rect 14323 4573 14335 4576
rect 14277 4567 14335 4573
rect 14366 4564 14372 4576
rect 14424 4564 14430 4616
rect 14476 4613 14504 4644
rect 14734 4632 14740 4684
rect 14792 4632 14798 4684
rect 15746 4632 15752 4684
rect 15804 4672 15810 4684
rect 15804 4644 16620 4672
rect 15804 4632 15810 4644
rect 14461 4607 14519 4613
rect 14461 4573 14473 4607
rect 14507 4573 14519 4607
rect 16301 4607 16359 4613
rect 16301 4604 16313 4607
rect 14461 4567 14519 4573
rect 14568 4576 16313 4604
rect 9760 4539 9818 4545
rect 9760 4505 9772 4539
rect 9806 4536 9818 4539
rect 9950 4536 9956 4548
rect 9806 4508 9956 4536
rect 9806 4505 9818 4508
rect 9760 4499 9818 4505
rect 9950 4496 9956 4508
rect 10008 4496 10014 4548
rect 11054 4536 11060 4548
rect 10060 4508 11060 4536
rect 10060 4468 10088 4508
rect 11054 4496 11060 4508
rect 11112 4496 11118 4548
rect 11876 4539 11934 4545
rect 11876 4505 11888 4539
rect 11922 4536 11934 4539
rect 12158 4536 12164 4548
rect 11922 4508 12164 4536
rect 11922 4505 11934 4508
rect 11876 4499 11934 4505
rect 12158 4496 12164 4508
rect 12216 4496 12222 4548
rect 13354 4496 13360 4548
rect 13412 4536 13418 4548
rect 14568 4536 14596 4576
rect 16301 4573 16313 4576
rect 16347 4573 16359 4607
rect 16301 4567 16359 4573
rect 16390 4564 16396 4616
rect 16448 4604 16454 4616
rect 16592 4613 16620 4644
rect 16684 4616 16712 4712
rect 16942 4632 16948 4684
rect 17000 4672 17006 4684
rect 17328 4681 17356 4780
rect 18046 4700 18052 4752
rect 18104 4740 18110 4752
rect 18417 4743 18475 4749
rect 18417 4740 18429 4743
rect 18104 4712 18429 4740
rect 18104 4700 18110 4712
rect 18417 4709 18429 4712
rect 18463 4709 18475 4743
rect 18892 4740 18920 4780
rect 18969 4777 18981 4811
rect 19015 4808 19027 4811
rect 21450 4808 21456 4820
rect 19015 4780 21456 4808
rect 19015 4777 19027 4780
rect 18969 4771 19027 4777
rect 19242 4740 19248 4752
rect 18892 4712 19248 4740
rect 18417 4703 18475 4709
rect 19242 4700 19248 4712
rect 19300 4700 19306 4752
rect 20533 4743 20591 4749
rect 20533 4709 20545 4743
rect 20579 4740 20591 4743
rect 20898 4740 20904 4752
rect 20579 4712 20904 4740
rect 20579 4709 20591 4712
rect 20533 4703 20591 4709
rect 20898 4700 20904 4712
rect 20956 4700 20962 4752
rect 17313 4675 17371 4681
rect 17000 4644 17172 4672
rect 17000 4632 17006 4644
rect 16485 4607 16543 4613
rect 16485 4604 16497 4607
rect 16448 4576 16497 4604
rect 16448 4564 16454 4576
rect 16485 4573 16497 4576
rect 16531 4573 16543 4607
rect 16485 4567 16543 4573
rect 16577 4607 16635 4613
rect 16577 4573 16589 4607
rect 16623 4573 16635 4607
rect 16577 4567 16635 4573
rect 16666 4564 16672 4616
rect 16724 4564 16730 4616
rect 17034 4564 17040 4616
rect 17092 4564 17098 4616
rect 13412 4508 14596 4536
rect 15004 4539 15062 4545
rect 13412 4496 13418 4508
rect 15004 4505 15016 4539
rect 15050 4536 15062 4539
rect 16945 4539 17003 4545
rect 16945 4536 16957 4539
rect 15050 4508 16957 4536
rect 15050 4505 15062 4508
rect 15004 4499 15062 4505
rect 16945 4505 16957 4508
rect 16991 4505 17003 4539
rect 17144 4536 17172 4644
rect 17313 4641 17325 4675
rect 17359 4641 17371 4675
rect 17313 4635 17371 4641
rect 19426 4632 19432 4684
rect 19484 4672 19490 4684
rect 19521 4675 19579 4681
rect 19521 4672 19533 4675
rect 19484 4644 19533 4672
rect 19484 4632 19490 4644
rect 19521 4641 19533 4644
rect 19567 4641 19579 4675
rect 19521 4635 19579 4641
rect 20622 4632 20628 4684
rect 20680 4672 20686 4684
rect 21100 4681 21128 4780
rect 21450 4768 21456 4780
rect 21508 4768 21514 4820
rect 22741 4811 22799 4817
rect 22741 4777 22753 4811
rect 22787 4808 22799 4811
rect 23106 4808 23112 4820
rect 22787 4780 23112 4808
rect 22787 4777 22799 4780
rect 22741 4771 22799 4777
rect 23106 4768 23112 4780
rect 23164 4768 23170 4820
rect 23293 4811 23351 4817
rect 23293 4777 23305 4811
rect 23339 4808 23351 4811
rect 23566 4808 23572 4820
rect 23339 4780 23572 4808
rect 23339 4777 23351 4780
rect 23293 4771 23351 4777
rect 23566 4768 23572 4780
rect 23624 4768 23630 4820
rect 23676 4780 26924 4808
rect 22922 4700 22928 4752
rect 22980 4740 22986 4752
rect 23676 4740 23704 4780
rect 22980 4712 23704 4740
rect 22980 4700 22986 4712
rect 23750 4700 23756 4752
rect 23808 4740 23814 4752
rect 26896 4740 26924 4780
rect 27154 4768 27160 4820
rect 27212 4808 27218 4820
rect 27249 4811 27307 4817
rect 27249 4808 27261 4811
rect 27212 4780 27261 4808
rect 27212 4768 27218 4780
rect 27249 4777 27261 4780
rect 27295 4777 27307 4811
rect 27249 4771 27307 4777
rect 27724 4780 28948 4808
rect 27062 4740 27068 4752
rect 23808 4712 25084 4740
rect 26896 4712 27068 4740
rect 23808 4700 23814 4712
rect 21085 4675 21143 4681
rect 20680 4644 20944 4672
rect 20680 4632 20686 4644
rect 17589 4607 17647 4613
rect 17589 4573 17601 4607
rect 17635 4573 17647 4607
rect 17589 4567 17647 4573
rect 17604 4536 17632 4567
rect 18230 4564 18236 4616
rect 18288 4604 18294 4616
rect 18601 4607 18659 4613
rect 18601 4604 18613 4607
rect 18288 4576 18613 4604
rect 18288 4564 18294 4576
rect 18601 4573 18613 4576
rect 18647 4573 18659 4607
rect 18601 4567 18659 4573
rect 18690 4564 18696 4616
rect 18748 4604 18754 4616
rect 18785 4607 18843 4613
rect 18785 4604 18797 4607
rect 18748 4576 18797 4604
rect 18748 4564 18754 4576
rect 18785 4573 18797 4576
rect 18831 4573 18843 4607
rect 18785 4567 18843 4573
rect 19245 4607 19303 4613
rect 19245 4573 19257 4607
rect 19291 4604 19303 4607
rect 19797 4607 19855 4613
rect 19797 4604 19809 4607
rect 19291 4576 19809 4604
rect 19291 4573 19303 4576
rect 19245 4567 19303 4573
rect 19797 4573 19809 4576
rect 19843 4604 19855 4607
rect 20438 4604 20444 4616
rect 19843 4576 20444 4604
rect 19843 4573 19855 4576
rect 19797 4567 19855 4573
rect 19260 4536 19288 4567
rect 20438 4564 20444 4576
rect 20496 4564 20502 4616
rect 20806 4564 20812 4616
rect 20864 4564 20870 4616
rect 20916 4613 20944 4644
rect 21085 4641 21097 4675
rect 21131 4641 21143 4675
rect 21085 4635 21143 4641
rect 21542 4632 21548 4684
rect 21600 4632 21606 4684
rect 21634 4632 21640 4684
rect 21692 4672 21698 4684
rect 21821 4675 21879 4681
rect 21821 4672 21833 4675
rect 21692 4644 21833 4672
rect 21692 4632 21698 4644
rect 21821 4641 21833 4644
rect 21867 4641 21879 4675
rect 21821 4635 21879 4641
rect 21910 4632 21916 4684
rect 21968 4681 21974 4684
rect 21968 4675 22017 4681
rect 21968 4641 21971 4675
rect 22005 4641 22017 4675
rect 21968 4635 22017 4641
rect 22097 4675 22155 4681
rect 22097 4641 22109 4675
rect 22143 4672 22155 4675
rect 22278 4672 22284 4684
rect 22143 4644 22284 4672
rect 22143 4641 22155 4644
rect 22097 4635 22155 4641
rect 21968 4632 21974 4635
rect 22278 4632 22284 4644
rect 22336 4632 22342 4684
rect 23845 4675 23903 4681
rect 23845 4672 23857 4675
rect 23584 4644 23857 4672
rect 23584 4616 23612 4644
rect 23845 4641 23857 4644
rect 23891 4641 23903 4675
rect 23845 4635 23903 4641
rect 23934 4632 23940 4684
rect 23992 4672 23998 4684
rect 24949 4675 25007 4681
rect 24949 4672 24961 4675
rect 23992 4644 24961 4672
rect 23992 4632 23998 4644
rect 24949 4641 24961 4644
rect 24995 4641 25007 4675
rect 24949 4635 25007 4641
rect 20901 4607 20959 4613
rect 20901 4573 20913 4607
rect 20947 4573 20959 4607
rect 20901 4567 20959 4573
rect 23566 4564 23572 4616
rect 23624 4564 23630 4616
rect 23661 4607 23719 4613
rect 23661 4573 23673 4607
rect 23707 4604 23719 4607
rect 24762 4604 24768 4616
rect 23707 4576 24768 4604
rect 23707 4573 23719 4576
rect 23661 4567 23719 4573
rect 24762 4564 24768 4576
rect 24820 4564 24826 4616
rect 24854 4564 24860 4616
rect 24912 4564 24918 4616
rect 25056 4604 25084 4712
rect 27062 4700 27068 4712
rect 27120 4740 27126 4752
rect 27614 4740 27620 4752
rect 27120 4712 27620 4740
rect 27120 4700 27126 4712
rect 27614 4700 27620 4712
rect 27672 4700 27678 4752
rect 25222 4632 25228 4684
rect 25280 4672 25286 4684
rect 25280 4644 26188 4672
rect 25280 4632 25286 4644
rect 25056 4576 25820 4604
rect 17144 4508 17632 4536
rect 18248 4508 19288 4536
rect 16945 4499 17003 4505
rect 9324 4440 10088 4468
rect 10686 4428 10692 4480
rect 10744 4468 10750 4480
rect 10873 4471 10931 4477
rect 10873 4468 10885 4471
rect 10744 4440 10885 4468
rect 10744 4428 10750 4440
rect 10873 4437 10885 4440
rect 10919 4437 10931 4471
rect 10873 4431 10931 4437
rect 12526 4428 12532 4480
rect 12584 4468 12590 4480
rect 14826 4468 14832 4480
rect 12584 4440 14832 4468
rect 12584 4428 12590 4440
rect 14826 4428 14832 4440
rect 14884 4428 14890 4480
rect 15378 4428 15384 4480
rect 15436 4468 15442 4480
rect 15562 4468 15568 4480
rect 15436 4440 15568 4468
rect 15436 4428 15442 4440
rect 15562 4428 15568 4440
rect 15620 4428 15626 4480
rect 16117 4471 16175 4477
rect 16117 4437 16129 4471
rect 16163 4468 16175 4471
rect 16298 4468 16304 4480
rect 16163 4440 16304 4468
rect 16163 4437 16175 4440
rect 16117 4431 16175 4437
rect 16298 4428 16304 4440
rect 16356 4428 16362 4480
rect 16390 4428 16396 4480
rect 16448 4468 16454 4480
rect 18248 4468 18276 4508
rect 23290 4496 23296 4548
rect 23348 4536 23354 4548
rect 23753 4539 23811 4545
rect 23753 4536 23765 4539
rect 23348 4508 23765 4536
rect 23348 4496 23354 4508
rect 23753 4505 23765 4508
rect 23799 4536 23811 4539
rect 25498 4536 25504 4548
rect 23799 4508 25504 4536
rect 23799 4505 23811 4508
rect 23753 4499 23811 4505
rect 25498 4496 25504 4508
rect 25556 4496 25562 4548
rect 16448 4440 18276 4468
rect 16448 4428 16454 4440
rect 18322 4428 18328 4480
rect 18380 4428 18386 4480
rect 19429 4471 19487 4477
rect 19429 4437 19441 4471
rect 19475 4468 19487 4471
rect 20438 4468 20444 4480
rect 19475 4440 20444 4468
rect 19475 4437 19487 4440
rect 19429 4431 19487 4437
rect 20438 4428 20444 4440
rect 20496 4428 20502 4480
rect 20530 4428 20536 4480
rect 20588 4468 20594 4480
rect 20625 4471 20683 4477
rect 20625 4468 20637 4471
rect 20588 4440 20637 4468
rect 20588 4428 20594 4440
rect 20625 4437 20637 4440
rect 20671 4437 20683 4471
rect 20625 4431 20683 4437
rect 20990 4428 20996 4480
rect 21048 4468 21054 4480
rect 21542 4468 21548 4480
rect 21048 4440 21548 4468
rect 21048 4428 21054 4440
rect 21542 4428 21548 4440
rect 21600 4428 21606 4480
rect 24394 4428 24400 4480
rect 24452 4428 24458 4480
rect 24765 4471 24823 4477
rect 24765 4437 24777 4471
rect 24811 4468 24823 4471
rect 25314 4468 25320 4480
rect 24811 4440 25320 4468
rect 24811 4437 24823 4440
rect 24765 4431 24823 4437
rect 25314 4428 25320 4440
rect 25372 4428 25378 4480
rect 25792 4468 25820 4576
rect 26160 4536 26188 4644
rect 26970 4632 26976 4684
rect 27028 4672 27034 4684
rect 27724 4672 27752 4780
rect 28920 4740 28948 4780
rect 28994 4768 29000 4820
rect 29052 4808 29058 4820
rect 29181 4811 29239 4817
rect 29181 4808 29193 4811
rect 29052 4780 29193 4808
rect 29052 4768 29058 4780
rect 29181 4777 29193 4780
rect 29227 4777 29239 4811
rect 30650 4808 30656 4820
rect 29181 4771 29239 4777
rect 29656 4780 30656 4808
rect 29656 4740 29684 4780
rect 30650 4768 30656 4780
rect 30708 4768 30714 4820
rect 34701 4811 34759 4817
rect 34701 4808 34713 4811
rect 31726 4780 34713 4808
rect 28920 4712 29684 4740
rect 29733 4743 29791 4749
rect 29733 4709 29745 4743
rect 29779 4709 29791 4743
rect 31726 4740 31754 4780
rect 34701 4777 34713 4780
rect 34747 4777 34759 4811
rect 34701 4771 34759 4777
rect 35084 4780 35940 4808
rect 29733 4703 29791 4709
rect 31588 4712 31754 4740
rect 31941 4743 31999 4749
rect 27028 4644 27752 4672
rect 27985 4675 28043 4681
rect 27028 4632 27034 4644
rect 27985 4641 27997 4675
rect 28031 4672 28043 4675
rect 28902 4672 28908 4684
rect 28031 4644 28908 4672
rect 28031 4641 28043 4644
rect 27985 4635 28043 4641
rect 28902 4632 28908 4644
rect 28960 4672 28966 4684
rect 29748 4672 29776 4703
rect 28960 4644 29776 4672
rect 28960 4632 28966 4644
rect 26234 4564 26240 4616
rect 26292 4564 26298 4616
rect 26513 4607 26571 4613
rect 26513 4573 26525 4607
rect 26559 4573 26571 4607
rect 26513 4567 26571 4573
rect 26528 4536 26556 4567
rect 26602 4564 26608 4616
rect 26660 4604 26666 4616
rect 27341 4607 27399 4613
rect 27341 4604 27353 4607
rect 26660 4576 27353 4604
rect 26660 4564 26666 4576
rect 27341 4573 27353 4576
rect 27387 4573 27399 4607
rect 27341 4567 27399 4573
rect 27430 4564 27436 4616
rect 27488 4604 27494 4616
rect 27525 4607 27583 4613
rect 27525 4604 27537 4607
rect 27488 4576 27537 4604
rect 27488 4564 27494 4576
rect 27525 4573 27537 4576
rect 27571 4573 27583 4607
rect 27525 4567 27583 4573
rect 28258 4564 28264 4616
rect 28316 4564 28322 4616
rect 28350 4564 28356 4616
rect 28408 4613 28414 4616
rect 28408 4607 28436 4613
rect 28424 4573 28436 4607
rect 28408 4567 28436 4573
rect 28408 4564 28414 4567
rect 28534 4564 28540 4616
rect 28592 4564 28598 4616
rect 30374 4564 30380 4616
rect 30432 4604 30438 4616
rect 30469 4607 30527 4613
rect 30469 4604 30481 4607
rect 30432 4576 30481 4604
rect 30432 4564 30438 4576
rect 30469 4573 30481 4576
rect 30515 4573 30527 4607
rect 30745 4607 30803 4613
rect 30745 4604 30757 4607
rect 30469 4567 30527 4573
rect 30576 4576 30757 4604
rect 26970 4536 26976 4548
rect 26160 4508 26976 4536
rect 26970 4496 26976 4508
rect 27028 4496 27034 4548
rect 29730 4496 29736 4548
rect 29788 4536 29794 4548
rect 30576 4536 30604 4576
rect 30745 4573 30757 4576
rect 30791 4573 30803 4607
rect 30745 4567 30803 4573
rect 30929 4607 30987 4613
rect 30929 4573 30941 4607
rect 30975 4604 30987 4607
rect 31110 4604 31116 4616
rect 30975 4576 31116 4604
rect 30975 4573 30987 4576
rect 30929 4567 30987 4573
rect 31110 4564 31116 4576
rect 31168 4564 31174 4616
rect 31205 4607 31263 4613
rect 31205 4573 31217 4607
rect 31251 4573 31263 4607
rect 31205 4567 31263 4573
rect 29788 4508 30604 4536
rect 29788 4496 29794 4508
rect 30650 4496 30656 4548
rect 30708 4536 30714 4548
rect 31220 4536 31248 4567
rect 30708 4508 31248 4536
rect 30708 4496 30714 4508
rect 31588 4468 31616 4712
rect 31941 4709 31953 4743
rect 31987 4740 31999 4743
rect 31987 4712 32720 4740
rect 31987 4709 31999 4712
rect 31941 4703 31999 4709
rect 31662 4632 31668 4684
rect 31720 4672 31726 4684
rect 32692 4681 32720 4712
rect 33594 4700 33600 4752
rect 33652 4740 33658 4752
rect 35084 4740 35112 4780
rect 33652 4712 35112 4740
rect 35912 4740 35940 4780
rect 35986 4768 35992 4820
rect 36044 4768 36050 4820
rect 36998 4768 37004 4820
rect 37056 4808 37062 4820
rect 37369 4811 37427 4817
rect 37369 4808 37381 4811
rect 37056 4780 37381 4808
rect 37056 4768 37062 4780
rect 37369 4777 37381 4780
rect 37415 4777 37427 4811
rect 37369 4771 37427 4777
rect 37642 4768 37648 4820
rect 37700 4808 37706 4820
rect 38381 4811 38439 4817
rect 38381 4808 38393 4811
rect 37700 4780 38393 4808
rect 37700 4768 37706 4780
rect 38381 4777 38393 4780
rect 38427 4777 38439 4811
rect 38381 4771 38439 4777
rect 38197 4743 38255 4749
rect 38197 4740 38209 4743
rect 35912 4712 38209 4740
rect 33652 4700 33658 4712
rect 38197 4709 38209 4712
rect 38243 4709 38255 4743
rect 38197 4703 38255 4709
rect 39390 4700 39396 4752
rect 39448 4700 39454 4752
rect 32585 4675 32643 4681
rect 32585 4672 32597 4675
rect 31720 4644 32597 4672
rect 31720 4632 31726 4644
rect 32585 4641 32597 4644
rect 32631 4641 32643 4675
rect 32585 4635 32643 4641
rect 32677 4675 32735 4681
rect 32677 4641 32689 4675
rect 32723 4641 32735 4675
rect 32677 4635 32735 4641
rect 32214 4564 32220 4616
rect 32272 4604 32278 4616
rect 32398 4604 32404 4616
rect 32272 4576 32404 4604
rect 32272 4564 32278 4576
rect 32398 4564 32404 4576
rect 32456 4564 32462 4616
rect 32490 4564 32496 4616
rect 32548 4564 32554 4616
rect 32600 4604 32628 4635
rect 33502 4632 33508 4684
rect 33560 4632 33566 4684
rect 38289 4675 38347 4681
rect 38289 4641 38301 4675
rect 38335 4672 38347 4675
rect 38335 4644 38700 4672
rect 38335 4641 38347 4644
rect 38289 4635 38347 4641
rect 33413 4607 33471 4613
rect 33413 4604 33425 4607
rect 32600 4576 33425 4604
rect 33413 4573 33425 4576
rect 33459 4573 33471 4607
rect 33413 4567 33471 4573
rect 35434 4564 35440 4616
rect 35492 4564 35498 4616
rect 35526 4564 35532 4616
rect 35584 4604 35590 4616
rect 38672 4613 38700 4644
rect 35713 4607 35771 4613
rect 35713 4604 35725 4607
rect 35584 4576 35725 4604
rect 35584 4564 35590 4576
rect 35713 4573 35725 4576
rect 35759 4573 35771 4607
rect 35713 4567 35771 4573
rect 35805 4607 35863 4613
rect 35805 4573 35817 4607
rect 35851 4573 35863 4607
rect 37553 4607 37611 4613
rect 37553 4604 37565 4607
rect 35805 4567 35863 4573
rect 35912 4576 37565 4604
rect 32582 4496 32588 4548
rect 32640 4536 32646 4548
rect 33321 4539 33379 4545
rect 33321 4536 33333 4539
rect 32640 4508 33333 4536
rect 32640 4496 32646 4508
rect 33321 4505 33333 4508
rect 33367 4505 33379 4539
rect 35452 4536 35480 4564
rect 35820 4536 35848 4567
rect 35452 4508 35848 4536
rect 33321 4499 33379 4505
rect 25792 4440 31616 4468
rect 32125 4471 32183 4477
rect 32125 4437 32137 4471
rect 32171 4468 32183 4471
rect 32398 4468 32404 4480
rect 32171 4440 32404 4468
rect 32171 4437 32183 4440
rect 32125 4431 32183 4437
rect 32398 4428 32404 4440
rect 32456 4428 32462 4480
rect 32858 4428 32864 4480
rect 32916 4468 32922 4480
rect 32953 4471 33011 4477
rect 32953 4468 32965 4471
rect 32916 4440 32965 4468
rect 32916 4428 32922 4440
rect 32953 4437 32965 4440
rect 32999 4437 33011 4471
rect 32953 4431 33011 4437
rect 35342 4428 35348 4480
rect 35400 4468 35406 4480
rect 35912 4468 35940 4576
rect 37553 4573 37565 4576
rect 37599 4573 37611 4607
rect 37553 4567 37611 4573
rect 38565 4607 38623 4613
rect 38565 4573 38577 4607
rect 38611 4573 38623 4607
rect 38565 4567 38623 4573
rect 38657 4607 38715 4613
rect 38657 4573 38669 4607
rect 38703 4573 38715 4607
rect 38657 4567 38715 4573
rect 39117 4607 39175 4613
rect 39117 4573 39129 4607
rect 39163 4604 39175 4607
rect 39209 4607 39267 4613
rect 39209 4604 39221 4607
rect 39163 4576 39221 4604
rect 39163 4573 39175 4576
rect 39117 4567 39175 4573
rect 39209 4573 39221 4576
rect 39255 4573 39267 4607
rect 39209 4567 39267 4573
rect 36446 4496 36452 4548
rect 36504 4536 36510 4548
rect 38580 4536 38608 4567
rect 39850 4536 39856 4548
rect 36504 4508 38608 4536
rect 38856 4508 39856 4536
rect 36504 4496 36510 4508
rect 38856 4477 38884 4508
rect 39850 4496 39856 4508
rect 39908 4496 39914 4548
rect 35400 4440 35940 4468
rect 38841 4471 38899 4477
rect 35400 4428 35406 4440
rect 38841 4437 38853 4471
rect 38887 4437 38899 4471
rect 38841 4431 38899 4437
rect 39117 4471 39175 4477
rect 39117 4437 39129 4471
rect 39163 4468 39175 4471
rect 39666 4468 39672 4480
rect 39163 4440 39672 4468
rect 39163 4437 39175 4440
rect 39117 4431 39175 4437
rect 39666 4428 39672 4440
rect 39724 4428 39730 4480
rect 1104 4378 39836 4400
rect 1104 4326 3010 4378
rect 3062 4326 3074 4378
rect 3126 4326 3138 4378
rect 3190 4326 3202 4378
rect 3254 4326 3266 4378
rect 3318 4326 9010 4378
rect 9062 4326 9074 4378
rect 9126 4326 9138 4378
rect 9190 4326 9202 4378
rect 9254 4326 9266 4378
rect 9318 4326 15010 4378
rect 15062 4326 15074 4378
rect 15126 4326 15138 4378
rect 15190 4326 15202 4378
rect 15254 4326 15266 4378
rect 15318 4326 21010 4378
rect 21062 4326 21074 4378
rect 21126 4326 21138 4378
rect 21190 4326 21202 4378
rect 21254 4326 21266 4378
rect 21318 4326 27010 4378
rect 27062 4326 27074 4378
rect 27126 4326 27138 4378
rect 27190 4326 27202 4378
rect 27254 4326 27266 4378
rect 27318 4326 33010 4378
rect 33062 4326 33074 4378
rect 33126 4326 33138 4378
rect 33190 4326 33202 4378
rect 33254 4326 33266 4378
rect 33318 4326 39010 4378
rect 39062 4326 39074 4378
rect 39126 4326 39138 4378
rect 39190 4326 39202 4378
rect 39254 4326 39266 4378
rect 39318 4326 39836 4378
rect 1104 4304 39836 4326
rect 3789 4267 3847 4273
rect 2746 4236 3004 4264
rect 2746 4208 2774 4236
rect 2682 4156 2688 4208
rect 2740 4168 2774 4208
rect 2740 4156 2746 4168
rect 2866 4156 2872 4208
rect 2924 4156 2930 4208
rect 2976 4196 3004 4236
rect 3789 4233 3801 4267
rect 3835 4264 3847 4267
rect 3878 4264 3884 4276
rect 3835 4236 3884 4264
rect 3835 4233 3847 4236
rect 3789 4227 3847 4233
rect 3878 4224 3884 4236
rect 3936 4224 3942 4276
rect 4338 4224 4344 4276
rect 4396 4264 4402 4276
rect 5537 4267 5595 4273
rect 5537 4264 5549 4267
rect 4396 4236 5549 4264
rect 4396 4224 4402 4236
rect 5537 4233 5549 4236
rect 5583 4233 5595 4267
rect 5537 4227 5595 4233
rect 6362 4224 6368 4276
rect 6420 4264 6426 4276
rect 6641 4267 6699 4273
rect 6641 4264 6653 4267
rect 6420 4236 6653 4264
rect 6420 4224 6426 4236
rect 6641 4233 6653 4236
rect 6687 4233 6699 4267
rect 6641 4227 6699 4233
rect 6733 4267 6791 4273
rect 6733 4233 6745 4267
rect 6779 4264 6791 4267
rect 6914 4264 6920 4276
rect 6779 4236 6920 4264
rect 6779 4233 6791 4236
rect 6733 4227 6791 4233
rect 6914 4224 6920 4236
rect 6972 4224 6978 4276
rect 7006 4224 7012 4276
rect 7064 4264 7070 4276
rect 7101 4267 7159 4273
rect 7101 4264 7113 4267
rect 7064 4236 7113 4264
rect 7064 4224 7070 4236
rect 7101 4233 7113 4236
rect 7147 4233 7159 4267
rect 7101 4227 7159 4233
rect 8570 4224 8576 4276
rect 8628 4264 8634 4276
rect 8849 4267 8907 4273
rect 8849 4264 8861 4267
rect 8628 4236 8861 4264
rect 8628 4224 8634 4236
rect 8849 4233 8861 4236
rect 8895 4233 8907 4267
rect 9401 4267 9459 4273
rect 8849 4227 8907 4233
rect 9048 4236 9352 4264
rect 7466 4196 7472 4208
rect 2976 4168 7472 4196
rect 7466 4156 7472 4168
rect 7524 4156 7530 4208
rect 8294 4156 8300 4208
rect 8352 4196 8358 4208
rect 9048 4196 9076 4236
rect 8352 4168 8596 4196
rect 8352 4156 8358 4168
rect 8568 4158 8596 4168
rect 8772 4168 9076 4196
rect 290 4088 296 4140
rect 348 4128 354 4140
rect 2501 4131 2559 4137
rect 2501 4128 2513 4131
rect 348 4100 2513 4128
rect 348 4088 354 4100
rect 2501 4097 2513 4100
rect 2547 4097 2559 4131
rect 2884 4128 2912 4156
rect 3053 4131 3111 4137
rect 3053 4128 3065 4131
rect 2884 4100 3065 4128
rect 2501 4091 2559 4097
rect 3053 4097 3065 4100
rect 3099 4128 3111 4131
rect 4157 4131 4215 4137
rect 4157 4128 4169 4131
rect 3099 4100 4169 4128
rect 3099 4097 3111 4100
rect 3053 4091 3111 4097
rect 4157 4097 4169 4100
rect 4203 4097 4215 4131
rect 4157 4091 4215 4097
rect 5166 4088 5172 4140
rect 5224 4088 5230 4140
rect 5258 4088 5264 4140
rect 5316 4088 5322 4140
rect 5350 4088 5356 4140
rect 5408 4128 5414 4140
rect 5721 4131 5779 4137
rect 5721 4128 5733 4131
rect 5408 4100 5733 4128
rect 5408 4088 5414 4100
rect 5721 4097 5733 4100
rect 5767 4097 5779 4131
rect 5721 4091 5779 4097
rect 5810 4088 5816 4140
rect 5868 4088 5874 4140
rect 6641 4131 6699 4137
rect 6641 4097 6653 4131
rect 6687 4128 6699 4131
rect 7006 4128 7012 4140
rect 6687 4100 7012 4128
rect 6687 4097 6699 4100
rect 6641 4091 6699 4097
rect 7006 4088 7012 4100
rect 7064 4128 7070 4140
rect 8110 4128 8116 4140
rect 7064 4100 8116 4128
rect 7064 4088 7070 4100
rect 8110 4088 8116 4100
rect 8168 4088 8174 4140
rect 8205 4131 8263 4137
rect 8205 4097 8217 4131
rect 8251 4097 8263 4131
rect 8205 4091 8263 4097
rect 8481 4131 8539 4137
rect 8481 4097 8493 4131
rect 8527 4097 8539 4131
rect 8568 4130 8616 4158
rect 8772 4137 8800 4168
rect 8588 4128 8616 4130
rect 8665 4131 8723 4137
rect 8665 4128 8677 4131
rect 8588 4100 8677 4128
rect 8481 4091 8539 4097
rect 8665 4097 8677 4100
rect 8711 4097 8723 4131
rect 8665 4091 8723 4097
rect 8757 4131 8815 4137
rect 8938 4135 8944 4138
rect 8757 4097 8769 4131
rect 8803 4097 8815 4131
rect 8932 4126 8944 4135
rect 8899 4098 8944 4126
rect 8757 4091 8815 4097
rect 750 4020 756 4072
rect 808 4060 814 4072
rect 1397 4063 1455 4069
rect 1397 4060 1409 4063
rect 808 4032 1409 4060
rect 808 4020 814 4032
rect 1397 4029 1409 4032
rect 1443 4029 1455 4063
rect 1397 4023 1455 4029
rect 1673 4063 1731 4069
rect 1673 4029 1685 4063
rect 1719 4029 1731 4063
rect 1673 4023 1731 4029
rect 1688 3992 1716 4023
rect 2682 4020 2688 4072
rect 2740 4060 2746 4072
rect 2777 4063 2835 4069
rect 2777 4060 2789 4063
rect 2740 4032 2789 4060
rect 2740 4020 2746 4032
rect 2777 4029 2789 4032
rect 2823 4029 2835 4063
rect 2777 4023 2835 4029
rect 3786 4020 3792 4072
rect 3844 4060 3850 4072
rect 3881 4063 3939 4069
rect 3881 4060 3893 4063
rect 3844 4032 3893 4060
rect 3844 4020 3850 4032
rect 3881 4029 3893 4032
rect 3927 4029 3939 4063
rect 6086 4060 6092 4072
rect 3881 4023 3939 4029
rect 4908 4032 6092 4060
rect 4908 4001 4936 4032
rect 6086 4020 6092 4032
rect 6144 4020 6150 4072
rect 6546 4020 6552 4072
rect 6604 4020 6610 4072
rect 8220 4060 8248 4091
rect 8386 4060 8392 4072
rect 8220 4032 8392 4060
rect 8386 4020 8392 4032
rect 8444 4020 8450 4072
rect 8505 4060 8533 4091
rect 8772 4060 8800 4091
rect 8932 4089 8944 4098
rect 8938 4086 8944 4089
rect 8996 4086 9002 4138
rect 9048 4137 9076 4168
rect 9324 4196 9352 4236
rect 9401 4233 9413 4267
rect 9447 4264 9459 4267
rect 9950 4264 9956 4276
rect 9447 4236 9956 4264
rect 9447 4233 9459 4236
rect 9401 4227 9459 4233
rect 9950 4224 9956 4236
rect 10008 4224 10014 4276
rect 10042 4224 10048 4276
rect 10100 4264 10106 4276
rect 10410 4264 10416 4276
rect 10100 4236 10416 4264
rect 10100 4224 10106 4236
rect 10410 4224 10416 4236
rect 10468 4224 10474 4276
rect 10873 4267 10931 4273
rect 10873 4233 10885 4267
rect 10919 4264 10931 4267
rect 12618 4264 12624 4276
rect 10919 4236 12624 4264
rect 10919 4233 10931 4236
rect 10873 4227 10931 4233
rect 12618 4224 12624 4236
rect 12676 4224 12682 4276
rect 12894 4224 12900 4276
rect 12952 4224 12958 4276
rect 13265 4267 13323 4273
rect 13265 4233 13277 4267
rect 13311 4264 13323 4267
rect 13354 4264 13360 4276
rect 13311 4236 13360 4264
rect 13311 4233 13323 4236
rect 13265 4227 13323 4233
rect 13354 4224 13360 4236
rect 13412 4224 13418 4276
rect 13446 4224 13452 4276
rect 13504 4224 13510 4276
rect 14001 4267 14059 4273
rect 14001 4233 14013 4267
rect 14047 4264 14059 4267
rect 14642 4264 14648 4276
rect 14047 4236 14648 4264
rect 14047 4233 14059 4236
rect 14001 4227 14059 4233
rect 14642 4224 14648 4236
rect 14700 4224 14706 4276
rect 15378 4224 15384 4276
rect 15436 4264 15442 4276
rect 15565 4267 15623 4273
rect 15565 4264 15577 4267
rect 15436 4236 15577 4264
rect 15436 4224 15442 4236
rect 15565 4233 15577 4236
rect 15611 4233 15623 4267
rect 15565 4227 15623 4233
rect 15657 4267 15715 4273
rect 15657 4233 15669 4267
rect 15703 4233 15715 4267
rect 15657 4227 15715 4233
rect 9766 4196 9772 4208
rect 9324 4168 9772 4196
rect 9033 4131 9091 4137
rect 9033 4097 9045 4131
rect 9079 4097 9091 4131
rect 9033 4091 9091 4097
rect 9214 4088 9220 4140
rect 9272 4088 9278 4140
rect 9324 4137 9352 4168
rect 9766 4156 9772 4168
rect 9824 4196 9830 4208
rect 9824 4168 10732 4196
rect 9824 4156 9830 4168
rect 9309 4131 9367 4137
rect 9309 4097 9321 4131
rect 9355 4097 9367 4131
rect 9309 4091 9367 4097
rect 9490 4088 9496 4140
rect 9548 4088 9554 4140
rect 10042 4128 10048 4140
rect 9646 4100 10048 4128
rect 9646 4060 9674 4100
rect 10042 4088 10048 4100
rect 10100 4088 10106 4140
rect 10336 4137 10364 4168
rect 10321 4131 10379 4137
rect 10321 4097 10333 4131
rect 10367 4097 10379 4131
rect 10321 4091 10379 4097
rect 10505 4131 10563 4137
rect 10505 4097 10517 4131
rect 10551 4128 10563 4131
rect 10594 4128 10600 4140
rect 10551 4100 10600 4128
rect 10551 4097 10563 4100
rect 10505 4091 10563 4097
rect 10594 4088 10600 4100
rect 10652 4088 10658 4140
rect 10704 4128 10732 4168
rect 10778 4156 10784 4208
rect 10836 4196 10842 4208
rect 10965 4199 11023 4205
rect 10965 4196 10977 4199
rect 10836 4168 10977 4196
rect 10836 4156 10842 4168
rect 10965 4165 10977 4168
rect 11011 4165 11023 4199
rect 10965 4159 11023 4165
rect 11330 4156 11336 4208
rect 11388 4196 11394 4208
rect 11762 4199 11820 4205
rect 11762 4196 11774 4199
rect 11388 4168 11774 4196
rect 11388 4156 11394 4168
rect 11762 4165 11774 4168
rect 11808 4165 11820 4199
rect 12912 4196 12940 4224
rect 13909 4199 13967 4205
rect 12912 4168 13676 4196
rect 11762 4159 11820 4165
rect 11422 4128 11428 4140
rect 10704 4100 11428 4128
rect 11422 4088 11428 4100
rect 11480 4088 11486 4140
rect 11514 4088 11520 4140
rect 11572 4088 11578 4140
rect 11624 4100 12572 4128
rect 8505 4032 8800 4060
rect 9140 4032 9674 4060
rect 4893 3995 4951 4001
rect 1688 3964 2912 3992
rect 566 3884 572 3936
rect 624 3924 630 3936
rect 2314 3924 2320 3936
rect 624 3896 2320 3924
rect 624 3884 630 3896
rect 2314 3884 2320 3896
rect 2372 3884 2378 3936
rect 2498 3884 2504 3936
rect 2556 3924 2562 3936
rect 2685 3927 2743 3933
rect 2685 3924 2697 3927
rect 2556 3896 2697 3924
rect 2556 3884 2562 3896
rect 2685 3893 2697 3896
rect 2731 3893 2743 3927
rect 2884 3924 2912 3964
rect 4893 3961 4905 3995
rect 4939 3961 4951 3995
rect 4893 3955 4951 3961
rect 4982 3952 4988 4004
rect 5040 3952 5046 4004
rect 5092 3964 5856 3992
rect 5092 3924 5120 3964
rect 2884 3896 5120 3924
rect 2685 3887 2743 3893
rect 5166 3884 5172 3936
rect 5224 3924 5230 3936
rect 5445 3927 5503 3933
rect 5445 3924 5457 3927
rect 5224 3896 5457 3924
rect 5224 3884 5230 3896
rect 5445 3893 5457 3896
rect 5491 3893 5503 3927
rect 5828 3924 5856 3964
rect 5902 3952 5908 4004
rect 5960 3992 5966 4004
rect 5997 3995 6055 4001
rect 5997 3992 6009 3995
rect 5960 3964 6009 3992
rect 5960 3952 5966 3964
rect 5997 3961 6009 3964
rect 6043 3961 6055 3995
rect 5997 3955 6055 3961
rect 7650 3952 7656 4004
rect 7708 3992 7714 4004
rect 8021 3995 8079 4001
rect 8021 3992 8033 3995
rect 7708 3964 8033 3992
rect 7708 3952 7714 3964
rect 8021 3961 8033 3964
rect 8067 3961 8079 3995
rect 8021 3955 8079 3961
rect 8570 3952 8576 4004
rect 8628 3952 8634 4004
rect 9030 3992 9036 4004
rect 8671 3964 9036 3992
rect 8671 3924 8699 3964
rect 9030 3952 9036 3964
rect 9088 3952 9094 4004
rect 9140 4001 9168 4032
rect 9858 4020 9864 4072
rect 9916 4060 9922 4072
rect 10229 4063 10287 4069
rect 10229 4060 10241 4063
rect 9916 4032 10241 4060
rect 9916 4020 9922 4032
rect 10229 4029 10241 4032
rect 10275 4029 10287 4063
rect 10229 4023 10287 4029
rect 9125 3995 9183 4001
rect 9125 3961 9137 3995
rect 9171 3961 9183 3995
rect 9125 3955 9183 3961
rect 9214 3952 9220 4004
rect 9272 3992 9278 4004
rect 9766 3992 9772 4004
rect 9272 3964 9772 3992
rect 9272 3952 9278 3964
rect 9766 3952 9772 3964
rect 9824 3952 9830 4004
rect 10244 3992 10272 4023
rect 10778 4020 10784 4072
rect 10836 4020 10842 4072
rect 11624 4060 11652 4100
rect 10888 4032 11652 4060
rect 10888 3992 10916 4032
rect 10244 3964 10916 3992
rect 12544 3992 12572 4100
rect 13078 4088 13084 4140
rect 13136 4088 13142 4140
rect 13262 4088 13268 4140
rect 13320 4088 13326 4140
rect 13538 4088 13544 4140
rect 13596 4088 13602 4140
rect 13648 4128 13676 4168
rect 13909 4165 13921 4199
rect 13955 4196 13967 4199
rect 14366 4196 14372 4208
rect 13955 4168 14372 4196
rect 13955 4165 13967 4168
rect 13909 4159 13967 4165
rect 14366 4156 14372 4168
rect 14424 4156 14430 4208
rect 14458 4156 14464 4208
rect 14516 4156 14522 4208
rect 14826 4156 14832 4208
rect 14884 4196 14890 4208
rect 15672 4196 15700 4227
rect 15746 4224 15752 4276
rect 15804 4264 15810 4276
rect 16390 4264 16396 4276
rect 15804 4236 16396 4264
rect 15804 4224 15810 4236
rect 16390 4224 16396 4236
rect 16448 4224 16454 4276
rect 16666 4224 16672 4276
rect 16724 4264 16730 4276
rect 18230 4264 18236 4276
rect 16724 4236 18236 4264
rect 16724 4224 16730 4236
rect 18230 4224 18236 4236
rect 18288 4224 18294 4276
rect 18877 4267 18935 4273
rect 18877 4233 18889 4267
rect 18923 4264 18935 4267
rect 22186 4264 22192 4276
rect 18923 4236 22192 4264
rect 18923 4233 18935 4236
rect 18877 4227 18935 4233
rect 22186 4224 22192 4236
rect 22244 4224 22250 4276
rect 22281 4267 22339 4273
rect 22281 4233 22293 4267
rect 22327 4264 22339 4267
rect 23106 4264 23112 4276
rect 22327 4236 23112 4264
rect 22327 4233 22339 4236
rect 22281 4227 22339 4233
rect 16758 4196 16764 4208
rect 14884 4168 15700 4196
rect 15764 4168 16068 4196
rect 14884 4156 14890 4168
rect 13648 4112 13952 4128
rect 13648 4100 14044 4112
rect 13924 4084 14044 4100
rect 14090 4088 14096 4140
rect 14148 4128 14154 4140
rect 14921 4131 14979 4137
rect 14921 4128 14933 4131
rect 14148 4100 14933 4128
rect 14148 4088 14154 4100
rect 14921 4097 14933 4100
rect 14967 4097 14979 4131
rect 14921 4091 14979 4097
rect 15381 4131 15439 4137
rect 15381 4097 15393 4131
rect 15427 4128 15439 4131
rect 15764 4128 15792 4168
rect 16040 4140 16068 4168
rect 16224 4168 16764 4196
rect 15427 4100 15792 4128
rect 15841 4131 15899 4137
rect 15427 4097 15439 4100
rect 15381 4091 15439 4097
rect 15841 4097 15853 4131
rect 15887 4097 15899 4131
rect 15841 4091 15899 4097
rect 13814 4020 13820 4072
rect 13872 4020 13878 4072
rect 14016 4060 14044 4084
rect 14737 4063 14795 4069
rect 14737 4060 14749 4063
rect 14016 4032 14749 4060
rect 14737 4029 14749 4032
rect 14783 4029 14795 4063
rect 14737 4023 14795 4029
rect 14826 4020 14832 4072
rect 14884 4060 14890 4072
rect 15197 4063 15255 4069
rect 15197 4060 15209 4063
rect 14884 4032 15209 4060
rect 14884 4020 14890 4032
rect 15197 4029 15209 4032
rect 15243 4029 15255 4063
rect 15856 4060 15884 4091
rect 16022 4088 16028 4140
rect 16080 4088 16086 4140
rect 16224 4137 16252 4168
rect 16758 4156 16764 4168
rect 16816 4156 16822 4208
rect 17678 4156 17684 4208
rect 17736 4196 17742 4208
rect 18417 4199 18475 4205
rect 18417 4196 18429 4199
rect 17736 4168 18429 4196
rect 17736 4156 17742 4168
rect 18417 4165 18429 4168
rect 18463 4196 18475 4199
rect 20714 4196 20720 4208
rect 18463 4168 20720 4196
rect 18463 4165 18475 4168
rect 18417 4159 18475 4165
rect 20714 4156 20720 4168
rect 20772 4156 20778 4208
rect 20809 4199 20867 4205
rect 20809 4165 20821 4199
rect 20855 4196 20867 4199
rect 22296 4196 22324 4227
rect 23106 4224 23112 4236
rect 23164 4224 23170 4276
rect 23201 4267 23259 4273
rect 23201 4233 23213 4267
rect 23247 4264 23259 4267
rect 24578 4264 24584 4276
rect 23247 4236 24584 4264
rect 23247 4233 23259 4236
rect 23201 4227 23259 4233
rect 24578 4224 24584 4236
rect 24636 4264 24642 4276
rect 25317 4267 25375 4273
rect 25317 4264 25329 4267
rect 24636 4236 25329 4264
rect 24636 4224 24642 4236
rect 25317 4233 25329 4236
rect 25363 4233 25375 4267
rect 25317 4227 25375 4233
rect 25406 4224 25412 4276
rect 25464 4224 25470 4276
rect 25498 4224 25504 4276
rect 25556 4264 25562 4276
rect 29914 4264 29920 4276
rect 25556 4236 29920 4264
rect 25556 4224 25562 4236
rect 29914 4224 29920 4236
rect 29972 4224 29978 4276
rect 30837 4267 30895 4273
rect 30837 4233 30849 4267
rect 30883 4264 30895 4267
rect 35802 4264 35808 4276
rect 30883 4236 35808 4264
rect 30883 4233 30895 4236
rect 30837 4227 30895 4233
rect 35802 4224 35808 4236
rect 35860 4224 35866 4276
rect 20855 4168 22324 4196
rect 20855 4165 20867 4168
rect 20809 4159 20867 4165
rect 23014 4156 23020 4208
rect 23072 4196 23078 4208
rect 26234 4196 26240 4208
rect 23072 4168 26240 4196
rect 23072 4156 23078 4168
rect 26234 4156 26240 4168
rect 26292 4196 26298 4208
rect 26786 4196 26792 4208
rect 26292 4168 26792 4196
rect 26292 4156 26298 4168
rect 26786 4156 26792 4168
rect 26844 4156 26850 4208
rect 27890 4196 27896 4208
rect 26896 4168 27896 4196
rect 16209 4131 16267 4137
rect 16209 4097 16221 4131
rect 16255 4097 16267 4131
rect 16209 4091 16267 4097
rect 16301 4131 16359 4137
rect 16301 4097 16313 4131
rect 16347 4128 16359 4131
rect 16482 4128 16488 4140
rect 16347 4100 16488 4128
rect 16347 4097 16359 4100
rect 16301 4091 16359 4097
rect 15197 4023 15255 4029
rect 15580 4032 15884 4060
rect 14369 3995 14427 4001
rect 12544 3964 13133 3992
rect 5828 3896 8699 3924
rect 5445 3887 5503 3893
rect 8938 3884 8944 3936
rect 8996 3924 9002 3936
rect 9582 3924 9588 3936
rect 8996 3896 9588 3924
rect 8996 3884 9002 3896
rect 9582 3884 9588 3896
rect 9640 3884 9646 3936
rect 10413 3927 10471 3933
rect 10413 3893 10425 3927
rect 10459 3924 10471 3927
rect 10962 3924 10968 3936
rect 10459 3896 10968 3924
rect 10459 3893 10471 3896
rect 10413 3887 10471 3893
rect 10962 3884 10968 3896
rect 11020 3884 11026 3936
rect 11333 3927 11391 3933
rect 11333 3893 11345 3927
rect 11379 3924 11391 3927
rect 11698 3924 11704 3936
rect 11379 3896 11704 3924
rect 11379 3893 11391 3896
rect 11333 3887 11391 3893
rect 11698 3884 11704 3896
rect 11756 3884 11762 3936
rect 13105 3924 13133 3964
rect 14369 3961 14381 3995
rect 14415 3992 14427 3995
rect 15580 3992 15608 4032
rect 16114 4020 16120 4072
rect 16172 4020 16178 4072
rect 14415 3964 15608 3992
rect 14415 3961 14427 3964
rect 14369 3955 14427 3961
rect 16022 3952 16028 4004
rect 16080 3992 16086 4004
rect 16224 3992 16252 4091
rect 16482 4088 16488 4100
rect 16540 4088 16546 4140
rect 18322 4088 18328 4140
rect 18380 4128 18386 4140
rect 18380 4100 19104 4128
rect 18380 4088 18386 4100
rect 17954 4060 17960 4072
rect 16592 4032 17960 4060
rect 16592 3992 16620 4032
rect 17954 4020 17960 4032
rect 18012 4020 18018 4072
rect 18230 4020 18236 4072
rect 18288 4060 18294 4072
rect 18874 4060 18880 4072
rect 18288 4032 18880 4060
rect 18288 4020 18294 4032
rect 18874 4020 18880 4032
rect 18932 4020 18938 4072
rect 18966 4020 18972 4072
rect 19024 4020 19030 4072
rect 19076 4069 19104 4100
rect 19518 4088 19524 4140
rect 19576 4128 19582 4140
rect 19576 4100 23244 4128
rect 19576 4088 19582 4100
rect 19061 4063 19119 4069
rect 19061 4029 19073 4063
rect 19107 4029 19119 4063
rect 19061 4023 19119 4029
rect 20714 4020 20720 4072
rect 20772 4060 20778 4072
rect 20901 4063 20959 4069
rect 20901 4060 20913 4063
rect 20772 4032 20913 4060
rect 20772 4020 20778 4032
rect 20901 4029 20913 4032
rect 20947 4029 20959 4063
rect 20901 4023 20959 4029
rect 16080 3964 16252 3992
rect 16408 3964 16620 3992
rect 17129 3995 17187 4001
rect 16080 3952 16086 3964
rect 14553 3927 14611 3933
rect 14553 3924 14565 3927
rect 13105 3896 14565 3924
rect 14553 3893 14565 3896
rect 14599 3893 14611 3927
rect 14553 3887 14611 3893
rect 15105 3927 15163 3933
rect 15105 3893 15117 3927
rect 15151 3924 15163 3927
rect 16408 3924 16436 3964
rect 17129 3961 17141 3995
rect 17175 3992 17187 3995
rect 17862 3992 17868 4004
rect 17175 3964 17868 3992
rect 17175 3961 17187 3964
rect 17129 3955 17187 3961
rect 17862 3952 17868 3964
rect 17920 3952 17926 4004
rect 18984 3992 19012 4020
rect 18340 3964 19012 3992
rect 20441 3995 20499 4001
rect 18340 3936 18368 3964
rect 20441 3961 20453 3995
rect 20487 3992 20499 3995
rect 20806 3992 20812 4004
rect 20487 3964 20812 3992
rect 20487 3961 20499 3964
rect 20441 3955 20499 3961
rect 20806 3952 20812 3964
rect 20864 3952 20870 4004
rect 20916 3992 20944 4023
rect 20990 4020 20996 4072
rect 21048 4020 21054 4072
rect 22370 4060 22376 4072
rect 21284 4032 22376 4060
rect 21284 3992 21312 4032
rect 22370 4020 22376 4032
rect 22428 4020 22434 4072
rect 22462 4020 22468 4072
rect 22520 4020 22526 4072
rect 23106 4020 23112 4072
rect 23164 4020 23170 4072
rect 23216 4060 23244 4100
rect 23290 4088 23296 4140
rect 23348 4088 23354 4140
rect 23750 4088 23756 4140
rect 23808 4128 23814 4140
rect 23937 4131 23995 4137
rect 23937 4128 23949 4131
rect 23808 4100 23949 4128
rect 23808 4088 23814 4100
rect 23937 4097 23949 4100
rect 23983 4097 23995 4131
rect 23937 4091 23995 4097
rect 24394 4088 24400 4140
rect 24452 4088 24458 4140
rect 24670 4088 24676 4140
rect 24728 4128 24734 4140
rect 26896 4128 26924 4168
rect 27890 4156 27896 4168
rect 27948 4156 27954 4208
rect 27982 4156 27988 4208
rect 28040 4196 28046 4208
rect 28350 4196 28356 4208
rect 28040 4168 28356 4196
rect 28040 4156 28046 4168
rect 28350 4156 28356 4168
rect 28408 4156 28414 4208
rect 28902 4156 28908 4208
rect 28960 4156 28966 4208
rect 31662 4196 31668 4208
rect 29012 4168 31668 4196
rect 24728 4100 26924 4128
rect 27525 4131 27583 4137
rect 24728 4088 24734 4100
rect 27525 4097 27537 4131
rect 27571 4097 27583 4131
rect 27525 4091 27583 4097
rect 23216 4032 23805 4060
rect 20916 3964 21312 3992
rect 21358 3952 21364 4004
rect 21416 3992 21422 4004
rect 21821 3995 21879 4001
rect 21821 3992 21833 3995
rect 21416 3964 21833 3992
rect 21416 3952 21422 3964
rect 21821 3961 21833 3964
rect 21867 3961 21879 3995
rect 21821 3955 21879 3961
rect 15151 3896 16436 3924
rect 15151 3893 15163 3896
rect 15105 3887 15163 3893
rect 16482 3884 16488 3936
rect 16540 3884 16546 3936
rect 18322 3884 18328 3936
rect 18380 3884 18386 3936
rect 18509 3927 18567 3933
rect 18509 3893 18521 3927
rect 18555 3924 18567 3927
rect 18782 3924 18788 3936
rect 18555 3896 18788 3924
rect 18555 3893 18567 3896
rect 18509 3887 18567 3893
rect 18782 3884 18788 3896
rect 18840 3884 18846 3936
rect 18874 3884 18880 3936
rect 18932 3924 18938 3936
rect 22922 3924 22928 3936
rect 18932 3896 22928 3924
rect 18932 3884 18938 3896
rect 22922 3884 22928 3896
rect 22980 3884 22986 3936
rect 23658 3884 23664 3936
rect 23716 3884 23722 3936
rect 23777 3933 23805 4032
rect 25222 4020 25228 4072
rect 25280 4020 25286 4072
rect 25314 4020 25320 4072
rect 25372 4020 25378 4072
rect 26326 4020 26332 4072
rect 26384 4060 26390 4072
rect 27338 4060 27344 4072
rect 26384 4032 27344 4060
rect 26384 4020 26390 4032
rect 27338 4020 27344 4032
rect 27396 4020 27402 4072
rect 27540 4060 27568 4091
rect 27614 4088 27620 4140
rect 27672 4128 27678 4140
rect 28077 4131 28135 4137
rect 28077 4128 28089 4131
rect 27672 4100 28089 4128
rect 27672 4088 27678 4100
rect 28077 4097 28089 4100
rect 28123 4128 28135 4131
rect 29012 4128 29040 4168
rect 31662 4156 31668 4168
rect 31720 4156 31726 4208
rect 34974 4156 34980 4208
rect 35032 4196 35038 4208
rect 36357 4199 36415 4205
rect 36357 4196 36369 4199
rect 35032 4168 36369 4196
rect 35032 4156 35038 4168
rect 36357 4165 36369 4168
rect 36403 4165 36415 4199
rect 36357 4159 36415 4165
rect 28123 4100 29040 4128
rect 28123 4097 28135 4100
rect 28077 4091 28135 4097
rect 29914 4088 29920 4140
rect 29972 4128 29978 4140
rect 30193 4131 30251 4137
rect 30193 4128 30205 4131
rect 29972 4100 30205 4128
rect 29972 4088 29978 4100
rect 30193 4097 30205 4100
rect 30239 4128 30251 4131
rect 30377 4131 30435 4137
rect 30377 4128 30389 4131
rect 30239 4100 30389 4128
rect 30239 4097 30251 4100
rect 30193 4091 30251 4097
rect 30377 4097 30389 4100
rect 30423 4097 30435 4131
rect 30377 4091 30435 4097
rect 30650 4088 30656 4140
rect 30708 4088 30714 4140
rect 32398 4088 32404 4140
rect 32456 4088 32462 4140
rect 32858 4088 32864 4140
rect 32916 4128 32922 4140
rect 32953 4131 33011 4137
rect 32953 4128 32965 4131
rect 32916 4100 32965 4128
rect 32916 4088 32922 4100
rect 32953 4097 32965 4100
rect 32999 4097 33011 4131
rect 32953 4091 33011 4097
rect 33410 4088 33416 4140
rect 33468 4128 33474 4140
rect 34882 4128 34888 4140
rect 33468 4100 34888 4128
rect 33468 4088 33474 4100
rect 34882 4088 34888 4100
rect 34940 4088 34946 4140
rect 35161 4131 35219 4137
rect 35161 4097 35173 4131
rect 35207 4128 35219 4131
rect 35434 4128 35440 4140
rect 35207 4100 35440 4128
rect 35207 4097 35219 4100
rect 35161 4091 35219 4097
rect 35434 4088 35440 4100
rect 35492 4088 35498 4140
rect 36262 4088 36268 4140
rect 36320 4128 36326 4140
rect 36449 4131 36507 4137
rect 36449 4128 36461 4131
rect 36320 4100 36461 4128
rect 36320 4088 36326 4100
rect 36449 4097 36461 4100
rect 36495 4097 36507 4131
rect 36449 4091 36507 4097
rect 36630 4088 36636 4140
rect 36688 4128 36694 4140
rect 37553 4131 37611 4137
rect 37553 4128 37565 4131
rect 36688 4100 37565 4128
rect 36688 4088 36694 4100
rect 37553 4097 37565 4100
rect 37599 4097 37611 4131
rect 37553 4091 37611 4097
rect 38838 4088 38844 4140
rect 38896 4088 38902 4140
rect 39209 4131 39267 4137
rect 39209 4097 39221 4131
rect 39255 4128 39267 4131
rect 39574 4128 39580 4140
rect 39255 4100 39580 4128
rect 39255 4097 39267 4100
rect 39209 4091 39267 4097
rect 39574 4088 39580 4100
rect 39632 4088 39638 4140
rect 27540 4032 27660 4060
rect 26694 3952 26700 4004
rect 26752 3992 26758 4004
rect 27632 4001 27660 4032
rect 28258 4020 28264 4072
rect 28316 4020 28322 4072
rect 28445 4063 28503 4069
rect 28445 4029 28457 4063
rect 28491 4060 28503 4063
rect 28718 4060 28724 4072
rect 28491 4032 28724 4060
rect 28491 4029 28503 4032
rect 28445 4023 28503 4029
rect 28718 4020 28724 4032
rect 28776 4020 28782 4072
rect 30098 4020 30104 4072
rect 30156 4060 30162 4072
rect 31294 4060 31300 4072
rect 30156 4032 31300 4060
rect 30156 4020 30162 4032
rect 31294 4020 31300 4032
rect 31352 4020 31358 4072
rect 32582 4020 32588 4072
rect 32640 4060 32646 4072
rect 33778 4060 33784 4072
rect 32640 4032 33784 4060
rect 32640 4020 32646 4032
rect 33778 4020 33784 4032
rect 33836 4020 33842 4072
rect 36541 4063 36599 4069
rect 36541 4029 36553 4063
rect 36587 4029 36599 4063
rect 36541 4023 36599 4029
rect 27617 3995 27675 4001
rect 26752 3964 27568 3992
rect 26752 3952 26758 3964
rect 23753 3927 23811 3933
rect 23753 3893 23765 3927
rect 23799 3893 23811 3927
rect 23753 3887 23811 3893
rect 23934 3884 23940 3936
rect 23992 3924 23998 3936
rect 24213 3927 24271 3933
rect 24213 3924 24225 3927
rect 23992 3896 24225 3924
rect 23992 3884 23998 3896
rect 24213 3893 24225 3896
rect 24259 3893 24271 3927
rect 24213 3887 24271 3893
rect 25498 3884 25504 3936
rect 25556 3924 25562 3936
rect 25777 3927 25835 3933
rect 25777 3924 25789 3927
rect 25556 3896 25789 3924
rect 25556 3884 25562 3896
rect 25777 3893 25789 3896
rect 25823 3893 25835 3927
rect 25777 3887 25835 3893
rect 27338 3884 27344 3936
rect 27396 3884 27402 3936
rect 27540 3924 27568 3964
rect 27617 3961 27629 3995
rect 27663 3961 27675 3995
rect 27617 3955 27675 3961
rect 28537 3995 28595 4001
rect 28537 3961 28549 3995
rect 28583 3961 28595 3995
rect 28537 3955 28595 3961
rect 28552 3924 28580 3955
rect 28902 3952 28908 4004
rect 28960 3992 28966 4004
rect 30650 3992 30656 4004
rect 28960 3964 30656 3992
rect 28960 3952 28966 3964
rect 30650 3952 30656 3964
rect 30708 3952 30714 4004
rect 31754 3952 31760 4004
rect 31812 3992 31818 4004
rect 32217 3995 32275 4001
rect 32217 3992 32229 3995
rect 31812 3964 32229 3992
rect 31812 3952 31818 3964
rect 32217 3961 32229 3964
rect 32263 3961 32275 3995
rect 32217 3955 32275 3961
rect 35897 3995 35955 4001
rect 35897 3961 35909 3995
rect 35943 3992 35955 3995
rect 36556 3992 36584 4023
rect 35943 3964 36584 3992
rect 37369 3995 37427 4001
rect 35943 3961 35955 3964
rect 35897 3955 35955 3961
rect 37369 3961 37381 3995
rect 37415 3992 37427 3995
rect 37458 3992 37464 4004
rect 37415 3964 37464 3992
rect 37415 3961 37427 3964
rect 37369 3955 37427 3961
rect 37458 3952 37464 3964
rect 37516 3952 37522 4004
rect 39390 3952 39396 4004
rect 39448 3952 39454 4004
rect 27540 3896 28580 3924
rect 29730 3884 29736 3936
rect 29788 3884 29794 3936
rect 30101 3927 30159 3933
rect 30101 3893 30113 3927
rect 30147 3924 30159 3927
rect 30374 3924 30380 3936
rect 30147 3896 30380 3924
rect 30147 3893 30159 3896
rect 30101 3887 30159 3893
rect 30374 3884 30380 3896
rect 30432 3884 30438 3936
rect 30561 3927 30619 3933
rect 30561 3893 30573 3927
rect 30607 3924 30619 3927
rect 31110 3924 31116 3936
rect 30607 3896 31116 3924
rect 30607 3893 30619 3896
rect 30561 3887 30619 3893
rect 31110 3884 31116 3896
rect 31168 3884 31174 3936
rect 32766 3884 32772 3936
rect 32824 3884 32830 3936
rect 35986 3884 35992 3936
rect 36044 3884 36050 3936
rect 39022 3884 39028 3936
rect 39080 3884 39086 3936
rect 1104 3834 39836 3856
rect 1104 3782 1950 3834
rect 2002 3782 2014 3834
rect 2066 3782 2078 3834
rect 2130 3782 2142 3834
rect 2194 3782 2206 3834
rect 2258 3782 7950 3834
rect 8002 3782 8014 3834
rect 8066 3782 8078 3834
rect 8130 3782 8142 3834
rect 8194 3782 8206 3834
rect 8258 3782 13950 3834
rect 14002 3782 14014 3834
rect 14066 3782 14078 3834
rect 14130 3782 14142 3834
rect 14194 3782 14206 3834
rect 14258 3782 19950 3834
rect 20002 3782 20014 3834
rect 20066 3782 20078 3834
rect 20130 3782 20142 3834
rect 20194 3782 20206 3834
rect 20258 3782 25950 3834
rect 26002 3782 26014 3834
rect 26066 3782 26078 3834
rect 26130 3782 26142 3834
rect 26194 3782 26206 3834
rect 26258 3782 31950 3834
rect 32002 3782 32014 3834
rect 32066 3782 32078 3834
rect 32130 3782 32142 3834
rect 32194 3782 32206 3834
rect 32258 3782 37950 3834
rect 38002 3782 38014 3834
rect 38066 3782 38078 3834
rect 38130 3782 38142 3834
rect 38194 3782 38206 3834
rect 38258 3782 39836 3834
rect 1104 3760 39836 3782
rect 1302 3680 1308 3732
rect 1360 3720 1366 3732
rect 2777 3723 2835 3729
rect 1360 3692 2452 3720
rect 1360 3680 1366 3692
rect 1118 3612 1124 3664
rect 1176 3652 1182 3664
rect 1176 3624 1900 3652
rect 1176 3612 1182 3624
rect 382 3544 388 3596
rect 440 3584 446 3596
rect 440 3556 1808 3584
rect 440 3544 446 3556
rect 750 3476 756 3528
rect 808 3516 814 3528
rect 1780 3525 1808 3556
rect 1489 3519 1547 3525
rect 1489 3516 1501 3519
rect 808 3488 1501 3516
rect 808 3476 814 3488
rect 1489 3485 1501 3488
rect 1535 3485 1547 3519
rect 1489 3479 1547 3485
rect 1765 3519 1823 3525
rect 1765 3485 1777 3519
rect 1811 3485 1823 3519
rect 1872 3516 1900 3624
rect 1946 3612 1952 3664
rect 2004 3612 2010 3664
rect 2041 3519 2099 3525
rect 2041 3516 2053 3519
rect 1872 3488 2053 3516
rect 1765 3479 1823 3485
rect 2041 3485 2053 3488
rect 2087 3485 2099 3519
rect 2041 3479 2099 3485
rect 2314 3476 2320 3528
rect 2372 3476 2378 3528
rect 2424 3516 2452 3692
rect 2777 3689 2789 3723
rect 2823 3720 2835 3723
rect 2823 3692 5396 3720
rect 2823 3689 2835 3692
rect 2777 3683 2835 3689
rect 2501 3655 2559 3661
rect 2501 3621 2513 3655
rect 2547 3621 2559 3655
rect 2501 3615 2559 3621
rect 2516 3584 2544 3615
rect 2682 3612 2688 3664
rect 2740 3652 2746 3664
rect 3421 3655 3479 3661
rect 3421 3652 3433 3655
rect 2740 3624 3433 3652
rect 2740 3612 2746 3624
rect 3421 3621 3433 3624
rect 3467 3621 3479 3655
rect 3421 3615 3479 3621
rect 3786 3612 3792 3664
rect 3844 3652 3850 3664
rect 4338 3652 4344 3664
rect 3844 3624 4344 3652
rect 3844 3612 3850 3624
rect 4338 3612 4344 3624
rect 4396 3652 4402 3664
rect 4396 3624 4476 3652
rect 4396 3612 4402 3624
rect 4448 3593 4476 3624
rect 4433 3587 4491 3593
rect 2516 3556 4384 3584
rect 2593 3519 2651 3525
rect 2593 3516 2605 3519
rect 2424 3488 2605 3516
rect 2593 3485 2605 3488
rect 2639 3485 2651 3519
rect 2593 3479 2651 3485
rect 2682 3476 2688 3528
rect 2740 3516 2746 3528
rect 2869 3519 2927 3525
rect 2869 3516 2881 3519
rect 2740 3488 2881 3516
rect 2740 3476 2746 3488
rect 2869 3485 2881 3488
rect 2915 3485 2927 3519
rect 2869 3479 2927 3485
rect 3605 3519 3663 3525
rect 3605 3485 3617 3519
rect 3651 3516 3663 3519
rect 4356 3516 4384 3556
rect 4433 3553 4445 3587
rect 4479 3553 4491 3587
rect 5368 3584 5396 3692
rect 5442 3680 5448 3732
rect 5500 3680 5506 3732
rect 5721 3723 5779 3729
rect 5721 3689 5733 3723
rect 5767 3720 5779 3723
rect 5810 3720 5816 3732
rect 5767 3692 5816 3720
rect 5767 3689 5779 3692
rect 5721 3683 5779 3689
rect 5810 3680 5816 3692
rect 5868 3680 5874 3732
rect 5902 3680 5908 3732
rect 5960 3720 5966 3732
rect 7190 3720 7196 3732
rect 5960 3692 7196 3720
rect 5960 3680 5966 3692
rect 7190 3680 7196 3692
rect 7248 3720 7254 3732
rect 7248 3692 8340 3720
rect 7248 3680 7254 3692
rect 6638 3612 6644 3664
rect 6696 3652 6702 3664
rect 6696 3624 7696 3652
rect 6696 3612 6702 3624
rect 7668 3596 7696 3624
rect 5368 3556 7328 3584
rect 4433 3547 4491 3553
rect 3651 3488 4292 3516
rect 4356 3488 4660 3516
rect 3651 3485 3663 3488
rect 3605 3479 3663 3485
rect 1673 3451 1731 3457
rect 1673 3417 1685 3451
rect 1719 3448 1731 3451
rect 2774 3448 2780 3460
rect 1719 3420 2780 3448
rect 1719 3417 1731 3420
rect 1673 3411 1731 3417
rect 2774 3408 2780 3420
rect 2832 3408 2838 3460
rect 3881 3451 3939 3457
rect 3881 3448 3893 3451
rect 2884 3420 3893 3448
rect 2884 3392 2912 3420
rect 3881 3417 3893 3420
rect 3927 3417 3939 3451
rect 3881 3411 3939 3417
rect 1762 3340 1768 3392
rect 1820 3380 1826 3392
rect 2225 3383 2283 3389
rect 2225 3380 2237 3383
rect 1820 3352 2237 3380
rect 1820 3340 1826 3352
rect 2225 3349 2237 3352
rect 2271 3349 2283 3383
rect 2225 3343 2283 3349
rect 2866 3340 2872 3392
rect 2924 3340 2930 3392
rect 3050 3340 3056 3392
rect 3108 3340 3114 3392
rect 3421 3383 3479 3389
rect 3421 3349 3433 3383
rect 3467 3380 3479 3383
rect 3694 3380 3700 3392
rect 3467 3352 3700 3380
rect 3467 3349 3479 3352
rect 3421 3343 3479 3349
rect 3694 3340 3700 3352
rect 3752 3340 3758 3392
rect 3970 3340 3976 3392
rect 4028 3340 4034 3392
rect 4264 3380 4292 3488
rect 4632 3448 4660 3488
rect 4706 3476 4712 3528
rect 4764 3476 4770 3528
rect 5534 3476 5540 3528
rect 5592 3476 5598 3528
rect 7190 3448 7196 3460
rect 4632 3420 7196 3448
rect 7190 3408 7196 3420
rect 7248 3408 7254 3460
rect 7300 3448 7328 3556
rect 7466 3544 7472 3596
rect 7524 3584 7530 3596
rect 7561 3587 7619 3593
rect 7561 3584 7573 3587
rect 7524 3556 7573 3584
rect 7524 3544 7530 3556
rect 7561 3553 7573 3556
rect 7607 3553 7619 3587
rect 7561 3547 7619 3553
rect 7650 3544 7656 3596
rect 7708 3544 7714 3596
rect 8312 3584 8340 3692
rect 8386 3680 8392 3732
rect 8444 3720 8450 3732
rect 8941 3723 8999 3729
rect 8941 3720 8953 3723
rect 8444 3692 8953 3720
rect 8444 3680 8450 3692
rect 8941 3689 8953 3692
rect 8987 3689 8999 3723
rect 8941 3683 8999 3689
rect 9030 3680 9036 3732
rect 9088 3720 9094 3732
rect 10134 3720 10140 3732
rect 9088 3692 10140 3720
rect 9088 3680 9094 3692
rect 10134 3680 10140 3692
rect 10192 3680 10198 3732
rect 10778 3680 10784 3732
rect 10836 3720 10842 3732
rect 11425 3723 11483 3729
rect 11425 3720 11437 3723
rect 10836 3692 11437 3720
rect 10836 3680 10842 3692
rect 11425 3689 11437 3692
rect 11471 3689 11483 3723
rect 11425 3683 11483 3689
rect 11606 3680 11612 3732
rect 11664 3680 11670 3732
rect 13170 3680 13176 3732
rect 13228 3720 13234 3732
rect 13357 3723 13415 3729
rect 13357 3720 13369 3723
rect 13228 3692 13369 3720
rect 13228 3680 13234 3692
rect 13357 3689 13369 3692
rect 13403 3689 13415 3723
rect 13357 3683 13415 3689
rect 13722 3680 13728 3732
rect 13780 3720 13786 3732
rect 13780 3692 14320 3720
rect 13780 3680 13786 3692
rect 8665 3655 8723 3661
rect 8665 3621 8677 3655
rect 8711 3652 8723 3655
rect 8711 3624 9536 3652
rect 8711 3621 8723 3624
rect 8665 3615 8723 3621
rect 9508 3593 9536 3624
rect 13262 3612 13268 3664
rect 13320 3652 13326 3664
rect 14185 3655 14243 3661
rect 14185 3652 14197 3655
rect 13320 3624 14197 3652
rect 13320 3612 13326 3624
rect 14185 3621 14197 3624
rect 14231 3621 14243 3655
rect 14292 3652 14320 3692
rect 14458 3680 14464 3732
rect 14516 3680 14522 3732
rect 14734 3680 14740 3732
rect 14792 3720 14798 3732
rect 20714 3720 20720 3732
rect 14792 3692 20720 3720
rect 14792 3680 14798 3692
rect 20714 3680 20720 3692
rect 20772 3680 20778 3732
rect 20990 3680 20996 3732
rect 21048 3680 21054 3732
rect 23014 3720 23020 3732
rect 22204 3692 23020 3720
rect 16022 3652 16028 3664
rect 14292 3624 16028 3652
rect 14185 3615 14243 3621
rect 16022 3612 16028 3624
rect 16080 3612 16086 3664
rect 18230 3612 18236 3664
rect 18288 3652 18294 3664
rect 18325 3655 18383 3661
rect 18325 3652 18337 3655
rect 18288 3624 18337 3652
rect 18288 3612 18294 3624
rect 18325 3621 18337 3624
rect 18371 3621 18383 3655
rect 18325 3615 18383 3621
rect 19150 3612 19156 3664
rect 19208 3652 19214 3664
rect 20346 3652 20352 3664
rect 19208 3624 20352 3652
rect 19208 3612 19214 3624
rect 20346 3612 20352 3624
rect 20404 3652 20410 3664
rect 22204 3652 22232 3692
rect 23014 3680 23020 3692
rect 23072 3680 23078 3732
rect 23106 3680 23112 3732
rect 23164 3680 23170 3732
rect 24213 3723 24271 3729
rect 24213 3689 24225 3723
rect 24259 3720 24271 3723
rect 26329 3723 26387 3729
rect 24259 3692 24900 3720
rect 24259 3689 24271 3692
rect 24213 3683 24271 3689
rect 20404 3624 22232 3652
rect 20404 3612 20410 3624
rect 24486 3612 24492 3664
rect 24544 3612 24550 3664
rect 24765 3655 24823 3661
rect 24765 3621 24777 3655
rect 24811 3621 24823 3655
rect 24765 3615 24823 3621
rect 9493 3587 9551 3593
rect 8312 3556 9444 3584
rect 7374 3476 7380 3528
rect 7432 3516 7438 3528
rect 7929 3519 7987 3525
rect 7432 3512 7880 3516
rect 7929 3512 7941 3519
rect 7432 3488 7941 3512
rect 7432 3476 7438 3488
rect 7852 3485 7941 3488
rect 7975 3485 7987 3519
rect 7852 3484 7987 3485
rect 7929 3479 7987 3484
rect 8294 3476 8300 3528
rect 8352 3516 8358 3528
rect 9214 3516 9220 3528
rect 8352 3488 9220 3516
rect 8352 3476 8358 3488
rect 9214 3476 9220 3488
rect 9272 3476 9278 3528
rect 9306 3476 9312 3528
rect 9364 3476 9370 3528
rect 9416 3516 9444 3556
rect 9493 3553 9505 3587
rect 9539 3553 9551 3587
rect 9674 3584 9680 3596
rect 9493 3547 9551 3553
rect 9600 3556 9680 3584
rect 9600 3516 9628 3556
rect 9674 3544 9680 3556
rect 9732 3584 9738 3596
rect 10413 3587 10471 3593
rect 10413 3584 10425 3587
rect 9732 3556 10425 3584
rect 9732 3544 9738 3556
rect 10413 3553 10425 3556
rect 10459 3553 10471 3587
rect 10413 3547 10471 3553
rect 11422 3544 11428 3596
rect 11480 3584 11486 3596
rect 11480 3556 11744 3584
rect 11480 3544 11486 3556
rect 10594 3516 10600 3528
rect 9416 3488 9628 3516
rect 10152 3488 10600 3516
rect 10152 3457 10180 3488
rect 10594 3476 10600 3488
rect 10652 3516 10658 3528
rect 10689 3519 10747 3525
rect 10689 3516 10701 3519
rect 10652 3488 10701 3516
rect 10652 3476 10658 3488
rect 10689 3485 10701 3488
rect 10735 3485 10747 3519
rect 10689 3479 10747 3485
rect 11054 3476 11060 3528
rect 11112 3516 11118 3528
rect 11716 3525 11744 3556
rect 11882 3544 11888 3596
rect 11940 3544 11946 3596
rect 13722 3584 13728 3596
rect 13096 3556 13728 3584
rect 13096 3528 13124 3556
rect 13722 3544 13728 3556
rect 13780 3544 13786 3596
rect 14458 3584 14464 3596
rect 13924 3556 14464 3584
rect 11517 3519 11575 3525
rect 11517 3516 11529 3519
rect 11112 3488 11529 3516
rect 11112 3476 11118 3488
rect 11517 3485 11529 3488
rect 11563 3485 11575 3519
rect 11517 3479 11575 3485
rect 11701 3519 11759 3525
rect 11701 3485 11713 3519
rect 11747 3516 11759 3519
rect 13078 3516 13084 3528
rect 11747 3488 13084 3516
rect 11747 3485 11759 3488
rect 11701 3479 11759 3485
rect 13078 3476 13084 3488
rect 13136 3476 13142 3528
rect 13446 3476 13452 3528
rect 13504 3516 13510 3528
rect 13924 3525 13952 3556
rect 14458 3544 14464 3556
rect 14516 3544 14522 3596
rect 15013 3587 15071 3593
rect 15013 3553 15025 3587
rect 15059 3553 15071 3587
rect 15013 3547 15071 3553
rect 13541 3519 13599 3525
rect 13541 3516 13553 3519
rect 13504 3488 13553 3516
rect 13504 3476 13510 3488
rect 13541 3485 13553 3488
rect 13587 3485 13599 3519
rect 13541 3479 13599 3485
rect 13909 3519 13967 3525
rect 13909 3485 13921 3519
rect 13955 3485 13967 3519
rect 13909 3479 13967 3485
rect 14274 3476 14280 3528
rect 14332 3516 14338 3528
rect 14369 3519 14427 3525
rect 14369 3516 14381 3519
rect 14332 3488 14381 3516
rect 14332 3476 14338 3488
rect 14369 3485 14381 3488
rect 14415 3516 14427 3519
rect 14734 3516 14740 3528
rect 14415 3488 14740 3516
rect 14415 3485 14427 3488
rect 14369 3479 14427 3485
rect 14734 3476 14740 3488
rect 14792 3476 14798 3528
rect 14826 3476 14832 3528
rect 14884 3476 14890 3528
rect 12158 3457 12164 3460
rect 10137 3451 10195 3457
rect 10137 3448 10149 3451
rect 7300 3420 10149 3448
rect 10137 3417 10149 3420
rect 10183 3417 10195 3451
rect 10137 3411 10195 3417
rect 10336 3420 12112 3448
rect 10336 3392 10364 3420
rect 5350 3380 5356 3392
rect 4264 3352 5356 3380
rect 5350 3340 5356 3352
rect 5408 3380 5414 3392
rect 7742 3380 7748 3392
rect 5408 3352 7748 3380
rect 5408 3340 5414 3352
rect 7742 3340 7748 3352
rect 7800 3380 7806 3392
rect 9306 3380 9312 3392
rect 7800 3352 9312 3380
rect 7800 3340 7806 3352
rect 9306 3340 9312 3352
rect 9364 3340 9370 3392
rect 9401 3383 9459 3389
rect 9401 3349 9413 3383
rect 9447 3380 9459 3383
rect 9490 3380 9496 3392
rect 9447 3352 9496 3380
rect 9447 3349 9459 3352
rect 9401 3343 9459 3349
rect 9490 3340 9496 3352
rect 9548 3340 9554 3392
rect 10226 3340 10232 3392
rect 10284 3340 10290 3392
rect 10318 3340 10324 3392
rect 10376 3340 10382 3392
rect 10778 3340 10784 3392
rect 10836 3380 10842 3392
rect 11974 3380 11980 3392
rect 10836 3352 11980 3380
rect 10836 3340 10842 3352
rect 11974 3340 11980 3352
rect 12032 3340 12038 3392
rect 12084 3380 12112 3420
rect 12152 3411 12164 3457
rect 12216 3448 12222 3460
rect 12216 3420 12252 3448
rect 12158 3408 12164 3411
rect 12216 3408 12222 3420
rect 12342 3408 12348 3460
rect 12400 3448 12406 3460
rect 12400 3420 13768 3448
rect 12400 3408 12406 3420
rect 12250 3380 12256 3392
rect 12084 3352 12256 3380
rect 12250 3340 12256 3352
rect 12308 3380 12314 3392
rect 13265 3383 13323 3389
rect 13265 3380 13277 3383
rect 12308 3352 13277 3380
rect 12308 3340 12314 3352
rect 13265 3349 13277 3352
rect 13311 3380 13323 3383
rect 13630 3380 13636 3392
rect 13311 3352 13636 3380
rect 13311 3349 13323 3352
rect 13265 3343 13323 3349
rect 13630 3340 13636 3352
rect 13688 3340 13694 3392
rect 13740 3389 13768 3420
rect 14090 3408 14096 3460
rect 14148 3448 14154 3460
rect 15028 3448 15056 3547
rect 15378 3544 15384 3596
rect 15436 3584 15442 3596
rect 17586 3584 17592 3596
rect 15436 3556 17592 3584
rect 15436 3544 15442 3556
rect 17586 3544 17592 3556
rect 17644 3544 17650 3596
rect 18966 3584 18972 3596
rect 18248 3556 18972 3584
rect 18248 3528 18276 3556
rect 18966 3544 18972 3556
rect 19024 3584 19030 3596
rect 19702 3584 19708 3596
rect 19024 3556 19708 3584
rect 19024 3544 19030 3556
rect 19702 3544 19708 3556
rect 19760 3544 19766 3596
rect 15102 3476 15108 3528
rect 15160 3516 15166 3528
rect 15289 3519 15347 3525
rect 15289 3516 15301 3519
rect 15160 3488 15301 3516
rect 15160 3476 15166 3488
rect 15289 3485 15301 3488
rect 15335 3485 15347 3519
rect 15289 3479 15347 3485
rect 14148 3420 15056 3448
rect 15304 3448 15332 3479
rect 15838 3476 15844 3528
rect 15896 3476 15902 3528
rect 16942 3476 16948 3528
rect 17000 3476 17006 3528
rect 17954 3476 17960 3528
rect 18012 3476 18018 3528
rect 18230 3476 18236 3528
rect 18288 3476 18294 3528
rect 18506 3476 18512 3528
rect 18564 3476 18570 3528
rect 18782 3476 18788 3528
rect 18840 3476 18846 3528
rect 19058 3476 19064 3528
rect 19116 3476 19122 3528
rect 20809 3519 20867 3525
rect 20809 3516 20821 3519
rect 19306 3488 20821 3516
rect 17972 3448 18000 3476
rect 19306 3448 19334 3488
rect 20809 3485 20821 3488
rect 20855 3485 20867 3519
rect 20809 3479 20867 3485
rect 21269 3519 21327 3525
rect 21269 3485 21281 3519
rect 21315 3516 21327 3519
rect 21358 3516 21364 3528
rect 21315 3488 21364 3516
rect 21315 3485 21327 3488
rect 21269 3479 21327 3485
rect 15304 3420 17908 3448
rect 17972 3420 19334 3448
rect 20824 3448 20852 3479
rect 21358 3476 21364 3488
rect 21416 3476 21422 3528
rect 21450 3476 21456 3528
rect 21508 3476 21514 3528
rect 22094 3476 22100 3528
rect 22152 3476 22158 3528
rect 22373 3519 22431 3525
rect 22373 3485 22385 3519
rect 22419 3485 22431 3519
rect 22373 3479 22431 3485
rect 23201 3519 23259 3525
rect 23201 3485 23213 3519
rect 23247 3485 23259 3519
rect 23201 3479 23259 3485
rect 22388 3448 22416 3479
rect 20824 3420 22416 3448
rect 23216 3448 23244 3479
rect 23474 3476 23480 3528
rect 23532 3476 23538 3528
rect 24673 3519 24731 3525
rect 24673 3485 24685 3519
rect 24719 3516 24731 3519
rect 24780 3516 24808 3615
rect 24872 3584 24900 3692
rect 26329 3689 26341 3723
rect 26375 3720 26387 3723
rect 27522 3720 27528 3732
rect 26375 3692 27528 3720
rect 26375 3689 26387 3692
rect 26329 3683 26387 3689
rect 27522 3680 27528 3692
rect 27580 3680 27586 3732
rect 28258 3680 28264 3732
rect 28316 3720 28322 3732
rect 28905 3723 28963 3729
rect 28905 3720 28917 3723
rect 28316 3692 28917 3720
rect 28316 3680 28322 3692
rect 28905 3689 28917 3692
rect 28951 3689 28963 3723
rect 28905 3683 28963 3689
rect 29181 3723 29239 3729
rect 29181 3689 29193 3723
rect 29227 3720 29239 3723
rect 38378 3720 38384 3732
rect 29227 3692 32444 3720
rect 29227 3689 29239 3692
rect 29181 3683 29239 3689
rect 25406 3612 25412 3664
rect 25464 3652 25470 3664
rect 25958 3652 25964 3664
rect 25464 3624 25964 3652
rect 25464 3612 25470 3624
rect 25958 3612 25964 3624
rect 26016 3612 26022 3664
rect 30650 3612 30656 3664
rect 30708 3652 30714 3664
rect 30929 3655 30987 3661
rect 30929 3652 30941 3655
rect 30708 3624 30941 3652
rect 30708 3612 30714 3624
rect 30929 3621 30941 3624
rect 30975 3621 30987 3655
rect 32416 3652 32444 3692
rect 32784 3692 38384 3720
rect 32784 3652 32812 3692
rect 38378 3680 38384 3692
rect 38436 3680 38442 3732
rect 32416 3624 32812 3652
rect 30929 3615 30987 3621
rect 32858 3612 32864 3664
rect 32916 3652 32922 3664
rect 38838 3652 38844 3664
rect 32916 3624 38844 3652
rect 32916 3612 32922 3624
rect 38838 3612 38844 3624
rect 38896 3612 38902 3664
rect 39390 3612 39396 3664
rect 39448 3612 39454 3664
rect 25317 3587 25375 3593
rect 25317 3584 25329 3587
rect 24872 3556 25329 3584
rect 25317 3553 25329 3556
rect 25363 3553 25375 3587
rect 25317 3547 25375 3553
rect 25774 3544 25780 3596
rect 25832 3544 25838 3596
rect 25869 3587 25927 3593
rect 25869 3553 25881 3587
rect 25915 3584 25927 3587
rect 26510 3584 26516 3596
rect 25915 3556 26516 3584
rect 25915 3553 25927 3556
rect 25869 3547 25927 3553
rect 24719 3488 24808 3516
rect 25133 3519 25191 3525
rect 24719 3485 24731 3488
rect 24673 3479 24731 3485
rect 25133 3485 25145 3519
rect 25179 3516 25191 3519
rect 25884 3516 25912 3547
rect 26510 3544 26516 3556
rect 26568 3544 26574 3596
rect 26786 3544 26792 3596
rect 26844 3544 26850 3596
rect 27706 3544 27712 3596
rect 27764 3584 27770 3596
rect 27893 3587 27951 3593
rect 27893 3584 27905 3587
rect 27764 3556 27905 3584
rect 27764 3544 27770 3556
rect 27893 3553 27905 3556
rect 27939 3553 27951 3587
rect 27893 3547 27951 3553
rect 30561 3587 30619 3593
rect 30561 3553 30573 3587
rect 30607 3584 30619 3587
rect 31110 3584 31116 3596
rect 30607 3556 31116 3584
rect 30607 3553 30619 3556
rect 30561 3547 30619 3553
rect 31110 3544 31116 3556
rect 31168 3544 31174 3596
rect 35250 3544 35256 3596
rect 35308 3584 35314 3596
rect 35308 3556 36124 3584
rect 35308 3544 35314 3556
rect 25179 3488 25912 3516
rect 25179 3485 25191 3488
rect 25133 3479 25191 3485
rect 25958 3476 25964 3528
rect 26016 3476 26022 3528
rect 27065 3519 27123 3525
rect 27065 3485 27077 3519
rect 27111 3485 27123 3519
rect 27065 3479 27123 3485
rect 24210 3448 24216 3460
rect 23216 3420 24216 3448
rect 14148 3408 14154 3420
rect 13725 3383 13783 3389
rect 13725 3349 13737 3383
rect 13771 3349 13783 3383
rect 13725 3343 13783 3349
rect 13998 3340 14004 3392
rect 14056 3380 14062 3392
rect 14921 3383 14979 3389
rect 14921 3380 14933 3383
rect 14056 3352 14933 3380
rect 14056 3340 14062 3352
rect 14921 3349 14933 3352
rect 14967 3380 14979 3383
rect 15378 3380 15384 3392
rect 14967 3352 15384 3380
rect 14967 3349 14979 3352
rect 14921 3343 14979 3349
rect 15378 3340 15384 3352
rect 15436 3340 15442 3392
rect 15470 3340 15476 3392
rect 15528 3340 15534 3392
rect 15654 3340 15660 3392
rect 15712 3340 15718 3392
rect 17126 3340 17132 3392
rect 17184 3340 17190 3392
rect 17218 3340 17224 3392
rect 17276 3340 17282 3392
rect 17880 3380 17908 3420
rect 18230 3380 18236 3392
rect 17880 3352 18236 3380
rect 18230 3340 18236 3352
rect 18288 3340 18294 3392
rect 18506 3340 18512 3392
rect 18564 3380 18570 3392
rect 18601 3383 18659 3389
rect 18601 3380 18613 3383
rect 18564 3352 18613 3380
rect 18564 3340 18570 3352
rect 18601 3349 18613 3352
rect 18647 3349 18659 3383
rect 18601 3343 18659 3349
rect 18690 3340 18696 3392
rect 18748 3380 18754 3392
rect 18877 3383 18935 3389
rect 18877 3380 18889 3383
rect 18748 3352 18889 3380
rect 18748 3340 18754 3352
rect 18877 3349 18889 3352
rect 18923 3349 18935 3383
rect 18877 3343 18935 3349
rect 19334 3340 19340 3392
rect 19392 3380 19398 3392
rect 21085 3383 21143 3389
rect 21085 3380 21097 3383
rect 19392 3352 21097 3380
rect 19392 3340 19398 3352
rect 21085 3349 21097 3352
rect 21131 3349 21143 3383
rect 21085 3343 21143 3349
rect 21634 3340 21640 3392
rect 21692 3340 21698 3392
rect 22094 3340 22100 3392
rect 22152 3380 22158 3392
rect 23216 3380 23244 3420
rect 24210 3408 24216 3420
rect 24268 3408 24274 3460
rect 25225 3451 25283 3457
rect 25225 3417 25237 3451
rect 25271 3448 25283 3451
rect 25314 3448 25320 3460
rect 25271 3420 25320 3448
rect 25271 3417 25283 3420
rect 25225 3411 25283 3417
rect 25314 3408 25320 3420
rect 25372 3408 25378 3460
rect 25406 3408 25412 3460
rect 25464 3448 25470 3460
rect 25464 3420 26096 3448
rect 25464 3408 25470 3420
rect 22152 3352 23244 3380
rect 26068 3380 26096 3420
rect 26142 3408 26148 3460
rect 26200 3448 26206 3460
rect 27080 3448 27108 3479
rect 28166 3476 28172 3528
rect 28224 3516 28230 3528
rect 28997 3519 29055 3525
rect 28997 3516 29009 3519
rect 28224 3488 29009 3516
rect 28224 3476 28230 3488
rect 28997 3485 29009 3488
rect 29043 3516 29055 3519
rect 30285 3519 30343 3525
rect 30285 3516 30297 3519
rect 29043 3488 30297 3516
rect 29043 3485 29055 3488
rect 28997 3479 29055 3485
rect 30285 3485 30297 3488
rect 30331 3485 30343 3519
rect 30285 3479 30343 3485
rect 31570 3476 31576 3528
rect 31628 3516 31634 3528
rect 31665 3519 31723 3525
rect 31665 3516 31677 3519
rect 31628 3488 31677 3516
rect 31628 3476 31634 3488
rect 31665 3485 31677 3488
rect 31711 3485 31723 3519
rect 31665 3479 31723 3485
rect 31938 3476 31944 3528
rect 31996 3476 32002 3528
rect 32306 3476 32312 3528
rect 32364 3516 32370 3528
rect 32677 3519 32735 3525
rect 32677 3516 32689 3519
rect 32364 3488 32689 3516
rect 32364 3476 32370 3488
rect 32677 3485 32689 3488
rect 32723 3485 32735 3519
rect 32677 3479 32735 3485
rect 35897 3519 35955 3525
rect 35897 3485 35909 3519
rect 35943 3516 35955 3519
rect 35986 3516 35992 3528
rect 35943 3488 35992 3516
rect 35943 3485 35955 3488
rect 35897 3479 35955 3485
rect 35986 3476 35992 3488
rect 36044 3476 36050 3528
rect 36096 3516 36124 3556
rect 37274 3544 37280 3596
rect 37332 3584 37338 3596
rect 37332 3556 39252 3584
rect 37332 3544 37338 3556
rect 39224 3525 39252 3556
rect 38841 3519 38899 3525
rect 38841 3516 38853 3519
rect 36096 3488 38853 3516
rect 38841 3485 38853 3488
rect 38887 3485 38899 3519
rect 38841 3479 38899 3485
rect 39209 3519 39267 3525
rect 39209 3485 39221 3519
rect 39255 3485 39267 3519
rect 39209 3479 39267 3485
rect 38470 3448 38476 3460
rect 26200 3420 27108 3448
rect 27172 3420 38476 3448
rect 26200 3408 26206 3420
rect 27172 3380 27200 3420
rect 38470 3408 38476 3420
rect 38528 3408 38534 3460
rect 26068 3352 27200 3380
rect 27801 3383 27859 3389
rect 22152 3340 22158 3352
rect 27801 3349 27813 3383
rect 27847 3380 27859 3383
rect 28442 3380 28448 3392
rect 27847 3352 28448 3380
rect 27847 3349 27859 3352
rect 27801 3343 27859 3349
rect 28442 3340 28448 3352
rect 28500 3340 28506 3392
rect 29549 3383 29607 3389
rect 29549 3349 29561 3383
rect 29595 3380 29607 3383
rect 29638 3380 29644 3392
rect 29595 3352 29644 3380
rect 29595 3349 29607 3352
rect 29549 3343 29607 3349
rect 29638 3340 29644 3352
rect 29696 3340 29702 3392
rect 30190 3340 30196 3392
rect 30248 3380 30254 3392
rect 32214 3380 32220 3392
rect 30248 3352 32220 3380
rect 30248 3340 30254 3352
rect 32214 3340 32220 3352
rect 32272 3340 32278 3392
rect 32493 3383 32551 3389
rect 32493 3349 32505 3383
rect 32539 3380 32551 3383
rect 32950 3380 32956 3392
rect 32539 3352 32956 3380
rect 32539 3349 32551 3352
rect 32493 3343 32551 3349
rect 32950 3340 32956 3352
rect 33008 3340 33014 3392
rect 33962 3340 33968 3392
rect 34020 3380 34026 3392
rect 34422 3380 34428 3392
rect 34020 3352 34428 3380
rect 34020 3340 34026 3352
rect 34422 3340 34428 3352
rect 34480 3340 34486 3392
rect 35802 3340 35808 3392
rect 35860 3340 35866 3392
rect 39025 3383 39083 3389
rect 39025 3349 39037 3383
rect 39071 3380 39083 3383
rect 39942 3380 39948 3392
rect 39071 3352 39948 3380
rect 39071 3349 39083 3352
rect 39025 3343 39083 3349
rect 39942 3340 39948 3352
rect 40000 3340 40006 3392
rect 1104 3290 39836 3312
rect 1104 3238 3010 3290
rect 3062 3238 3074 3290
rect 3126 3238 3138 3290
rect 3190 3238 3202 3290
rect 3254 3238 3266 3290
rect 3318 3238 9010 3290
rect 9062 3238 9074 3290
rect 9126 3238 9138 3290
rect 9190 3238 9202 3290
rect 9254 3238 9266 3290
rect 9318 3238 15010 3290
rect 15062 3238 15074 3290
rect 15126 3238 15138 3290
rect 15190 3238 15202 3290
rect 15254 3238 15266 3290
rect 15318 3238 21010 3290
rect 21062 3238 21074 3290
rect 21126 3238 21138 3290
rect 21190 3238 21202 3290
rect 21254 3238 21266 3290
rect 21318 3238 27010 3290
rect 27062 3238 27074 3290
rect 27126 3238 27138 3290
rect 27190 3238 27202 3290
rect 27254 3238 27266 3290
rect 27318 3238 33010 3290
rect 33062 3238 33074 3290
rect 33126 3238 33138 3290
rect 33190 3238 33202 3290
rect 33254 3238 33266 3290
rect 33318 3238 39010 3290
rect 39062 3238 39074 3290
rect 39126 3238 39138 3290
rect 39190 3238 39202 3290
rect 39254 3238 39266 3290
rect 39318 3238 39836 3290
rect 1104 3216 39836 3238
rect 1673 3179 1731 3185
rect 1673 3145 1685 3179
rect 1719 3145 1731 3179
rect 1673 3139 1731 3145
rect 1026 3068 1032 3120
rect 1084 3108 1090 3120
rect 1688 3108 1716 3139
rect 1946 3136 1952 3188
rect 2004 3176 2010 3188
rect 6733 3179 6791 3185
rect 2004 3148 6684 3176
rect 2004 3136 2010 3148
rect 4706 3108 4712 3120
rect 1084 3080 1624 3108
rect 1688 3080 4712 3108
rect 1084 3068 1090 3080
rect 566 3000 572 3052
rect 624 3040 630 3052
rect 1489 3043 1547 3049
rect 1489 3040 1501 3043
rect 624 3012 1501 3040
rect 624 3000 630 3012
rect 1489 3009 1501 3012
rect 1535 3009 1547 3043
rect 1596 3040 1624 3080
rect 4706 3068 4712 3080
rect 4764 3068 4770 3120
rect 6656 3108 6684 3148
rect 6733 3145 6745 3179
rect 6779 3176 6791 3179
rect 6822 3176 6828 3188
rect 6779 3148 6828 3176
rect 6779 3145 6791 3148
rect 6733 3139 6791 3145
rect 6822 3136 6828 3148
rect 6880 3136 6886 3188
rect 7190 3136 7196 3188
rect 7248 3176 7254 3188
rect 7926 3176 7932 3188
rect 7248 3148 7932 3176
rect 7248 3136 7254 3148
rect 7926 3136 7932 3148
rect 7984 3136 7990 3188
rect 8478 3136 8484 3188
rect 8536 3176 8542 3188
rect 8536 3148 9674 3176
rect 8536 3136 8542 3148
rect 9646 3108 9674 3148
rect 9950 3136 9956 3188
rect 10008 3136 10014 3188
rect 10134 3136 10140 3188
rect 10192 3176 10198 3188
rect 10778 3176 10784 3188
rect 10192 3148 10784 3176
rect 10192 3136 10198 3148
rect 10778 3136 10784 3148
rect 10836 3136 10842 3188
rect 11517 3179 11575 3185
rect 11517 3145 11529 3179
rect 11563 3176 11575 3179
rect 11790 3176 11796 3188
rect 11563 3148 11796 3176
rect 11563 3145 11575 3148
rect 11517 3139 11575 3145
rect 11790 3136 11796 3148
rect 11848 3136 11854 3188
rect 11882 3136 11888 3188
rect 11940 3176 11946 3188
rect 13630 3176 13636 3188
rect 11940 3148 13636 3176
rect 11940 3136 11946 3148
rect 13630 3136 13636 3148
rect 13688 3136 13694 3188
rect 13814 3136 13820 3188
rect 13872 3176 13878 3188
rect 13909 3179 13967 3185
rect 13909 3176 13921 3179
rect 13872 3148 13921 3176
rect 13872 3136 13878 3148
rect 13909 3145 13921 3148
rect 13955 3145 13967 3179
rect 13909 3139 13967 3145
rect 13998 3136 14004 3188
rect 14056 3176 14062 3188
rect 14550 3176 14556 3188
rect 14056 3148 14556 3176
rect 14056 3136 14062 3148
rect 14550 3136 14556 3148
rect 14608 3136 14614 3188
rect 16022 3136 16028 3188
rect 16080 3176 16086 3188
rect 17037 3179 17095 3185
rect 17037 3176 17049 3179
rect 16080 3148 17049 3176
rect 16080 3136 16086 3148
rect 17037 3145 17049 3148
rect 17083 3145 17095 3179
rect 17037 3139 17095 3145
rect 17129 3179 17187 3185
rect 17129 3145 17141 3179
rect 17175 3176 17187 3179
rect 23842 3176 23848 3188
rect 17175 3148 23848 3176
rect 17175 3145 17187 3148
rect 17129 3139 17187 3145
rect 23842 3136 23848 3148
rect 23900 3136 23906 3188
rect 24118 3136 24124 3188
rect 24176 3136 24182 3188
rect 25222 3136 25228 3188
rect 25280 3136 25286 3188
rect 25317 3179 25375 3185
rect 25317 3145 25329 3179
rect 25363 3145 25375 3179
rect 25317 3139 25375 3145
rect 6656 3080 9076 3108
rect 9646 3080 10732 3108
rect 1765 3043 1823 3049
rect 1765 3040 1777 3043
rect 1596 3012 1777 3040
rect 1489 3003 1547 3009
rect 1765 3009 1777 3012
rect 1811 3009 1823 3043
rect 2041 3043 2099 3049
rect 2041 3040 2053 3043
rect 1765 3003 1823 3009
rect 1872 3012 2053 3040
rect 474 2932 480 2984
rect 532 2972 538 2984
rect 1872 2972 1900 3012
rect 2041 3009 2053 3012
rect 2087 3009 2099 3043
rect 2041 3003 2099 3009
rect 2314 3000 2320 3052
rect 2372 3000 2378 3052
rect 2590 3000 2596 3052
rect 2648 3000 2654 3052
rect 2682 3000 2688 3052
rect 2740 3040 2746 3052
rect 2869 3043 2927 3049
rect 2869 3040 2881 3043
rect 2740 3012 2881 3040
rect 2740 3000 2746 3012
rect 2869 3009 2881 3012
rect 2915 3009 2927 3043
rect 4724 3040 4752 3068
rect 5261 3043 5319 3049
rect 5261 3040 5273 3043
rect 4724 3012 5273 3040
rect 2869 3003 2927 3009
rect 5261 3009 5273 3012
rect 5307 3009 5319 3043
rect 5261 3003 5319 3009
rect 6825 3043 6883 3049
rect 6825 3009 6837 3043
rect 6871 3040 6883 3043
rect 7466 3040 7472 3052
rect 6871 3012 7472 3040
rect 6871 3009 6883 3012
rect 6825 3003 6883 3009
rect 7466 3000 7472 3012
rect 7524 3000 7530 3052
rect 7561 3043 7619 3049
rect 7561 3009 7573 3043
rect 7607 3040 7619 3043
rect 7742 3040 7748 3052
rect 7607 3012 7748 3040
rect 7607 3009 7619 3012
rect 7561 3003 7619 3009
rect 7742 3000 7748 3012
rect 7800 3000 7806 3052
rect 7837 3043 7895 3049
rect 7837 3009 7849 3043
rect 7883 3040 7895 3043
rect 7926 3040 7932 3052
rect 7883 3012 7932 3040
rect 7883 3009 7895 3012
rect 7837 3003 7895 3009
rect 7926 3000 7932 3012
rect 7984 3040 7990 3052
rect 8570 3040 8576 3052
rect 7984 3012 8576 3040
rect 7984 3000 7990 3012
rect 8570 3000 8576 3012
rect 8628 3040 8634 3052
rect 8941 3043 8999 3049
rect 8941 3040 8953 3043
rect 8628 3012 8953 3040
rect 8628 3000 8634 3012
rect 8941 3009 8953 3012
rect 8987 3009 8999 3043
rect 9048 3040 9076 3080
rect 9048 3012 9674 3040
rect 8941 3003 8999 3009
rect 3602 2972 3608 2984
rect 532 2944 1900 2972
rect 1964 2944 3608 2972
rect 532 2932 538 2944
rect 1964 2913 1992 2944
rect 3602 2932 3608 2944
rect 3660 2932 3666 2984
rect 3694 2932 3700 2984
rect 3752 2972 3758 2984
rect 4985 2975 5043 2981
rect 4985 2972 4997 2975
rect 3752 2944 4997 2972
rect 3752 2932 3758 2944
rect 4985 2941 4997 2944
rect 5031 2941 5043 2975
rect 4985 2935 5043 2941
rect 1949 2907 2007 2913
rect 1949 2873 1961 2907
rect 1995 2873 2007 2907
rect 1949 2867 2007 2873
rect 2225 2907 2283 2913
rect 2225 2873 2237 2907
rect 2271 2904 2283 2907
rect 2406 2904 2412 2916
rect 2271 2876 2412 2904
rect 2271 2873 2283 2876
rect 2225 2867 2283 2873
rect 2406 2864 2412 2876
rect 2464 2864 2470 2916
rect 2501 2907 2559 2913
rect 2501 2873 2513 2907
rect 2547 2904 2559 2907
rect 4062 2904 4068 2916
rect 2547 2876 4068 2904
rect 2547 2873 2559 2876
rect 2501 2867 2559 2873
rect 4062 2864 4068 2876
rect 4120 2864 4126 2916
rect 4890 2864 4896 2916
rect 4948 2864 4954 2916
rect 5000 2904 5028 2935
rect 6914 2932 6920 2984
rect 6972 2932 6978 2984
rect 8478 2932 8484 2984
rect 8536 2972 8542 2984
rect 8665 2975 8723 2981
rect 8665 2972 8677 2975
rect 8536 2944 8677 2972
rect 8536 2932 8542 2944
rect 8665 2941 8677 2944
rect 8711 2941 8723 2975
rect 9646 2972 9674 3012
rect 9766 3000 9772 3052
rect 9824 3000 9830 3052
rect 10321 3043 10379 3049
rect 10321 3009 10333 3043
rect 10367 3040 10379 3043
rect 10502 3040 10508 3052
rect 10367 3012 10508 3040
rect 10367 3009 10379 3012
rect 10321 3003 10379 3009
rect 10502 3000 10508 3012
rect 10560 3000 10566 3052
rect 10594 3000 10600 3052
rect 10652 3000 10658 3052
rect 10704 3040 10732 3080
rect 12084 3080 14320 3108
rect 11606 3040 11612 3052
rect 10704 3012 11612 3040
rect 11606 3000 11612 3012
rect 11664 3000 11670 3052
rect 11698 3000 11704 3052
rect 11756 3000 11762 3052
rect 11790 3000 11796 3052
rect 11848 3000 11854 3052
rect 11974 3000 11980 3052
rect 12032 3040 12038 3052
rect 12084 3049 12112 3080
rect 12069 3043 12127 3049
rect 12069 3040 12081 3043
rect 12032 3012 12081 3040
rect 12032 3000 12038 3012
rect 12069 3009 12081 3012
rect 12115 3009 12127 3043
rect 12069 3003 12127 3009
rect 12894 3000 12900 3052
rect 12952 3000 12958 3052
rect 13170 3000 13176 3052
rect 13228 3000 13234 3052
rect 14292 3049 14320 3080
rect 14642 3068 14648 3120
rect 14700 3108 14706 3120
rect 16114 3108 16120 3120
rect 14700 3080 16120 3108
rect 14700 3068 14706 3080
rect 16114 3068 16120 3080
rect 16172 3068 16178 3120
rect 17218 3108 17224 3120
rect 17052 3080 17224 3108
rect 14277 3043 14335 3049
rect 14277 3009 14289 3043
rect 14323 3009 14335 3043
rect 14277 3003 14335 3009
rect 14826 3000 14832 3052
rect 14884 3040 14890 3052
rect 15381 3043 15439 3049
rect 15381 3040 15393 3043
rect 14884 3012 15393 3040
rect 14884 3000 14890 3012
rect 15381 3009 15393 3012
rect 15427 3009 15439 3043
rect 17052 3040 17080 3080
rect 17218 3068 17224 3080
rect 17276 3068 17282 3120
rect 19426 3068 19432 3120
rect 19484 3108 19490 3120
rect 19484 3080 20852 3108
rect 19484 3068 19490 3080
rect 15381 3003 15439 3009
rect 16960 3012 17080 3040
rect 17236 3012 17724 3040
rect 10134 2972 10140 2984
rect 9646 2944 10140 2972
rect 8665 2935 8723 2941
rect 10134 2932 10140 2944
rect 10192 2932 10198 2984
rect 13538 2932 13544 2984
rect 13596 2972 13602 2984
rect 13906 2972 13912 2984
rect 13596 2944 13912 2972
rect 13596 2932 13602 2944
rect 13906 2932 13912 2944
rect 13964 2932 13970 2984
rect 13998 2932 14004 2984
rect 14056 2932 14062 2984
rect 14918 2932 14924 2984
rect 14976 2972 14982 2984
rect 16960 2981 16988 3012
rect 15105 2975 15163 2981
rect 15105 2972 15117 2975
rect 14976 2944 15117 2972
rect 14976 2932 14982 2944
rect 15105 2941 15117 2944
rect 15151 2941 15163 2975
rect 15105 2935 15163 2941
rect 16945 2975 17003 2981
rect 16945 2941 16957 2975
rect 16991 2941 17003 2975
rect 16945 2935 17003 2941
rect 17037 2975 17095 2981
rect 17037 2941 17049 2975
rect 17083 2972 17095 2975
rect 17236 2972 17264 3012
rect 17083 2944 17264 2972
rect 17083 2941 17095 2944
rect 17037 2935 17095 2941
rect 17494 2932 17500 2984
rect 17552 2932 17558 2984
rect 17586 2932 17592 2984
rect 17644 2932 17650 2984
rect 5997 2907 6055 2913
rect 5000 2876 5120 2904
rect 2777 2839 2835 2845
rect 2777 2805 2789 2839
rect 2823 2836 2835 2839
rect 2866 2836 2872 2848
rect 2823 2808 2872 2836
rect 2823 2805 2835 2808
rect 2777 2799 2835 2805
rect 2866 2796 2872 2808
rect 2924 2796 2930 2848
rect 3053 2839 3111 2845
rect 3053 2805 3065 2839
rect 3099 2836 3111 2839
rect 3786 2836 3792 2848
rect 3099 2808 3792 2836
rect 3099 2805 3111 2808
rect 3053 2799 3111 2805
rect 3786 2796 3792 2808
rect 3844 2796 3850 2848
rect 5092 2836 5120 2876
rect 5997 2873 6009 2907
rect 6043 2904 6055 2907
rect 6043 2876 6500 2904
rect 6043 2873 6055 2876
rect 5997 2867 6055 2873
rect 5902 2836 5908 2848
rect 5092 2808 5908 2836
rect 5902 2796 5908 2808
rect 5960 2796 5966 2848
rect 6178 2796 6184 2848
rect 6236 2836 6242 2848
rect 6365 2839 6423 2845
rect 6365 2836 6377 2839
rect 6236 2808 6377 2836
rect 6236 2796 6242 2808
rect 6365 2805 6377 2808
rect 6411 2805 6423 2839
rect 6472 2836 6500 2876
rect 13630 2864 13636 2916
rect 13688 2904 13694 2916
rect 13688 2876 14136 2904
rect 13688 2864 13694 2876
rect 6914 2836 6920 2848
rect 6472 2808 6920 2836
rect 6365 2799 6423 2805
rect 6914 2796 6920 2808
rect 6972 2796 6978 2848
rect 8573 2839 8631 2845
rect 8573 2805 8585 2839
rect 8619 2836 8631 2839
rect 9030 2836 9036 2848
rect 8619 2808 9036 2836
rect 8619 2805 8631 2808
rect 8573 2799 8631 2805
rect 9030 2796 9036 2808
rect 9088 2796 9094 2848
rect 9677 2839 9735 2845
rect 9677 2805 9689 2839
rect 9723 2836 9735 2839
rect 11054 2836 11060 2848
rect 9723 2808 11060 2836
rect 9723 2805 9735 2808
rect 9677 2799 9735 2805
rect 11054 2796 11060 2808
rect 11112 2796 11118 2848
rect 11330 2796 11336 2848
rect 11388 2796 11394 2848
rect 12805 2839 12863 2845
rect 12805 2805 12817 2839
rect 12851 2836 12863 2839
rect 13722 2836 13728 2848
rect 12851 2808 13728 2836
rect 12851 2805 12863 2808
rect 12805 2799 12863 2805
rect 13722 2796 13728 2808
rect 13780 2796 13786 2848
rect 14108 2836 14136 2876
rect 14734 2836 14740 2848
rect 14108 2808 14740 2836
rect 14734 2796 14740 2808
rect 14792 2836 14798 2848
rect 14945 2836 14973 2932
rect 16117 2907 16175 2913
rect 16117 2873 16129 2907
rect 16163 2904 16175 2907
rect 17512 2904 17540 2932
rect 16163 2876 17540 2904
rect 16163 2873 16175 2876
rect 16117 2867 16175 2873
rect 14792 2808 14973 2836
rect 14792 2796 14798 2808
rect 15010 2796 15016 2848
rect 15068 2796 15074 2848
rect 17494 2796 17500 2848
rect 17552 2796 17558 2848
rect 17696 2836 17724 3012
rect 17770 3000 17776 3052
rect 17828 3000 17834 3052
rect 18782 3000 18788 3052
rect 18840 3000 18846 3052
rect 19702 3000 19708 3052
rect 19760 3040 19766 3052
rect 19797 3043 19855 3049
rect 19797 3040 19809 3043
rect 19760 3012 19809 3040
rect 19760 3000 19766 3012
rect 19797 3009 19809 3012
rect 19843 3009 19855 3043
rect 19797 3003 19855 3009
rect 20346 3000 20352 3052
rect 20404 3040 20410 3052
rect 20441 3043 20499 3049
rect 20441 3040 20453 3043
rect 20404 3012 20453 3040
rect 20404 3000 20410 3012
rect 20441 3009 20453 3012
rect 20487 3009 20499 3043
rect 20441 3003 20499 3009
rect 20714 3000 20720 3052
rect 20772 3000 20778 3052
rect 20824 3040 20852 3080
rect 20898 3068 20904 3120
rect 20956 3108 20962 3120
rect 21818 3108 21824 3120
rect 20956 3080 21824 3108
rect 20956 3068 20962 3080
rect 21818 3068 21824 3080
rect 21876 3108 21882 3120
rect 21876 3080 23980 3108
rect 21876 3068 21882 3080
rect 21450 3040 21456 3052
rect 20824 3012 21456 3040
rect 21450 3000 21456 3012
rect 21508 3040 21514 3052
rect 22281 3043 22339 3049
rect 22281 3040 22293 3043
rect 21508 3012 22293 3040
rect 21508 3000 21514 3012
rect 22281 3009 22293 3012
rect 22327 3009 22339 3043
rect 22281 3003 22339 3009
rect 23382 3000 23388 3052
rect 23440 3040 23446 3052
rect 23952 3049 23980 3080
rect 25130 3068 25136 3120
rect 25188 3108 25194 3120
rect 25332 3108 25360 3139
rect 25774 3136 25780 3188
rect 25832 3176 25838 3188
rect 28534 3176 28540 3188
rect 25832 3148 28540 3176
rect 25832 3136 25838 3148
rect 28534 3136 28540 3148
rect 28592 3136 28598 3188
rect 29917 3179 29975 3185
rect 29917 3145 29929 3179
rect 29963 3176 29975 3179
rect 30098 3176 30104 3188
rect 29963 3148 30104 3176
rect 29963 3145 29975 3148
rect 29917 3139 29975 3145
rect 30098 3136 30104 3148
rect 30156 3136 30162 3188
rect 30285 3179 30343 3185
rect 30285 3145 30297 3179
rect 30331 3145 30343 3179
rect 30285 3139 30343 3145
rect 30377 3179 30435 3185
rect 30377 3145 30389 3179
rect 30423 3176 30435 3179
rect 30558 3176 30564 3188
rect 30423 3148 30564 3176
rect 30423 3145 30435 3148
rect 30377 3139 30435 3145
rect 25188 3080 25360 3108
rect 25188 3068 25194 3080
rect 26142 3068 26148 3120
rect 26200 3108 26206 3120
rect 26200 3080 27752 3108
rect 26200 3068 26206 3080
rect 23477 3043 23535 3049
rect 23477 3040 23489 3043
rect 23440 3012 23489 3040
rect 23440 3000 23446 3012
rect 23477 3009 23489 3012
rect 23523 3009 23535 3043
rect 23477 3003 23535 3009
rect 23937 3043 23995 3049
rect 23937 3009 23949 3043
rect 23983 3040 23995 3043
rect 24489 3043 24547 3049
rect 24489 3040 24501 3043
rect 23983 3012 24501 3040
rect 23983 3009 23995 3012
rect 23937 3003 23995 3009
rect 24489 3009 24501 3012
rect 24535 3009 24547 3043
rect 24489 3003 24547 3009
rect 25498 3000 25504 3052
rect 25556 3000 25562 3052
rect 25774 3000 25780 3052
rect 25832 3040 25838 3052
rect 26326 3040 26332 3052
rect 25832 3012 26332 3040
rect 25832 3000 25838 3012
rect 26326 3000 26332 3012
rect 26384 3000 26390 3052
rect 26786 3000 26792 3052
rect 26844 3000 26850 3052
rect 27724 3049 27752 3080
rect 28626 3068 28632 3120
rect 28684 3108 28690 3120
rect 29825 3111 29883 3117
rect 29825 3108 29837 3111
rect 28684 3080 29837 3108
rect 28684 3068 28690 3080
rect 29825 3077 29837 3080
rect 29871 3077 29883 3111
rect 29825 3071 29883 3077
rect 27709 3043 27767 3049
rect 27709 3009 27721 3043
rect 27755 3040 27767 3043
rect 28077 3043 28135 3049
rect 28077 3040 28089 3043
rect 27755 3012 28089 3040
rect 27755 3009 27767 3012
rect 27709 3003 27767 3009
rect 28077 3009 28089 3012
rect 28123 3009 28135 3043
rect 28077 3003 28135 3009
rect 28534 3000 28540 3052
rect 28592 3040 28598 3052
rect 30300 3040 30328 3139
rect 30558 3136 30564 3148
rect 30616 3136 30622 3188
rect 30742 3136 30748 3188
rect 30800 3176 30806 3188
rect 32858 3176 32864 3188
rect 30800 3148 32864 3176
rect 30800 3136 30806 3148
rect 32858 3136 32864 3148
rect 32916 3136 32922 3188
rect 34885 3179 34943 3185
rect 34885 3176 34897 3179
rect 32968 3148 34897 3176
rect 31202 3068 31208 3120
rect 31260 3108 31266 3120
rect 31478 3108 31484 3120
rect 31260 3080 31484 3108
rect 31260 3068 31266 3080
rect 31478 3068 31484 3080
rect 31536 3108 31542 3120
rect 31938 3108 31944 3120
rect 31536 3080 31944 3108
rect 31536 3068 31542 3080
rect 31938 3068 31944 3080
rect 31996 3068 32002 3120
rect 32214 3068 32220 3120
rect 32272 3108 32278 3120
rect 32272 3080 32904 3108
rect 32272 3068 32278 3080
rect 32876 3052 32904 3080
rect 30561 3043 30619 3049
rect 30561 3040 30573 3043
rect 28592 3012 29960 3040
rect 30300 3012 30573 3040
rect 28592 3000 28598 3012
rect 18322 2932 18328 2984
rect 18380 2972 18386 2984
rect 18509 2975 18567 2981
rect 18509 2972 18521 2975
rect 18380 2944 18521 2972
rect 18380 2932 18386 2944
rect 18509 2941 18521 2944
rect 18555 2941 18567 2975
rect 18509 2935 18567 2941
rect 18647 2975 18705 2981
rect 18647 2941 18659 2975
rect 18693 2972 18705 2975
rect 19521 2975 19579 2981
rect 18693 2944 19196 2972
rect 18693 2941 18705 2944
rect 18647 2935 18705 2941
rect 18230 2864 18236 2916
rect 18288 2864 18294 2916
rect 19168 2836 19196 2944
rect 19521 2941 19533 2975
rect 19567 2941 19579 2975
rect 19521 2935 19579 2941
rect 19242 2864 19248 2916
rect 19300 2904 19306 2916
rect 19536 2904 19564 2935
rect 22002 2932 22008 2984
rect 22060 2932 22066 2984
rect 23566 2932 23572 2984
rect 23624 2932 23630 2984
rect 23661 2975 23719 2981
rect 23661 2941 23673 2975
rect 23707 2941 23719 2975
rect 23661 2935 23719 2941
rect 20346 2904 20352 2916
rect 19300 2876 20352 2904
rect 19300 2864 19306 2876
rect 20346 2864 20352 2876
rect 20404 2864 20410 2916
rect 23017 2907 23075 2913
rect 23017 2873 23029 2907
rect 23063 2904 23075 2907
rect 23676 2904 23704 2935
rect 24210 2932 24216 2984
rect 24268 2932 24274 2984
rect 27985 2975 28043 2981
rect 27985 2941 27997 2975
rect 28031 2941 28043 2975
rect 27985 2935 28043 2941
rect 23063 2876 23704 2904
rect 24228 2904 24256 2932
rect 24228 2876 24348 2904
rect 23063 2873 23075 2876
rect 23017 2867 23075 2873
rect 17696 2808 19196 2836
rect 19426 2796 19432 2848
rect 19484 2796 19490 2848
rect 21450 2796 21456 2848
rect 21508 2796 21514 2848
rect 23109 2839 23167 2845
rect 23109 2805 23121 2839
rect 23155 2836 23167 2839
rect 23198 2836 23204 2848
rect 23155 2808 23204 2836
rect 23155 2805 23167 2808
rect 23109 2799 23167 2805
rect 23198 2796 23204 2808
rect 23256 2796 23262 2848
rect 24320 2836 24348 2876
rect 24872 2876 27384 2904
rect 24872 2836 24900 2876
rect 24320 2808 24900 2836
rect 25958 2796 25964 2848
rect 26016 2796 26022 2848
rect 26602 2796 26608 2848
rect 26660 2796 26666 2848
rect 26973 2839 27031 2845
rect 26973 2805 26985 2839
rect 27019 2836 27031 2839
rect 27246 2836 27252 2848
rect 27019 2808 27252 2836
rect 27019 2805 27031 2808
rect 26973 2799 27031 2805
rect 27246 2796 27252 2808
rect 27304 2796 27310 2848
rect 27356 2836 27384 2876
rect 28000 2836 28028 2935
rect 29638 2932 29644 2984
rect 29696 2932 29702 2984
rect 29932 2972 29960 3012
rect 30561 3009 30573 3012
rect 30607 3009 30619 3043
rect 30561 3003 30619 3009
rect 31570 3000 31576 3052
rect 31628 3000 31634 3052
rect 31662 3000 31668 3052
rect 31720 3040 31726 3052
rect 32401 3043 32459 3049
rect 32401 3040 32413 3043
rect 31720 3012 32413 3040
rect 31720 3000 31726 3012
rect 32401 3009 32413 3012
rect 32447 3009 32459 3043
rect 32401 3003 32459 3009
rect 32858 3000 32864 3052
rect 32916 3000 32922 3052
rect 31849 2975 31907 2981
rect 29932 2944 30880 2972
rect 28261 2907 28319 2913
rect 28261 2873 28273 2907
rect 28307 2904 28319 2907
rect 30742 2904 30748 2916
rect 28307 2876 30748 2904
rect 28307 2873 28319 2876
rect 28261 2867 28319 2873
rect 30742 2864 30748 2876
rect 30800 2864 30806 2916
rect 30852 2913 30880 2944
rect 31849 2941 31861 2975
rect 31895 2972 31907 2975
rect 31938 2972 31944 2984
rect 31895 2944 31944 2972
rect 31895 2941 31907 2944
rect 31849 2935 31907 2941
rect 31938 2932 31944 2944
rect 31996 2932 32002 2984
rect 32122 2932 32128 2984
rect 32180 2932 32186 2984
rect 32968 2972 32996 3148
rect 34885 3145 34897 3148
rect 34931 3145 34943 3179
rect 34885 3139 34943 3145
rect 34977 3179 35035 3185
rect 34977 3145 34989 3179
rect 35023 3176 35035 3179
rect 36262 3176 36268 3188
rect 35023 3148 36268 3176
rect 35023 3145 35035 3148
rect 34977 3139 35035 3145
rect 36262 3136 36268 3148
rect 36320 3136 36326 3188
rect 36817 3179 36875 3185
rect 36817 3145 36829 3179
rect 36863 3176 36875 3179
rect 37366 3176 37372 3188
rect 36863 3148 37372 3176
rect 36863 3145 36875 3148
rect 36817 3139 36875 3145
rect 37366 3136 37372 3148
rect 37424 3136 37430 3188
rect 39390 3136 39396 3188
rect 39448 3136 39454 3188
rect 33042 3068 33048 3120
rect 33100 3108 33106 3120
rect 33100 3080 33824 3108
rect 33100 3068 33106 3080
rect 33410 3000 33416 3052
rect 33468 3000 33474 3052
rect 33686 3000 33692 3052
rect 33744 3000 33750 3052
rect 33796 3040 33824 3080
rect 34238 3068 34244 3120
rect 34296 3108 34302 3120
rect 34296 3080 35388 3108
rect 34296 3068 34302 3080
rect 35360 3049 35388 3080
rect 36372 3080 39252 3108
rect 35345 3043 35403 3049
rect 33796 3012 35204 3040
rect 34977 2975 35035 2981
rect 34977 2972 34989 2975
rect 32784 2944 32996 2972
rect 34072 2944 34989 2972
rect 30837 2907 30895 2913
rect 30837 2873 30849 2907
rect 30883 2873 30895 2907
rect 30837 2867 30895 2873
rect 30374 2836 30380 2848
rect 27356 2808 30380 2836
rect 30374 2796 30380 2808
rect 30432 2796 30438 2848
rect 30466 2796 30472 2848
rect 30524 2836 30530 2848
rect 32784 2836 32812 2944
rect 32858 2864 32864 2916
rect 32916 2904 32922 2916
rect 32916 2876 33272 2904
rect 32916 2864 32922 2876
rect 30524 2808 32812 2836
rect 30524 2796 30530 2808
rect 33042 2796 33048 2848
rect 33100 2836 33106 2848
rect 33137 2839 33195 2845
rect 33137 2836 33149 2839
rect 33100 2808 33149 2836
rect 33100 2796 33106 2808
rect 33137 2805 33149 2808
rect 33183 2805 33195 2839
rect 33244 2836 33272 2876
rect 34072 2836 34100 2944
rect 34977 2941 34989 2944
rect 35023 2941 35035 2975
rect 34977 2935 35035 2941
rect 35069 2975 35127 2981
rect 35069 2941 35081 2975
rect 35115 2941 35127 2975
rect 35176 2972 35204 3012
rect 35345 3009 35357 3043
rect 35391 3009 35403 3043
rect 35345 3003 35403 3009
rect 36372 2972 36400 3080
rect 36633 3043 36691 3049
rect 36633 3009 36645 3043
rect 36679 3009 36691 3043
rect 36633 3003 36691 3009
rect 38749 3043 38807 3049
rect 38749 3009 38761 3043
rect 38795 3009 38807 3043
rect 38749 3003 38807 3009
rect 35176 2944 36400 2972
rect 35069 2935 35127 2941
rect 34330 2864 34336 2916
rect 34388 2904 34394 2916
rect 34517 2907 34575 2913
rect 34517 2904 34529 2907
rect 34388 2876 34529 2904
rect 34388 2864 34394 2876
rect 34517 2873 34529 2876
rect 34563 2873 34575 2907
rect 35084 2904 35112 2935
rect 34517 2867 34575 2873
rect 34624 2876 35112 2904
rect 35529 2907 35587 2913
rect 33244 2808 34100 2836
rect 34425 2839 34483 2845
rect 33137 2799 33195 2805
rect 34425 2805 34437 2839
rect 34471 2836 34483 2839
rect 34624 2836 34652 2876
rect 35529 2873 35541 2907
rect 35575 2904 35587 2907
rect 35710 2904 35716 2916
rect 35575 2876 35716 2904
rect 35575 2873 35587 2876
rect 35529 2867 35587 2873
rect 35710 2864 35716 2876
rect 35768 2864 35774 2916
rect 36648 2904 36676 3003
rect 38764 2972 38792 3003
rect 38838 3000 38844 3052
rect 38896 3000 38902 3052
rect 39224 3049 39252 3080
rect 39209 3043 39267 3049
rect 39209 3009 39221 3043
rect 39255 3009 39267 3043
rect 39209 3003 39267 3009
rect 39482 2972 39488 2984
rect 38764 2944 39488 2972
rect 39482 2932 39488 2944
rect 39540 2932 39546 2984
rect 39758 2904 39764 2916
rect 36648 2876 39764 2904
rect 39758 2864 39764 2876
rect 39816 2864 39822 2916
rect 34471 2808 34652 2836
rect 34471 2805 34483 2808
rect 34425 2799 34483 2805
rect 34698 2796 34704 2848
rect 34756 2836 34762 2848
rect 38565 2839 38623 2845
rect 38565 2836 38577 2839
rect 34756 2808 38577 2836
rect 34756 2796 34762 2808
rect 38565 2805 38577 2808
rect 38611 2805 38623 2839
rect 38565 2799 38623 2805
rect 39022 2796 39028 2848
rect 39080 2796 39086 2848
rect 1104 2746 39836 2768
rect 1104 2694 1950 2746
rect 2002 2694 2014 2746
rect 2066 2694 2078 2746
rect 2130 2694 2142 2746
rect 2194 2694 2206 2746
rect 2258 2694 7950 2746
rect 8002 2694 8014 2746
rect 8066 2694 8078 2746
rect 8130 2694 8142 2746
rect 8194 2694 8206 2746
rect 8258 2694 13950 2746
rect 14002 2694 14014 2746
rect 14066 2694 14078 2746
rect 14130 2694 14142 2746
rect 14194 2694 14206 2746
rect 14258 2694 19950 2746
rect 20002 2694 20014 2746
rect 20066 2694 20078 2746
rect 20130 2694 20142 2746
rect 20194 2694 20206 2746
rect 20258 2694 25950 2746
rect 26002 2694 26014 2746
rect 26066 2694 26078 2746
rect 26130 2694 26142 2746
rect 26194 2694 26206 2746
rect 26258 2694 31950 2746
rect 32002 2694 32014 2746
rect 32066 2694 32078 2746
rect 32130 2694 32142 2746
rect 32194 2694 32206 2746
rect 32258 2694 37950 2746
rect 38002 2694 38014 2746
rect 38066 2694 38078 2746
rect 38130 2694 38142 2746
rect 38194 2694 38206 2746
rect 38258 2694 39836 2746
rect 1104 2672 39836 2694
rect 1578 2592 1584 2644
rect 1636 2632 1642 2644
rect 1762 2632 1768 2644
rect 1636 2604 1768 2632
rect 1636 2592 1642 2604
rect 1762 2592 1768 2604
rect 1820 2592 1826 2644
rect 1949 2635 2007 2641
rect 1949 2601 1961 2635
rect 1995 2632 2007 2635
rect 4706 2632 4712 2644
rect 1995 2604 4712 2632
rect 1995 2601 2007 2604
rect 1949 2595 2007 2601
rect 4706 2592 4712 2604
rect 4764 2592 4770 2644
rect 5994 2592 6000 2644
rect 6052 2592 6058 2644
rect 10505 2635 10563 2641
rect 10505 2632 10517 2635
rect 7484 2604 10517 2632
rect 1118 2524 1124 2576
rect 1176 2564 1182 2576
rect 1176 2536 3004 2564
rect 1176 2524 1182 2536
rect 1302 2456 1308 2508
rect 1360 2496 1366 2508
rect 1360 2468 2728 2496
rect 1360 2456 1366 2468
rect 934 2388 940 2440
rect 992 2428 998 2440
rect 1857 2431 1915 2437
rect 1857 2428 1869 2431
rect 992 2400 1869 2428
rect 992 2388 998 2400
rect 1857 2397 1869 2400
rect 1903 2397 1915 2431
rect 1857 2391 1915 2397
rect 2225 2431 2283 2437
rect 2225 2397 2237 2431
rect 2271 2428 2283 2431
rect 2590 2428 2596 2440
rect 2271 2400 2596 2428
rect 2271 2397 2283 2400
rect 2225 2391 2283 2397
rect 2590 2388 2596 2400
rect 2648 2388 2654 2440
rect 2700 2437 2728 2468
rect 2976 2437 3004 2536
rect 3878 2524 3884 2576
rect 3936 2564 3942 2576
rect 7484 2564 7512 2604
rect 10505 2601 10517 2604
rect 10551 2601 10563 2635
rect 10505 2595 10563 2601
rect 11054 2592 11060 2644
rect 11112 2632 11118 2644
rect 11517 2635 11575 2641
rect 11517 2632 11529 2635
rect 11112 2604 11529 2632
rect 11112 2592 11118 2604
rect 11517 2601 11529 2604
rect 11563 2601 11575 2635
rect 11517 2595 11575 2601
rect 13173 2635 13231 2641
rect 13173 2601 13185 2635
rect 13219 2632 13231 2635
rect 13446 2632 13452 2644
rect 13219 2604 13452 2632
rect 13219 2601 13231 2604
rect 13173 2595 13231 2601
rect 13446 2592 13452 2604
rect 13504 2592 13510 2644
rect 14550 2632 14556 2644
rect 13556 2604 14556 2632
rect 10318 2564 10324 2576
rect 3936 2536 7512 2564
rect 8036 2536 10324 2564
rect 3936 2524 3942 2536
rect 4522 2456 4528 2508
rect 4580 2496 4586 2508
rect 4706 2496 4712 2508
rect 4580 2468 4712 2496
rect 4580 2456 4586 2468
rect 4706 2456 4712 2468
rect 4764 2456 4770 2508
rect 2685 2431 2743 2437
rect 2685 2397 2697 2431
rect 2731 2397 2743 2431
rect 2685 2391 2743 2397
rect 2961 2431 3019 2437
rect 2961 2397 2973 2431
rect 3007 2397 3019 2431
rect 2961 2391 3019 2397
rect 4062 2388 4068 2440
rect 4120 2388 4126 2440
rect 4798 2388 4804 2440
rect 4856 2388 4862 2440
rect 5902 2388 5908 2440
rect 5960 2388 5966 2440
rect 6178 2388 6184 2440
rect 6236 2388 6242 2440
rect 7006 2388 7012 2440
rect 7064 2388 7070 2440
rect 7466 2388 7472 2440
rect 7524 2428 7530 2440
rect 8036 2437 8064 2536
rect 10318 2524 10324 2536
rect 10376 2524 10382 2576
rect 10962 2524 10968 2576
rect 11020 2524 11026 2576
rect 11606 2524 11612 2576
rect 11664 2564 11670 2576
rect 13556 2564 13584 2604
rect 14550 2592 14556 2604
rect 14608 2592 14614 2644
rect 14642 2592 14648 2644
rect 14700 2632 14706 2644
rect 15470 2632 15476 2644
rect 14700 2604 15476 2632
rect 14700 2592 14706 2604
rect 15470 2592 15476 2604
rect 15528 2592 15534 2644
rect 15749 2635 15807 2641
rect 15749 2601 15761 2635
rect 15795 2632 15807 2635
rect 15838 2632 15844 2644
rect 15795 2604 15844 2632
rect 15795 2601 15807 2604
rect 15749 2595 15807 2601
rect 15838 2592 15844 2604
rect 15896 2592 15902 2644
rect 17957 2635 18015 2641
rect 17957 2601 17969 2635
rect 18003 2632 18015 2635
rect 18230 2632 18236 2644
rect 18003 2604 18236 2632
rect 18003 2601 18015 2604
rect 17957 2595 18015 2601
rect 18230 2592 18236 2604
rect 18288 2592 18294 2644
rect 21358 2592 21364 2644
rect 21416 2632 21422 2644
rect 21545 2635 21603 2641
rect 21545 2632 21557 2635
rect 21416 2604 21557 2632
rect 21416 2592 21422 2604
rect 21545 2601 21557 2604
rect 21591 2601 21603 2635
rect 21545 2595 21603 2601
rect 22922 2592 22928 2644
rect 22980 2592 22986 2644
rect 26786 2592 26792 2644
rect 26844 2632 26850 2644
rect 26973 2635 27031 2641
rect 26973 2632 26985 2635
rect 26844 2604 26985 2632
rect 26844 2592 26850 2604
rect 26973 2601 26985 2604
rect 27019 2601 27031 2635
rect 29454 2632 29460 2644
rect 26973 2595 27031 2601
rect 27080 2604 29460 2632
rect 17034 2564 17040 2576
rect 11664 2536 13584 2564
rect 14016 2536 17040 2564
rect 11664 2524 11670 2536
rect 8404 2468 8984 2496
rect 8404 2437 8432 2468
rect 8021 2431 8079 2437
rect 7524 2400 7972 2428
rect 7524 2388 7530 2400
rect 382 2320 388 2372
rect 440 2360 446 2372
rect 1489 2363 1547 2369
rect 1489 2360 1501 2363
rect 440 2332 1501 2360
rect 440 2320 446 2332
rect 1489 2329 1501 2332
rect 1535 2329 1547 2363
rect 7650 2360 7656 2372
rect 1489 2323 1547 2329
rect 3160 2332 7656 2360
rect 1578 2252 1584 2304
rect 1636 2252 1642 2304
rect 2222 2252 2228 2304
rect 2280 2292 2286 2304
rect 2409 2295 2467 2301
rect 2409 2292 2421 2295
rect 2280 2264 2421 2292
rect 2280 2252 2286 2264
rect 2409 2261 2421 2264
rect 2455 2261 2467 2295
rect 2409 2255 2467 2261
rect 2866 2252 2872 2304
rect 2924 2252 2930 2304
rect 3160 2301 3188 2332
rect 7650 2320 7656 2332
rect 7708 2320 7714 2372
rect 7944 2360 7972 2400
rect 8021 2397 8033 2431
rect 8067 2397 8079 2431
rect 8021 2391 8079 2397
rect 8389 2431 8447 2437
rect 8389 2397 8401 2431
rect 8435 2397 8447 2431
rect 8389 2391 8447 2397
rect 8570 2388 8576 2440
rect 8628 2388 8634 2440
rect 8956 2428 8984 2468
rect 9030 2456 9036 2508
rect 9088 2456 9094 2508
rect 9490 2456 9496 2508
rect 9548 2496 9554 2508
rect 9548 2468 10456 2496
rect 9548 2456 9554 2468
rect 10134 2428 10140 2440
rect 8956 2400 10140 2428
rect 10134 2388 10140 2400
rect 10192 2388 10198 2440
rect 10318 2388 10324 2440
rect 10376 2388 10382 2440
rect 7944 2332 8708 2360
rect 3145 2295 3203 2301
rect 3145 2261 3157 2295
rect 3191 2261 3203 2295
rect 3145 2255 3203 2261
rect 3418 2252 3424 2304
rect 3476 2292 3482 2304
rect 3881 2295 3939 2301
rect 3881 2292 3893 2295
rect 3476 2264 3893 2292
rect 3476 2252 3482 2264
rect 3881 2261 3893 2264
rect 3927 2261 3939 2295
rect 3881 2255 3939 2261
rect 4430 2252 4436 2304
rect 4488 2292 4494 2304
rect 4617 2295 4675 2301
rect 4617 2292 4629 2295
rect 4488 2264 4629 2292
rect 4488 2252 4494 2264
rect 4617 2261 4629 2264
rect 4663 2261 4675 2295
rect 4617 2255 4675 2261
rect 5534 2252 5540 2304
rect 5592 2292 5598 2304
rect 5721 2295 5779 2301
rect 5721 2292 5733 2295
rect 5592 2264 5733 2292
rect 5592 2252 5598 2264
rect 5721 2261 5733 2264
rect 5767 2261 5779 2295
rect 5721 2255 5779 2261
rect 6638 2252 6644 2304
rect 6696 2292 6702 2304
rect 6825 2295 6883 2301
rect 6825 2292 6837 2295
rect 6696 2264 6837 2292
rect 6696 2252 6702 2264
rect 6825 2261 6837 2264
rect 6871 2261 6883 2295
rect 6825 2255 6883 2261
rect 7742 2252 7748 2304
rect 7800 2292 7806 2304
rect 7837 2295 7895 2301
rect 7837 2292 7849 2295
rect 7800 2264 7849 2292
rect 7800 2252 7806 2264
rect 7837 2261 7849 2264
rect 7883 2261 7895 2295
rect 7837 2255 7895 2261
rect 8205 2295 8263 2301
rect 8205 2261 8217 2295
rect 8251 2292 8263 2295
rect 8570 2292 8576 2304
rect 8251 2264 8576 2292
rect 8251 2261 8263 2264
rect 8205 2255 8263 2261
rect 8570 2252 8576 2264
rect 8628 2252 8634 2304
rect 8680 2292 8708 2332
rect 8754 2320 8760 2372
rect 8812 2320 8818 2372
rect 9490 2360 9496 2372
rect 9232 2332 9496 2360
rect 9232 2301 9260 2332
rect 9490 2320 9496 2332
rect 9548 2320 9554 2372
rect 10428 2360 10456 2468
rect 11330 2456 11336 2508
rect 11388 2496 11394 2508
rect 12069 2499 12127 2505
rect 12069 2496 12081 2499
rect 11388 2468 12081 2496
rect 11388 2456 11394 2468
rect 12069 2465 12081 2468
rect 12115 2465 12127 2499
rect 12069 2459 12127 2465
rect 12342 2456 12348 2508
rect 12400 2496 12406 2508
rect 13170 2496 13176 2508
rect 12400 2468 13176 2496
rect 12400 2456 12406 2468
rect 10594 2388 10600 2440
rect 10652 2428 10658 2440
rect 10689 2431 10747 2437
rect 10689 2428 10701 2431
rect 10652 2400 10701 2428
rect 10652 2388 10658 2400
rect 10689 2397 10701 2400
rect 10735 2397 10747 2431
rect 10689 2391 10747 2397
rect 10778 2388 10784 2440
rect 10836 2388 10842 2440
rect 11063 2431 11121 2437
rect 11063 2398 11075 2431
rect 10888 2397 11075 2398
rect 11109 2397 11121 2431
rect 10888 2391 11121 2397
rect 10888 2370 11100 2391
rect 11882 2388 11888 2440
rect 11940 2388 11946 2440
rect 12912 2437 12940 2468
rect 13170 2456 13176 2468
rect 13228 2456 13234 2508
rect 13722 2456 13728 2508
rect 13780 2456 13786 2508
rect 12621 2431 12679 2437
rect 12621 2397 12633 2431
rect 12667 2397 12679 2431
rect 12621 2391 12679 2397
rect 12897 2431 12955 2437
rect 12897 2397 12909 2431
rect 12943 2397 12955 2431
rect 12897 2391 12955 2397
rect 13541 2431 13599 2437
rect 13541 2397 13553 2431
rect 13587 2428 13599 2431
rect 14016 2428 14044 2536
rect 17034 2524 17040 2536
rect 17092 2524 17098 2576
rect 20165 2567 20223 2573
rect 20165 2533 20177 2567
rect 20211 2564 20223 2567
rect 27080 2564 27108 2604
rect 29454 2592 29460 2604
rect 29512 2592 29518 2644
rect 30837 2635 30895 2641
rect 30837 2601 30849 2635
rect 30883 2632 30895 2635
rect 30926 2632 30932 2644
rect 30883 2604 30932 2632
rect 30883 2601 30895 2604
rect 30837 2595 30895 2601
rect 30926 2592 30932 2604
rect 30984 2592 30990 2644
rect 31386 2592 31392 2644
rect 31444 2632 31450 2644
rect 31444 2604 31616 2632
rect 31444 2592 31450 2604
rect 20211 2536 27108 2564
rect 20211 2533 20223 2536
rect 20165 2527 20223 2533
rect 30374 2524 30380 2576
rect 30432 2564 30438 2576
rect 31478 2564 31484 2576
rect 30432 2536 31484 2564
rect 30432 2524 30438 2536
rect 15010 2456 15016 2508
rect 15068 2496 15074 2508
rect 15197 2499 15255 2505
rect 15197 2496 15209 2499
rect 15068 2468 15209 2496
rect 15068 2456 15074 2468
rect 15197 2465 15209 2468
rect 15243 2465 15255 2499
rect 15197 2459 15255 2465
rect 15289 2499 15347 2505
rect 15289 2465 15301 2499
rect 15335 2496 15347 2499
rect 15562 2496 15568 2508
rect 15335 2468 15568 2496
rect 15335 2465 15347 2468
rect 15289 2459 15347 2465
rect 15562 2456 15568 2468
rect 15620 2496 15626 2508
rect 18322 2496 18328 2508
rect 15620 2468 18328 2496
rect 15620 2456 15626 2468
rect 13587 2400 14044 2428
rect 14093 2431 14151 2437
rect 13587 2397 13599 2400
rect 13541 2391 13599 2397
rect 14093 2397 14105 2431
rect 14139 2428 14151 2431
rect 14550 2428 14556 2440
rect 14139 2400 14556 2428
rect 14139 2397 14151 2400
rect 14093 2391 14151 2397
rect 10888 2360 10916 2370
rect 10428 2332 10916 2360
rect 11974 2320 11980 2372
rect 12032 2320 12038 2372
rect 12066 2320 12072 2372
rect 12124 2360 12130 2372
rect 12636 2360 12664 2391
rect 14550 2388 14556 2400
rect 14608 2388 14614 2440
rect 14734 2388 14740 2440
rect 14792 2388 14798 2440
rect 15838 2428 15844 2440
rect 14844 2400 15844 2428
rect 13633 2363 13691 2369
rect 13633 2360 13645 2363
rect 12124 2332 13645 2360
rect 12124 2320 12130 2332
rect 13633 2329 13645 2332
rect 13679 2360 13691 2363
rect 14844 2360 14872 2400
rect 15838 2388 15844 2400
rect 15896 2388 15902 2440
rect 15930 2388 15936 2440
rect 15988 2428 15994 2440
rect 16960 2437 16988 2468
rect 18322 2456 18328 2468
rect 18380 2456 18386 2508
rect 18966 2456 18972 2508
rect 19024 2456 19030 2508
rect 20993 2499 21051 2505
rect 20993 2465 21005 2499
rect 21039 2496 21051 2499
rect 21450 2496 21456 2508
rect 21039 2468 21456 2496
rect 21039 2465 21051 2468
rect 20993 2459 21051 2465
rect 21450 2456 21456 2468
rect 21508 2456 21514 2508
rect 21634 2456 21640 2508
rect 21692 2496 21698 2508
rect 21692 2468 26832 2496
rect 21692 2456 21698 2468
rect 16117 2431 16175 2437
rect 16117 2428 16129 2431
rect 15988 2400 16129 2428
rect 15988 2388 15994 2400
rect 16117 2397 16129 2400
rect 16163 2397 16175 2431
rect 16117 2391 16175 2397
rect 16945 2431 17003 2437
rect 16945 2397 16957 2431
rect 16991 2397 17003 2431
rect 16945 2391 17003 2397
rect 17494 2388 17500 2440
rect 17552 2428 17558 2440
rect 17681 2431 17739 2437
rect 17681 2428 17693 2431
rect 17552 2400 17693 2428
rect 17552 2388 17558 2400
rect 17681 2397 17693 2400
rect 17727 2397 17739 2431
rect 17681 2391 17739 2397
rect 18690 2388 18696 2440
rect 18748 2388 18754 2440
rect 19426 2388 19432 2440
rect 19484 2388 19490 2440
rect 19886 2388 19892 2440
rect 19944 2428 19950 2440
rect 19981 2431 20039 2437
rect 19981 2428 19993 2431
rect 19944 2400 19993 2428
rect 19944 2388 19950 2400
rect 19981 2397 19993 2400
rect 20027 2397 20039 2431
rect 19981 2391 20039 2397
rect 20898 2388 20904 2440
rect 20956 2428 20962 2440
rect 21821 2431 21879 2437
rect 21821 2428 21833 2431
rect 20956 2400 21833 2428
rect 20956 2388 20962 2400
rect 21821 2397 21833 2400
rect 21867 2397 21879 2431
rect 21821 2391 21879 2397
rect 23109 2431 23167 2437
rect 23109 2397 23121 2431
rect 23155 2428 23167 2431
rect 23198 2428 23204 2440
rect 23155 2400 23204 2428
rect 23155 2397 23167 2400
rect 23109 2391 23167 2397
rect 23198 2388 23204 2400
rect 23256 2388 23262 2440
rect 25884 2400 26188 2428
rect 13679 2332 14872 2360
rect 15381 2363 15439 2369
rect 13679 2329 13691 2332
rect 13633 2323 13691 2329
rect 15381 2329 15393 2363
rect 15427 2360 15439 2363
rect 25884 2360 25912 2400
rect 15427 2332 25912 2360
rect 15427 2329 15439 2332
rect 15381 2323 15439 2329
rect 9217 2295 9275 2301
rect 9217 2292 9229 2295
rect 8680 2264 9229 2292
rect 9217 2261 9229 2264
rect 9263 2261 9275 2295
rect 9217 2255 9275 2261
rect 9309 2295 9367 2301
rect 9309 2261 9321 2295
rect 9355 2292 9367 2295
rect 9582 2292 9588 2304
rect 9355 2264 9588 2292
rect 9355 2261 9367 2264
rect 9309 2255 9367 2261
rect 9582 2252 9588 2264
rect 9640 2252 9646 2304
rect 9677 2295 9735 2301
rect 9677 2261 9689 2295
rect 9723 2292 9735 2295
rect 9766 2292 9772 2304
rect 9723 2264 9772 2292
rect 9723 2261 9735 2264
rect 9677 2255 9735 2261
rect 9766 2252 9772 2264
rect 9824 2252 9830 2304
rect 9950 2252 9956 2304
rect 10008 2292 10014 2304
rect 10137 2295 10195 2301
rect 10137 2292 10149 2295
rect 10008 2264 10149 2292
rect 10008 2252 10014 2264
rect 10137 2261 10149 2264
rect 10183 2261 10195 2295
rect 10137 2255 10195 2261
rect 11054 2252 11060 2304
rect 11112 2292 11118 2304
rect 11241 2295 11299 2301
rect 11241 2292 11253 2295
rect 11112 2264 11253 2292
rect 11112 2252 11118 2264
rect 11241 2261 11253 2264
rect 11287 2261 11299 2295
rect 11241 2255 11299 2261
rect 11698 2252 11704 2304
rect 11756 2292 11762 2304
rect 12342 2292 12348 2304
rect 11756 2264 12348 2292
rect 11756 2252 11762 2264
rect 12342 2252 12348 2264
rect 12400 2252 12406 2304
rect 12434 2252 12440 2304
rect 12492 2252 12498 2304
rect 13078 2252 13084 2304
rect 13136 2252 13142 2304
rect 14277 2295 14335 2301
rect 14277 2261 14289 2295
rect 14323 2292 14335 2295
rect 14366 2292 14372 2304
rect 14323 2264 14372 2292
rect 14323 2261 14335 2264
rect 14277 2255 14335 2261
rect 14366 2252 14372 2264
rect 14424 2252 14430 2304
rect 15470 2252 15476 2304
rect 15528 2292 15534 2304
rect 15933 2295 15991 2301
rect 15933 2292 15945 2295
rect 15528 2264 15945 2292
rect 15528 2252 15534 2264
rect 15933 2261 15945 2264
rect 15979 2261 15991 2295
rect 15933 2255 15991 2261
rect 16574 2252 16580 2304
rect 16632 2292 16638 2304
rect 16761 2295 16819 2301
rect 16761 2292 16773 2295
rect 16632 2264 16773 2292
rect 16632 2252 16638 2264
rect 16761 2261 16773 2264
rect 16807 2261 16819 2295
rect 16761 2255 16819 2261
rect 17494 2252 17500 2304
rect 17552 2252 17558 2304
rect 19242 2252 19248 2304
rect 19300 2252 19306 2304
rect 20806 2252 20812 2304
rect 20864 2292 20870 2304
rect 21082 2292 21088 2304
rect 20864 2264 21088 2292
rect 20864 2252 20870 2264
rect 21082 2252 21088 2264
rect 21140 2252 21146 2304
rect 21177 2295 21235 2301
rect 21177 2261 21189 2295
rect 21223 2292 21235 2295
rect 21542 2292 21548 2304
rect 21223 2264 21548 2292
rect 21223 2261 21235 2264
rect 21177 2255 21235 2261
rect 21542 2252 21548 2264
rect 21600 2252 21606 2304
rect 22005 2295 22063 2301
rect 22005 2261 22017 2295
rect 22051 2292 22063 2295
rect 25866 2292 25872 2304
rect 22051 2264 25872 2292
rect 22051 2261 22063 2264
rect 22005 2255 22063 2261
rect 25866 2252 25872 2264
rect 25924 2252 25930 2304
rect 26160 2292 26188 2400
rect 26804 2360 26832 2468
rect 26878 2456 26884 2508
rect 26936 2496 26942 2508
rect 27433 2499 27491 2505
rect 27433 2496 27445 2499
rect 26936 2468 27445 2496
rect 26936 2456 26942 2468
rect 27433 2465 27445 2468
rect 27479 2465 27491 2499
rect 27433 2459 27491 2465
rect 27522 2456 27528 2508
rect 27580 2456 27586 2508
rect 27341 2431 27399 2437
rect 27341 2397 27353 2431
rect 27387 2428 27399 2431
rect 27798 2428 27804 2440
rect 27387 2400 27804 2428
rect 27387 2397 27399 2400
rect 27341 2391 27399 2397
rect 27798 2388 27804 2400
rect 27856 2388 27862 2440
rect 30668 2437 30696 2536
rect 31478 2524 31484 2536
rect 31536 2524 31542 2576
rect 31588 2564 31616 2604
rect 32306 2592 32312 2644
rect 32364 2632 32370 2644
rect 32493 2635 32551 2641
rect 32493 2632 32505 2635
rect 32364 2604 32505 2632
rect 32364 2592 32370 2604
rect 32493 2601 32505 2604
rect 32539 2601 32551 2635
rect 32493 2595 32551 2601
rect 33689 2635 33747 2641
rect 33689 2601 33701 2635
rect 33735 2632 33747 2635
rect 38286 2632 38292 2644
rect 33735 2604 38292 2632
rect 33735 2601 33747 2604
rect 33689 2595 33747 2601
rect 38286 2592 38292 2604
rect 38344 2592 38350 2644
rect 31588 2536 38516 2564
rect 31570 2456 31576 2508
rect 31628 2496 31634 2508
rect 31628 2468 32996 2496
rect 31628 2456 31634 2468
rect 30653 2431 30711 2437
rect 30653 2397 30665 2431
rect 30699 2397 30711 2431
rect 30653 2391 30711 2397
rect 31662 2388 31668 2440
rect 31720 2428 31726 2440
rect 31757 2431 31815 2437
rect 31757 2428 31769 2431
rect 31720 2400 31769 2428
rect 31720 2388 31726 2400
rect 31757 2397 31769 2400
rect 31803 2397 31815 2431
rect 32674 2428 32680 2440
rect 31757 2391 31815 2397
rect 31864 2400 32680 2428
rect 31386 2360 31392 2372
rect 26804 2332 31392 2360
rect 31386 2320 31392 2332
rect 31444 2320 31450 2372
rect 31864 2292 31892 2400
rect 32674 2388 32680 2400
rect 32732 2388 32738 2440
rect 32766 2388 32772 2440
rect 32824 2428 32830 2440
rect 32861 2431 32919 2437
rect 32861 2428 32873 2431
rect 32824 2400 32873 2428
rect 32824 2388 32830 2400
rect 32861 2397 32873 2400
rect 32907 2397 32919 2431
rect 32968 2428 32996 2468
rect 33042 2456 33048 2508
rect 33100 2456 33106 2508
rect 37826 2496 37832 2508
rect 33888 2468 37832 2496
rect 33505 2431 33563 2437
rect 33505 2428 33517 2431
rect 32968 2400 33517 2428
rect 32861 2391 32919 2397
rect 33505 2397 33517 2400
rect 33551 2428 33563 2431
rect 33686 2428 33692 2440
rect 33551 2400 33692 2428
rect 33551 2397 33563 2400
rect 33505 2391 33563 2397
rect 33686 2388 33692 2400
rect 33744 2388 33750 2440
rect 33888 2360 33916 2468
rect 37826 2456 37832 2468
rect 37884 2456 37890 2508
rect 34333 2431 34391 2437
rect 34333 2397 34345 2431
rect 34379 2428 34391 2431
rect 34514 2428 34520 2440
rect 34379 2400 34520 2428
rect 34379 2397 34391 2400
rect 34333 2391 34391 2397
rect 34514 2388 34520 2400
rect 34572 2388 34578 2440
rect 34606 2388 34612 2440
rect 34664 2428 34670 2440
rect 37737 2431 37795 2437
rect 37737 2428 37749 2431
rect 34664 2400 37749 2428
rect 34664 2388 34670 2400
rect 37737 2397 37749 2400
rect 37783 2397 37795 2431
rect 37737 2391 37795 2397
rect 38102 2388 38108 2440
rect 38160 2388 38166 2440
rect 38488 2437 38516 2536
rect 39390 2524 39396 2576
rect 39448 2524 39454 2576
rect 38473 2431 38531 2437
rect 38473 2397 38485 2431
rect 38519 2397 38531 2431
rect 38473 2391 38531 2397
rect 38838 2388 38844 2440
rect 38896 2388 38902 2440
rect 39209 2431 39267 2437
rect 39209 2397 39221 2431
rect 39255 2397 39267 2431
rect 39209 2391 39267 2397
rect 31956 2332 33916 2360
rect 31956 2301 31984 2332
rect 37458 2320 37464 2372
rect 37516 2360 37522 2372
rect 39224 2360 39252 2391
rect 37516 2332 39252 2360
rect 37516 2320 37522 2332
rect 26160 2264 31892 2292
rect 31941 2295 31999 2301
rect 31941 2261 31953 2295
rect 31987 2261 31999 2295
rect 31941 2255 31999 2261
rect 32858 2252 32864 2304
rect 32916 2292 32922 2304
rect 32953 2295 33011 2301
rect 32953 2292 32965 2295
rect 32916 2264 32965 2292
rect 32916 2252 32922 2264
rect 32953 2261 32965 2264
rect 32999 2261 33011 2295
rect 32953 2255 33011 2261
rect 33410 2252 33416 2304
rect 33468 2292 33474 2304
rect 34241 2295 34299 2301
rect 34241 2292 34253 2295
rect 33468 2264 34253 2292
rect 33468 2252 33474 2264
rect 34241 2261 34253 2264
rect 34287 2261 34299 2295
rect 34241 2255 34299 2261
rect 37918 2252 37924 2304
rect 37976 2252 37982 2304
rect 38286 2252 38292 2304
rect 38344 2252 38350 2304
rect 38657 2295 38715 2301
rect 38657 2261 38669 2295
rect 38703 2292 38715 2295
rect 38930 2292 38936 2304
rect 38703 2264 38936 2292
rect 38703 2261 38715 2264
rect 38657 2255 38715 2261
rect 38930 2252 38936 2264
rect 38988 2252 38994 2304
rect 39025 2295 39083 2301
rect 39025 2261 39037 2295
rect 39071 2292 39083 2295
rect 39942 2292 39948 2304
rect 39071 2264 39948 2292
rect 39071 2261 39083 2264
rect 39025 2255 39083 2261
rect 39942 2252 39948 2264
rect 40000 2252 40006 2304
rect 1104 2202 39836 2224
rect 1104 2150 3010 2202
rect 3062 2150 3074 2202
rect 3126 2150 3138 2202
rect 3190 2150 3202 2202
rect 3254 2150 3266 2202
rect 3318 2150 9010 2202
rect 9062 2150 9074 2202
rect 9126 2150 9138 2202
rect 9190 2150 9202 2202
rect 9254 2150 9266 2202
rect 9318 2150 15010 2202
rect 15062 2150 15074 2202
rect 15126 2150 15138 2202
rect 15190 2150 15202 2202
rect 15254 2150 15266 2202
rect 15318 2150 21010 2202
rect 21062 2150 21074 2202
rect 21126 2150 21138 2202
rect 21190 2150 21202 2202
rect 21254 2150 21266 2202
rect 21318 2150 27010 2202
rect 27062 2150 27074 2202
rect 27126 2150 27138 2202
rect 27190 2150 27202 2202
rect 27254 2150 27266 2202
rect 27318 2150 33010 2202
rect 33062 2150 33074 2202
rect 33126 2150 33138 2202
rect 33190 2150 33202 2202
rect 33254 2150 33266 2202
rect 33318 2150 39010 2202
rect 39062 2150 39074 2202
rect 39126 2150 39138 2202
rect 39190 2150 39202 2202
rect 39254 2150 39266 2202
rect 39318 2150 39836 2202
rect 1104 2128 39836 2150
rect 1578 2048 1584 2100
rect 1636 2088 1642 2100
rect 7558 2088 7564 2100
rect 1636 2060 7564 2088
rect 1636 2048 1642 2060
rect 7558 2048 7564 2060
rect 7616 2048 7622 2100
rect 9490 2048 9496 2100
rect 9548 2088 9554 2100
rect 10686 2088 10692 2100
rect 9548 2060 10692 2088
rect 9548 2048 9554 2060
rect 10686 2048 10692 2060
rect 10744 2088 10750 2100
rect 12066 2088 12072 2100
rect 10744 2060 12072 2088
rect 10744 2048 10750 2060
rect 12066 2048 12072 2060
rect 12124 2048 12130 2100
rect 12158 2048 12164 2100
rect 12216 2088 12222 2100
rect 17862 2088 17868 2100
rect 12216 2060 17868 2088
rect 12216 2048 12222 2060
rect 17862 2048 17868 2060
rect 17920 2048 17926 2100
rect 18322 2048 18328 2100
rect 18380 2088 18386 2100
rect 26786 2088 26792 2100
rect 18380 2060 26792 2088
rect 18380 2048 18386 2060
rect 26786 2048 26792 2060
rect 26844 2048 26850 2100
rect 27706 2048 27712 2100
rect 27764 2088 27770 2100
rect 37458 2088 37464 2100
rect 27764 2060 37464 2088
rect 27764 2048 27770 2060
rect 37458 2048 37464 2060
rect 37516 2048 37522 2100
rect 2866 1980 2872 2032
rect 2924 2020 2930 2032
rect 11698 2020 11704 2032
rect 2924 1992 11704 2020
rect 2924 1980 2930 1992
rect 11698 1980 11704 1992
rect 11756 1980 11762 2032
rect 15746 2020 15752 2032
rect 11808 1992 15752 2020
rect 3786 1912 3792 1964
rect 3844 1952 3850 1964
rect 11808 1952 11836 1992
rect 15746 1980 15752 1992
rect 15804 1980 15810 2032
rect 26878 1980 26884 2032
rect 26936 2020 26942 2032
rect 34606 2020 34612 2032
rect 26936 1992 34612 2020
rect 26936 1980 26942 1992
rect 34606 1980 34612 1992
rect 34664 1980 34670 2032
rect 3844 1924 11836 1952
rect 3844 1912 3850 1924
rect 11974 1912 11980 1964
rect 12032 1952 12038 1964
rect 12032 1924 19334 1952
rect 12032 1912 12038 1924
rect 5902 1844 5908 1896
rect 5960 1884 5966 1896
rect 13814 1884 13820 1896
rect 5960 1856 13820 1884
rect 5960 1844 5966 1856
rect 13814 1844 13820 1856
rect 13872 1844 13878 1896
rect 19306 1884 19334 1924
rect 20438 1912 20444 1964
rect 20496 1952 20502 1964
rect 32582 1952 32588 1964
rect 20496 1924 32588 1952
rect 20496 1912 20502 1924
rect 32582 1912 32588 1924
rect 32640 1912 32646 1964
rect 20806 1884 20812 1896
rect 19306 1856 20812 1884
rect 20806 1844 20812 1856
rect 20864 1844 20870 1896
rect 28074 1844 28080 1896
rect 28132 1884 28138 1896
rect 38102 1884 38108 1896
rect 28132 1856 38108 1884
rect 28132 1844 28138 1856
rect 38102 1844 38108 1856
rect 38160 1844 38166 1896
rect 4798 1776 4804 1828
rect 4856 1816 4862 1828
rect 16298 1816 16304 1828
rect 4856 1788 16304 1816
rect 4856 1776 4862 1788
rect 16298 1776 16304 1788
rect 16356 1776 16362 1828
rect 17126 1776 17132 1828
rect 17184 1816 17190 1828
rect 36906 1816 36912 1828
rect 17184 1788 36912 1816
rect 17184 1776 17190 1788
rect 36906 1776 36912 1788
rect 36964 1776 36970 1828
rect 11146 1708 11152 1760
rect 11204 1748 11210 1760
rect 33410 1748 33416 1760
rect 11204 1720 33416 1748
rect 11204 1708 11210 1720
rect 33410 1708 33416 1720
rect 33468 1708 33474 1760
rect 10134 1640 10140 1692
rect 10192 1680 10198 1692
rect 11238 1680 11244 1692
rect 10192 1652 11244 1680
rect 10192 1640 10198 1652
rect 11238 1640 11244 1652
rect 11296 1680 11302 1692
rect 11974 1680 11980 1692
rect 11296 1652 11980 1680
rect 11296 1640 11302 1652
rect 11974 1640 11980 1652
rect 12032 1640 12038 1692
rect 12526 1640 12532 1692
rect 12584 1680 12590 1692
rect 31570 1680 31576 1692
rect 12584 1652 31576 1680
rect 12584 1640 12590 1652
rect 31570 1640 31576 1652
rect 31628 1640 31634 1692
rect 1762 1572 1768 1624
rect 1820 1612 1826 1624
rect 17954 1612 17960 1624
rect 1820 1584 17960 1612
rect 1820 1572 1826 1584
rect 17954 1572 17960 1584
rect 18012 1572 18018 1624
rect 25866 1572 25872 1624
rect 25924 1612 25930 1624
rect 30006 1612 30012 1624
rect 25924 1584 30012 1612
rect 25924 1572 25930 1584
rect 30006 1572 30012 1584
rect 30064 1572 30070 1624
rect 7650 1504 7656 1556
rect 7708 1544 7714 1556
rect 12802 1544 12808 1556
rect 7708 1516 12808 1544
rect 7708 1504 7714 1516
rect 12802 1504 12808 1516
rect 12860 1504 12866 1556
rect 11146 1436 11152 1488
rect 11204 1476 11210 1488
rect 32490 1476 32496 1488
rect 11204 1448 32496 1476
rect 11204 1436 11210 1448
rect 32490 1436 32496 1448
rect 32548 1436 32554 1488
rect 6730 1300 6736 1352
rect 6788 1340 6794 1352
rect 35066 1340 35072 1352
rect 6788 1312 35072 1340
rect 6788 1300 6794 1312
rect 35066 1300 35072 1312
rect 35124 1300 35130 1352
rect 10962 1232 10968 1284
rect 11020 1272 11026 1284
rect 39574 1272 39580 1284
rect 11020 1244 39580 1272
rect 11020 1232 11026 1244
rect 39574 1232 39580 1244
rect 39632 1232 39638 1284
rect 13078 1164 13084 1216
rect 13136 1204 13142 1216
rect 38838 1204 38844 1216
rect 13136 1176 38844 1204
rect 13136 1164 13142 1176
rect 38838 1164 38844 1176
rect 38896 1164 38902 1216
rect 7558 1096 7564 1148
rect 7616 1136 7622 1148
rect 17310 1136 17316 1148
rect 7616 1108 17316 1136
rect 7616 1096 7622 1108
rect 17310 1096 17316 1108
rect 17368 1096 17374 1148
rect 3510 1028 3516 1080
rect 3568 1068 3574 1080
rect 28166 1068 28172 1080
rect 3568 1040 28172 1068
rect 3568 1028 3574 1040
rect 28166 1028 28172 1040
rect 28224 1028 28230 1080
rect 10226 960 10232 1012
rect 10284 1000 10290 1012
rect 33870 1000 33876 1012
rect 10284 972 33876 1000
rect 10284 960 10290 972
rect 33870 960 33876 972
rect 33928 960 33934 1012
rect 8754 892 8760 944
rect 8812 932 8818 944
rect 29822 932 29828 944
rect 8812 904 29828 932
rect 8812 892 8818 904
rect 29822 892 29828 904
rect 29880 892 29886 944
rect 7374 824 7380 876
rect 7432 864 7438 876
rect 23474 864 23480 876
rect 7432 836 23480 864
rect 7432 824 7438 836
rect 23474 824 23480 836
rect 23532 824 23538 876
rect 4522 756 4528 808
rect 4580 796 4586 808
rect 18414 796 18420 808
rect 4580 768 18420 796
rect 4580 756 4586 768
rect 18414 756 18420 768
rect 18472 756 18478 808
rect 7466 688 7472 740
rect 7524 728 7530 740
rect 27522 728 27528 740
rect 7524 700 27528 728
rect 7524 688 7530 700
rect 27522 688 27528 700
rect 27580 688 27586 740
rect 1486 620 1492 672
rect 1544 660 1550 672
rect 18046 660 18052 672
rect 1544 632 18052 660
rect 1544 620 1550 632
rect 18046 620 18052 632
rect 18104 620 18110 672
rect 7282 552 7288 604
rect 7340 592 7346 604
rect 23934 592 23940 604
rect 7340 564 23940 592
rect 7340 552 7346 564
rect 23934 552 23940 564
rect 23992 552 23998 604
rect 4706 484 4712 536
rect 4764 524 4770 536
rect 29546 524 29552 536
rect 4764 496 29552 524
rect 4764 484 4770 496
rect 29546 484 29552 496
rect 29604 484 29610 536
rect 2498 416 2504 468
rect 2556 456 2562 468
rect 16942 456 16948 468
rect 2556 428 16948 456
rect 2556 416 2562 428
rect 16942 416 16948 428
rect 17000 416 17006 468
rect 23198 144 23204 196
rect 23256 144 23262 196
rect 24302 144 24308 196
rect 24360 184 24366 196
rect 38562 184 38568 196
rect 24360 156 38568 184
rect 24360 144 24366 156
rect 38562 144 38568 156
rect 38620 144 38626 196
rect 23216 116 23244 144
rect 37734 116 37740 128
rect 23216 88 37740 116
rect 37734 76 37740 88
rect 37792 76 37798 128
rect 22186 8 22192 60
rect 22244 48 22250 60
rect 39482 48 39488 60
rect 22244 20 39488 48
rect 22244 8 22250 20
rect 39482 8 39488 20
rect 39540 8 39546 60
<< via1 >>
rect 6644 11160 6696 11212
rect 12900 11160 12952 11212
rect 17224 10820 17276 10872
rect 18420 10820 18472 10872
rect 12992 10684 13044 10736
rect 14556 10684 14608 10736
rect 12900 10480 12952 10532
rect 20996 10480 21048 10532
rect 1492 10412 1544 10464
rect 3516 10412 3568 10464
rect 2044 10208 2096 10260
rect 23020 10412 23072 10464
rect 7288 10344 7340 10396
rect 22376 10344 22428 10396
rect 8944 10276 8996 10328
rect 17132 10276 17184 10328
rect 28908 10276 28960 10328
rect 32404 10276 32456 10328
rect 9496 10208 9548 10260
rect 17500 10208 17552 10260
rect 6460 10140 6512 10192
rect 8760 10140 8812 10192
rect 12808 10140 12860 10192
rect 19064 10140 19116 10192
rect 23572 10140 23624 10192
rect 30472 10140 30524 10192
rect 7012 10072 7064 10124
rect 7840 10004 7892 10056
rect 9588 10004 9640 10056
rect 10232 10072 10284 10124
rect 3700 9936 3752 9988
rect 6552 9936 6604 9988
rect 8392 9936 8444 9988
rect 13728 9936 13780 9988
rect 6092 9868 6144 9920
rect 11796 9868 11848 9920
rect 11888 9868 11940 9920
rect 12624 9868 12676 9920
rect 19156 10072 19208 10124
rect 20904 10072 20956 10124
rect 20996 10072 21048 10124
rect 30748 10072 30800 10124
rect 17500 10004 17552 10056
rect 26608 10004 26660 10056
rect 27988 9936 28040 9988
rect 26792 9868 26844 9920
rect 6184 9800 6236 9852
rect 7932 9800 7984 9852
rect 9588 9800 9640 9852
rect 14004 9800 14056 9852
rect 16948 9800 17000 9852
rect 18972 9800 19024 9852
rect 19064 9800 19116 9852
rect 23572 9800 23624 9852
rect 24124 9800 24176 9852
rect 35624 9868 35676 9920
rect 1768 9732 1820 9784
rect 4344 9732 4396 9784
rect 8576 9732 8628 9784
rect 12348 9732 12400 9784
rect 3424 9664 3476 9716
rect 4620 9664 4672 9716
rect 7196 9664 7248 9716
rect 12072 9664 12124 9716
rect 6368 9596 6420 9648
rect 8944 9596 8996 9648
rect 9036 9596 9088 9648
rect 17132 9664 17184 9716
rect 24124 9664 24176 9716
rect 33784 9732 33836 9784
rect 27804 9664 27856 9716
rect 32312 9664 32364 9716
rect 5908 9528 5960 9580
rect 11796 9528 11848 9580
rect 1676 9460 1728 9512
rect 9772 9460 9824 9512
rect 9864 9460 9916 9512
rect 17132 9460 17184 9512
rect 17500 9460 17552 9512
rect 24400 9460 24452 9512
rect 10784 9392 10836 9444
rect 4252 9324 4304 9376
rect 10324 9324 10376 9376
rect 10508 9324 10560 9376
rect 17960 9392 18012 9444
rect 23664 9392 23716 9444
rect 26424 9392 26476 9444
rect 27344 9392 27396 9444
rect 29552 9460 29604 9512
rect 29000 9392 29052 9444
rect 34244 9392 34296 9444
rect 2136 9188 2188 9240
rect 5632 9256 5684 9308
rect 16304 9256 16356 9308
rect 16856 9256 16908 9308
rect 22744 9324 22796 9376
rect 29828 9324 29880 9376
rect 30012 9324 30064 9376
rect 31300 9324 31352 9376
rect 31392 9324 31444 9376
rect 32588 9324 32640 9376
rect 18604 9256 18656 9308
rect 22836 9256 22888 9308
rect 23664 9256 23716 9308
rect 25412 9256 25464 9308
rect 38568 9256 38620 9308
rect 5540 9188 5592 9240
rect 11704 9188 11756 9240
rect 11796 9188 11848 9240
rect 1860 9120 1912 9172
rect 9680 9120 9732 9172
rect 11336 9120 11388 9172
rect 18052 9120 18104 9172
rect 26148 9188 26200 9240
rect 28816 9188 28868 9240
rect 29736 9188 29788 9240
rect 31576 9188 31628 9240
rect 31944 9188 31996 9240
rect 33968 9188 34020 9240
rect 26332 9120 26384 9172
rect 27804 9120 27856 9172
rect 30932 9120 30984 9172
rect 5448 9052 5500 9104
rect 16856 9052 16908 9104
rect 23848 9052 23900 9104
rect 3608 8984 3660 9036
rect 6000 8984 6052 9036
rect 8024 8984 8076 9036
rect 12072 8984 12124 9036
rect 13084 8984 13136 9036
rect 20536 8984 20588 9036
rect 1400 8916 1452 8968
rect 6920 8916 6972 8968
rect 7748 8916 7800 8968
rect 1584 8848 1636 8900
rect 8116 8848 8168 8900
rect 8852 8916 8904 8968
rect 13084 8848 13136 8900
rect 13268 8848 13320 8900
rect 15200 8848 15252 8900
rect 3884 8780 3936 8832
rect 9036 8780 9088 8832
rect 11796 8780 11848 8832
rect 14740 8780 14792 8832
rect 16028 8780 16080 8832
rect 16488 8780 16540 8832
rect 18236 8916 18288 8968
rect 24032 8916 24084 8968
rect 18972 8848 19024 8900
rect 27896 9052 27948 9104
rect 29368 9052 29420 9104
rect 34980 9052 35032 9104
rect 24308 8984 24360 9036
rect 30104 8984 30156 9036
rect 32220 8984 32272 9036
rect 34796 8984 34848 9036
rect 26516 8916 26568 8968
rect 31760 8916 31812 8968
rect 33048 8916 33100 8968
rect 34520 8916 34572 8968
rect 35348 8916 35400 8968
rect 38384 8916 38436 8968
rect 25596 8848 25648 8900
rect 26884 8848 26936 8900
rect 27528 8848 27580 8900
rect 32128 8848 32180 8900
rect 34336 8848 34388 8900
rect 36544 8848 36596 8900
rect 21548 8780 21600 8832
rect 22836 8780 22888 8832
rect 23848 8780 23900 8832
rect 25320 8780 25372 8832
rect 30196 8780 30248 8832
rect 33324 8780 33376 8832
rect 33784 8780 33836 8832
rect 35716 8780 35768 8832
rect 37372 8780 37424 8832
rect 3010 8678 3062 8730
rect 3074 8678 3126 8730
rect 3138 8678 3190 8730
rect 3202 8678 3254 8730
rect 3266 8678 3318 8730
rect 9010 8678 9062 8730
rect 9074 8678 9126 8730
rect 9138 8678 9190 8730
rect 9202 8678 9254 8730
rect 9266 8678 9318 8730
rect 15010 8678 15062 8730
rect 15074 8678 15126 8730
rect 15138 8678 15190 8730
rect 15202 8678 15254 8730
rect 15266 8678 15318 8730
rect 21010 8678 21062 8730
rect 21074 8678 21126 8730
rect 21138 8678 21190 8730
rect 21202 8678 21254 8730
rect 21266 8678 21318 8730
rect 27010 8678 27062 8730
rect 27074 8678 27126 8730
rect 27138 8678 27190 8730
rect 27202 8678 27254 8730
rect 27266 8678 27318 8730
rect 33010 8678 33062 8730
rect 33074 8678 33126 8730
rect 33138 8678 33190 8730
rect 33202 8678 33254 8730
rect 33266 8678 33318 8730
rect 39010 8678 39062 8730
rect 39074 8678 39126 8730
rect 39138 8678 39190 8730
rect 39202 8678 39254 8730
rect 39266 8678 39318 8730
rect 1584 8619 1636 8628
rect 1584 8585 1593 8619
rect 1593 8585 1627 8619
rect 1627 8585 1636 8619
rect 1584 8576 1636 8585
rect 3516 8619 3568 8628
rect 3516 8585 3525 8619
rect 3525 8585 3559 8619
rect 3559 8585 3568 8619
rect 3516 8576 3568 8585
rect 4436 8619 4488 8628
rect 4436 8585 4445 8619
rect 4445 8585 4479 8619
rect 4479 8585 4488 8619
rect 4436 8576 4488 8585
rect 5448 8619 5500 8628
rect 5448 8585 5457 8619
rect 5457 8585 5491 8619
rect 5491 8585 5500 8619
rect 5448 8576 5500 8585
rect 5816 8576 5868 8628
rect 6092 8619 6144 8628
rect 6092 8585 6101 8619
rect 6101 8585 6135 8619
rect 6135 8585 6144 8619
rect 6092 8576 6144 8585
rect 6644 8576 6696 8628
rect 7012 8576 7064 8628
rect 7196 8576 7248 8628
rect 7748 8576 7800 8628
rect 8392 8576 8444 8628
rect 8576 8619 8628 8628
rect 8576 8585 8585 8619
rect 8585 8585 8619 8619
rect 8619 8585 8628 8619
rect 8576 8576 8628 8585
rect 9588 8576 9640 8628
rect 1400 8483 1452 8492
rect 1400 8449 1409 8483
rect 1409 8449 1443 8483
rect 1443 8449 1452 8483
rect 1400 8440 1452 8449
rect 1676 8483 1728 8492
rect 1676 8449 1685 8483
rect 1685 8449 1719 8483
rect 1719 8449 1728 8483
rect 1676 8440 1728 8449
rect 1860 8483 1912 8492
rect 1860 8449 1869 8483
rect 1869 8449 1903 8483
rect 1903 8449 1912 8483
rect 1860 8440 1912 8449
rect 3976 8508 4028 8560
rect 2136 8483 2188 8492
rect 2136 8449 2145 8483
rect 2145 8449 2179 8483
rect 2179 8449 2188 8483
rect 2136 8440 2188 8449
rect 2504 8483 2556 8492
rect 2504 8449 2513 8483
rect 2513 8449 2547 8483
rect 2547 8449 2556 8483
rect 2504 8440 2556 8449
rect 3884 8440 3936 8492
rect 1124 8372 1176 8424
rect 9496 8508 9548 8560
rect 11244 8576 11296 8628
rect 11612 8576 11664 8628
rect 11796 8619 11848 8628
rect 11796 8585 11805 8619
rect 11805 8585 11839 8619
rect 11839 8585 11848 8619
rect 11796 8576 11848 8585
rect 12992 8576 13044 8628
rect 14924 8576 14976 8628
rect 12072 8508 12124 8560
rect 4804 8440 4856 8492
rect 6000 8440 6052 8492
rect 7656 8483 7708 8492
rect 7656 8449 7665 8483
rect 7665 8449 7699 8483
rect 7699 8449 7708 8483
rect 7656 8440 7708 8449
rect 8116 8483 8168 8492
rect 8116 8449 8125 8483
rect 8125 8449 8159 8483
rect 8159 8449 8168 8483
rect 8116 8440 8168 8449
rect 8760 8483 8812 8492
rect 8760 8449 8769 8483
rect 8769 8449 8803 8483
rect 8803 8449 8812 8483
rect 8760 8440 8812 8449
rect 2596 8236 2648 8288
rect 2688 8236 2740 8288
rect 4712 8415 4764 8424
rect 4712 8381 4721 8415
rect 4721 8381 4755 8415
rect 4755 8381 4764 8415
rect 4712 8372 4764 8381
rect 6092 8304 6144 8356
rect 6644 8236 6696 8288
rect 7472 8236 7524 8288
rect 7932 8347 7984 8356
rect 7932 8313 7941 8347
rect 7941 8313 7975 8347
rect 7975 8313 7984 8347
rect 7932 8304 7984 8313
rect 8392 8372 8444 8424
rect 8944 8372 8996 8424
rect 9220 8372 9272 8424
rect 9588 8372 9640 8424
rect 9956 8415 10008 8424
rect 9956 8381 9965 8415
rect 9965 8381 9999 8415
rect 9999 8381 10008 8415
rect 9956 8372 10008 8381
rect 10324 8483 10376 8492
rect 10324 8449 10333 8483
rect 10333 8449 10367 8483
rect 10367 8449 10376 8483
rect 10324 8440 10376 8449
rect 10968 8440 11020 8492
rect 11244 8372 11296 8424
rect 11428 8372 11480 8424
rect 11704 8440 11756 8492
rect 11980 8483 12032 8492
rect 11980 8449 11989 8483
rect 11989 8449 12023 8483
rect 12023 8449 12032 8483
rect 11980 8440 12032 8449
rect 12716 8440 12768 8492
rect 12808 8483 12860 8492
rect 12808 8449 12817 8483
rect 12817 8449 12851 8483
rect 12851 8449 12860 8483
rect 12808 8440 12860 8449
rect 13544 8483 13596 8492
rect 13544 8449 13553 8483
rect 13553 8449 13587 8483
rect 13587 8449 13596 8483
rect 13544 8440 13596 8449
rect 13728 8508 13780 8560
rect 14648 8508 14700 8560
rect 14740 8551 14792 8560
rect 14740 8517 14749 8551
rect 14749 8517 14783 8551
rect 14783 8517 14792 8551
rect 14740 8508 14792 8517
rect 16212 8576 16264 8628
rect 16764 8576 16816 8628
rect 17040 8576 17092 8628
rect 18328 8619 18380 8628
rect 18328 8585 18337 8619
rect 18337 8585 18371 8619
rect 18371 8585 18380 8619
rect 18328 8576 18380 8585
rect 18420 8576 18472 8628
rect 15936 8508 15988 8560
rect 12992 8372 13044 8424
rect 11520 8304 11572 8356
rect 11980 8304 12032 8356
rect 14096 8415 14148 8424
rect 14096 8381 14105 8415
rect 14105 8381 14139 8415
rect 14139 8381 14148 8415
rect 14096 8372 14148 8381
rect 14832 8440 14884 8492
rect 15292 8440 15344 8492
rect 15568 8440 15620 8492
rect 15752 8483 15804 8492
rect 15752 8449 15761 8483
rect 15761 8449 15795 8483
rect 15795 8449 15804 8483
rect 15752 8440 15804 8449
rect 16856 8508 16908 8560
rect 17500 8440 17552 8492
rect 8392 8236 8444 8288
rect 8760 8236 8812 8288
rect 9404 8236 9456 8288
rect 9772 8236 9824 8288
rect 10508 8236 10560 8288
rect 10784 8236 10836 8288
rect 11060 8236 11112 8288
rect 11888 8236 11940 8288
rect 12624 8279 12676 8288
rect 12624 8245 12633 8279
rect 12633 8245 12667 8279
rect 12667 8245 12676 8279
rect 12624 8236 12676 8245
rect 15660 8304 15712 8356
rect 14464 8236 14516 8288
rect 14832 8279 14884 8288
rect 14832 8245 14841 8279
rect 14841 8245 14875 8279
rect 14875 8245 14884 8279
rect 14832 8236 14884 8245
rect 14924 8236 14976 8288
rect 16028 8304 16080 8356
rect 16396 8372 16448 8424
rect 16672 8372 16724 8424
rect 17408 8415 17460 8424
rect 17408 8381 17417 8415
rect 17417 8381 17451 8415
rect 17451 8381 17460 8415
rect 17408 8372 17460 8381
rect 18236 8483 18288 8492
rect 18236 8449 18245 8483
rect 18245 8449 18279 8483
rect 18279 8449 18288 8483
rect 18236 8440 18288 8449
rect 18696 8415 18748 8424
rect 18696 8381 18705 8415
rect 18705 8381 18739 8415
rect 18739 8381 18748 8415
rect 18696 8372 18748 8381
rect 18972 8483 19024 8492
rect 18972 8449 18981 8483
rect 18981 8449 19015 8483
rect 19015 8449 19024 8483
rect 18972 8440 19024 8449
rect 19064 8483 19116 8492
rect 19064 8449 19073 8483
rect 19073 8449 19107 8483
rect 19107 8449 19116 8483
rect 19064 8440 19116 8449
rect 20904 8440 20956 8492
rect 21456 8483 21508 8492
rect 21456 8449 21465 8483
rect 21465 8449 21499 8483
rect 21499 8449 21508 8483
rect 21456 8440 21508 8449
rect 18604 8304 18656 8356
rect 18972 8304 19024 8356
rect 19524 8304 19576 8356
rect 20352 8415 20404 8424
rect 20352 8381 20361 8415
rect 20361 8381 20395 8415
rect 20395 8381 20404 8415
rect 20352 8372 20404 8381
rect 21088 8372 21140 8424
rect 21364 8372 21416 8424
rect 21640 8372 21692 8424
rect 22836 8440 22888 8492
rect 23204 8508 23256 8560
rect 24124 8576 24176 8628
rect 25228 8619 25280 8628
rect 25228 8585 25237 8619
rect 25237 8585 25271 8619
rect 25271 8585 25280 8619
rect 25228 8576 25280 8585
rect 23756 8508 23808 8560
rect 24492 8508 24544 8560
rect 24584 8508 24636 8560
rect 25872 8508 25924 8560
rect 22928 8372 22980 8424
rect 23204 8372 23256 8424
rect 23572 8372 23624 8424
rect 24308 8372 24360 8424
rect 21732 8304 21784 8356
rect 23388 8304 23440 8356
rect 24676 8372 24728 8424
rect 25688 8440 25740 8492
rect 27068 8483 27120 8492
rect 27068 8449 27077 8483
rect 27077 8449 27111 8483
rect 27111 8449 27120 8483
rect 27068 8440 27120 8449
rect 25780 8415 25832 8424
rect 25780 8381 25789 8415
rect 25789 8381 25823 8415
rect 25823 8381 25832 8415
rect 25780 8372 25832 8381
rect 26884 8372 26936 8424
rect 27252 8372 27304 8424
rect 28264 8576 28316 8628
rect 28908 8576 28960 8628
rect 29000 8576 29052 8628
rect 28080 8508 28132 8560
rect 28264 8440 28316 8492
rect 29828 8508 29880 8560
rect 29000 8440 29052 8492
rect 29092 8483 29144 8492
rect 29092 8449 29101 8483
rect 29101 8449 29135 8483
rect 29135 8449 29144 8483
rect 29092 8440 29144 8449
rect 29552 8440 29604 8492
rect 20904 8236 20956 8288
rect 23112 8236 23164 8288
rect 23204 8279 23256 8288
rect 23204 8245 23213 8279
rect 23213 8245 23247 8279
rect 23247 8245 23256 8279
rect 23204 8236 23256 8245
rect 23848 8236 23900 8288
rect 24860 8304 24912 8356
rect 25228 8304 25280 8356
rect 25320 8304 25372 8356
rect 24676 8236 24728 8288
rect 24768 8236 24820 8288
rect 25688 8236 25740 8288
rect 28264 8347 28316 8356
rect 28264 8313 28273 8347
rect 28273 8313 28307 8347
rect 28307 8313 28316 8347
rect 28264 8304 28316 8313
rect 28908 8304 28960 8356
rect 29092 8304 29144 8356
rect 29368 8347 29420 8356
rect 29368 8313 29377 8347
rect 29377 8313 29411 8347
rect 29411 8313 29420 8347
rect 29368 8304 29420 8313
rect 30104 8508 30156 8560
rect 30656 8551 30708 8560
rect 30656 8517 30665 8551
rect 30665 8517 30699 8551
rect 30699 8517 30708 8551
rect 30656 8508 30708 8517
rect 30932 8508 30984 8560
rect 30196 8483 30248 8492
rect 30196 8449 30205 8483
rect 30205 8449 30239 8483
rect 30239 8449 30248 8483
rect 30196 8440 30248 8449
rect 30380 8440 30432 8492
rect 30012 8372 30064 8424
rect 31392 8440 31444 8492
rect 31576 8483 31628 8492
rect 31576 8449 31585 8483
rect 31585 8449 31619 8483
rect 31619 8449 31628 8483
rect 31576 8440 31628 8449
rect 31760 8440 31812 8492
rect 32128 8483 32180 8492
rect 32128 8449 32137 8483
rect 32137 8449 32171 8483
rect 32171 8449 32180 8483
rect 32128 8440 32180 8449
rect 31116 8415 31168 8424
rect 31116 8381 31125 8415
rect 31125 8381 31159 8415
rect 31159 8381 31168 8415
rect 31116 8372 31168 8381
rect 31024 8347 31076 8356
rect 31024 8313 31033 8347
rect 31033 8313 31067 8347
rect 31067 8313 31076 8347
rect 31024 8304 31076 8313
rect 31208 8304 31260 8356
rect 31944 8304 31996 8356
rect 26792 8279 26844 8288
rect 26792 8245 26801 8279
rect 26801 8245 26835 8279
rect 26835 8245 26844 8279
rect 26792 8236 26844 8245
rect 27712 8236 27764 8288
rect 28724 8279 28776 8288
rect 28724 8245 28733 8279
rect 28733 8245 28767 8279
rect 28767 8245 28776 8279
rect 28724 8236 28776 8245
rect 29552 8279 29604 8288
rect 29552 8245 29561 8279
rect 29561 8245 29595 8279
rect 29595 8245 29604 8279
rect 29552 8236 29604 8245
rect 29736 8279 29788 8288
rect 29736 8245 29745 8279
rect 29745 8245 29779 8279
rect 29779 8245 29788 8279
rect 29736 8236 29788 8245
rect 29920 8236 29972 8288
rect 31760 8236 31812 8288
rect 32404 8372 32456 8424
rect 32496 8372 32548 8424
rect 32864 8576 32916 8628
rect 34520 8576 34572 8628
rect 33876 8508 33928 8560
rect 33048 8440 33100 8492
rect 33876 8372 33928 8424
rect 34152 8440 34204 8492
rect 34336 8483 34388 8492
rect 34336 8449 34345 8483
rect 34345 8449 34379 8483
rect 34379 8449 34388 8483
rect 34336 8440 34388 8449
rect 34888 8440 34940 8492
rect 35808 8576 35860 8628
rect 36912 8576 36964 8628
rect 37464 8508 37516 8560
rect 38568 8508 38620 8560
rect 35348 8483 35400 8492
rect 35348 8449 35357 8483
rect 35357 8449 35391 8483
rect 35391 8449 35400 8483
rect 35348 8440 35400 8449
rect 35716 8483 35768 8492
rect 35716 8449 35725 8483
rect 35725 8449 35759 8483
rect 35759 8449 35768 8483
rect 35716 8440 35768 8449
rect 35900 8440 35952 8492
rect 36728 8440 36780 8492
rect 36820 8483 36872 8492
rect 36820 8449 36829 8483
rect 36829 8449 36863 8483
rect 36863 8449 36872 8483
rect 36820 8440 36872 8449
rect 37280 8483 37332 8492
rect 37280 8449 37289 8483
rect 37289 8449 37323 8483
rect 37323 8449 37332 8483
rect 37280 8440 37332 8449
rect 37648 8440 37700 8492
rect 35164 8372 35216 8424
rect 32772 8304 32824 8356
rect 33600 8304 33652 8356
rect 34704 8304 34756 8356
rect 37832 8372 37884 8424
rect 38752 8440 38804 8492
rect 38844 8483 38896 8492
rect 38844 8449 38853 8483
rect 38853 8449 38887 8483
rect 38887 8449 38896 8483
rect 38844 8440 38896 8449
rect 36360 8304 36412 8356
rect 32864 8236 32916 8288
rect 33784 8279 33836 8288
rect 33784 8245 33793 8279
rect 33793 8245 33827 8279
rect 33827 8245 33836 8279
rect 33784 8236 33836 8245
rect 35256 8236 35308 8288
rect 37188 8304 37240 8356
rect 39028 8347 39080 8356
rect 39028 8313 39037 8347
rect 39037 8313 39071 8347
rect 39071 8313 39080 8347
rect 39028 8304 39080 8313
rect 39396 8347 39448 8356
rect 39396 8313 39405 8347
rect 39405 8313 39439 8347
rect 39439 8313 39448 8347
rect 39396 8304 39448 8313
rect 1950 8134 2002 8186
rect 2014 8134 2066 8186
rect 2078 8134 2130 8186
rect 2142 8134 2194 8186
rect 2206 8134 2258 8186
rect 7950 8134 8002 8186
rect 8014 8134 8066 8186
rect 8078 8134 8130 8186
rect 8142 8134 8194 8186
rect 8206 8134 8258 8186
rect 13950 8134 14002 8186
rect 14014 8134 14066 8186
rect 14078 8134 14130 8186
rect 14142 8134 14194 8186
rect 14206 8134 14258 8186
rect 19950 8134 20002 8186
rect 20014 8134 20066 8186
rect 20078 8134 20130 8186
rect 20142 8134 20194 8186
rect 20206 8134 20258 8186
rect 25950 8134 26002 8186
rect 26014 8134 26066 8186
rect 26078 8134 26130 8186
rect 26142 8134 26194 8186
rect 26206 8134 26258 8186
rect 31950 8134 32002 8186
rect 32014 8134 32066 8186
rect 32078 8134 32130 8186
rect 32142 8134 32194 8186
rect 32206 8134 32258 8186
rect 37950 8134 38002 8186
rect 38014 8134 38066 8186
rect 38078 8134 38130 8186
rect 38142 8134 38194 8186
rect 38206 8134 38258 8186
rect 4712 8032 4764 8084
rect 6920 8075 6972 8084
rect 6920 8041 6929 8075
rect 6929 8041 6963 8075
rect 6963 8041 6972 8075
rect 6920 8032 6972 8041
rect 11060 8032 11112 8084
rect 11152 8032 11204 8084
rect 12348 8032 12400 8084
rect 16580 8032 16632 8084
rect 16672 8075 16724 8084
rect 16672 8041 16681 8075
rect 16681 8041 16715 8075
rect 16715 8041 16724 8075
rect 16672 8032 16724 8041
rect 17316 8032 17368 8084
rect 18328 8032 18380 8084
rect 18604 8032 18656 8084
rect 20168 8032 20220 8084
rect 4896 7964 4948 8016
rect 1216 7896 1268 7948
rect 756 7828 808 7880
rect 2412 7828 2464 7880
rect 2596 7871 2648 7880
rect 2596 7837 2605 7871
rect 2605 7837 2639 7871
rect 2639 7837 2648 7871
rect 2596 7828 2648 7837
rect 2504 7760 2556 7812
rect 4068 7871 4120 7880
rect 4068 7837 4077 7871
rect 4077 7837 4111 7871
rect 4111 7837 4120 7871
rect 4068 7828 4120 7837
rect 5172 7896 5224 7948
rect 7656 7964 7708 8016
rect 3884 7760 3936 7812
rect 5632 7828 5684 7880
rect 5908 7828 5960 7880
rect 7932 7896 7984 7948
rect 7748 7828 7800 7880
rect 8116 7871 8168 7880
rect 8116 7837 8125 7871
rect 8125 7837 8159 7871
rect 8159 7837 8168 7871
rect 8116 7828 8168 7837
rect 8392 7871 8444 7880
rect 8392 7837 8401 7871
rect 8401 7837 8435 7871
rect 8435 7837 8444 7871
rect 8392 7828 8444 7837
rect 8944 7939 8996 7948
rect 8944 7905 8953 7939
rect 8953 7905 8987 7939
rect 8987 7905 8996 7939
rect 8944 7896 8996 7905
rect 13452 7896 13504 7948
rect 14648 7964 14700 8016
rect 2780 7692 2832 7744
rect 6644 7760 6696 7812
rect 4896 7735 4948 7744
rect 4896 7701 4905 7735
rect 4905 7701 4939 7735
rect 4939 7701 4948 7735
rect 4896 7692 4948 7701
rect 6552 7692 6604 7744
rect 7748 7692 7800 7744
rect 10508 7871 10560 7880
rect 10508 7837 10517 7871
rect 10517 7837 10551 7871
rect 10551 7837 10560 7871
rect 10508 7828 10560 7837
rect 10600 7828 10652 7880
rect 8944 7760 8996 7812
rect 9680 7760 9732 7812
rect 12440 7828 12492 7880
rect 12624 7871 12676 7880
rect 12624 7837 12658 7871
rect 12658 7837 12676 7871
rect 12624 7828 12676 7837
rect 13176 7828 13228 7880
rect 13728 7828 13780 7880
rect 11060 7803 11112 7812
rect 11060 7769 11094 7803
rect 11094 7769 11112 7803
rect 11060 7760 11112 7769
rect 10324 7735 10376 7744
rect 10324 7701 10333 7735
rect 10333 7701 10367 7735
rect 10367 7701 10376 7735
rect 10324 7692 10376 7701
rect 13912 7760 13964 7812
rect 13728 7735 13780 7744
rect 13728 7701 13737 7735
rect 13737 7701 13771 7735
rect 13771 7701 13780 7735
rect 13728 7692 13780 7701
rect 14188 7760 14240 7812
rect 14464 7828 14516 7880
rect 14648 7871 14700 7880
rect 14648 7837 14657 7871
rect 14657 7837 14691 7871
rect 14691 7837 14700 7871
rect 14648 7828 14700 7837
rect 15108 7871 15160 7880
rect 15108 7837 15117 7871
rect 15117 7837 15151 7871
rect 15151 7837 15160 7871
rect 15108 7828 15160 7837
rect 15752 7828 15804 7880
rect 17040 7964 17092 8016
rect 17408 7828 17460 7880
rect 18052 7871 18104 7880
rect 18052 7837 18061 7871
rect 18061 7837 18095 7871
rect 18095 7837 18104 7871
rect 18052 7828 18104 7837
rect 22376 7964 22428 8016
rect 23020 7964 23072 8016
rect 18512 7896 18564 7948
rect 21456 7896 21508 7948
rect 18604 7871 18656 7880
rect 18604 7837 18613 7871
rect 18613 7837 18647 7871
rect 18647 7837 18656 7871
rect 18604 7828 18656 7837
rect 15844 7760 15896 7812
rect 18880 7871 18932 7880
rect 18880 7837 18889 7871
rect 18889 7837 18923 7871
rect 18923 7837 18932 7871
rect 18880 7828 18932 7837
rect 20260 7828 20312 7880
rect 21916 7828 21968 7880
rect 24584 7896 24636 7948
rect 25044 8032 25096 8084
rect 28908 8032 28960 8084
rect 29736 8032 29788 8084
rect 29828 8032 29880 8084
rect 30196 8075 30248 8084
rect 30196 8041 30205 8075
rect 30205 8041 30239 8075
rect 30239 8041 30248 8075
rect 30196 8032 30248 8041
rect 27804 7964 27856 8016
rect 28724 8007 28776 8016
rect 28724 7973 28733 8007
rect 28733 7973 28767 8007
rect 28767 7973 28776 8007
rect 28724 7964 28776 7973
rect 25044 7896 25096 7948
rect 25504 7896 25556 7948
rect 24124 7828 24176 7880
rect 27068 7828 27120 7880
rect 27528 7828 27580 7880
rect 29184 8007 29236 8016
rect 29184 7973 29193 8007
rect 29193 7973 29227 8007
rect 29227 7973 29236 8007
rect 29184 7964 29236 7973
rect 29368 7964 29420 8016
rect 31208 8032 31260 8084
rect 31576 8032 31628 8084
rect 33048 8032 33100 8084
rect 33416 8032 33468 8084
rect 34520 8032 34572 8084
rect 35532 8032 35584 8084
rect 36084 8032 36136 8084
rect 36636 8032 36688 8084
rect 37740 8032 37792 8084
rect 38660 8075 38712 8084
rect 38660 8041 38669 8075
rect 38669 8041 38703 8075
rect 38703 8041 38712 8075
rect 38660 8032 38712 8041
rect 31760 7964 31812 8016
rect 32496 7964 32548 8016
rect 32772 7964 32824 8016
rect 30472 7939 30524 7948
rect 30472 7905 30481 7939
rect 30481 7905 30515 7939
rect 30515 7905 30524 7939
rect 30472 7896 30524 7905
rect 19340 7760 19392 7812
rect 19432 7760 19484 7812
rect 15476 7692 15528 7744
rect 16580 7692 16632 7744
rect 17960 7692 18012 7744
rect 18972 7692 19024 7744
rect 19800 7692 19852 7744
rect 20168 7803 20220 7812
rect 20168 7769 20177 7803
rect 20177 7769 20211 7803
rect 20211 7769 20220 7803
rect 20168 7760 20220 7769
rect 20352 7803 20404 7812
rect 20352 7769 20361 7803
rect 20361 7769 20395 7803
rect 20395 7769 20404 7803
rect 20352 7760 20404 7769
rect 22560 7760 22612 7812
rect 24492 7803 24544 7812
rect 24492 7769 24501 7803
rect 24501 7769 24535 7803
rect 24535 7769 24544 7803
rect 24492 7760 24544 7769
rect 24952 7760 25004 7812
rect 25872 7760 25924 7812
rect 26240 7803 26292 7812
rect 26240 7769 26249 7803
rect 26249 7769 26283 7803
rect 26283 7769 26292 7803
rect 26240 7760 26292 7769
rect 20996 7692 21048 7744
rect 21088 7692 21140 7744
rect 22744 7692 22796 7744
rect 27988 7692 28040 7744
rect 28356 7871 28408 7880
rect 28356 7837 28365 7871
rect 28365 7837 28399 7871
rect 28399 7837 28408 7871
rect 28356 7828 28408 7837
rect 28448 7828 28500 7880
rect 28908 7871 28960 7880
rect 28908 7837 28917 7871
rect 28917 7837 28951 7871
rect 28951 7837 28960 7871
rect 28908 7828 28960 7837
rect 28816 7760 28868 7812
rect 29644 7828 29696 7880
rect 30564 7828 30616 7880
rect 31484 7828 31536 7880
rect 31760 7828 31812 7880
rect 32220 7871 32272 7880
rect 32220 7837 32229 7871
rect 32229 7837 32263 7871
rect 32263 7837 32272 7871
rect 32220 7828 32272 7837
rect 32588 7828 32640 7880
rect 33232 7828 33284 7880
rect 33508 7828 33560 7880
rect 29368 7692 29420 7744
rect 30564 7692 30616 7744
rect 31392 7692 31444 7744
rect 32772 7760 32824 7812
rect 32956 7760 33008 7812
rect 33692 7760 33744 7812
rect 36360 7828 36412 7880
rect 36452 7871 36504 7880
rect 36452 7837 36461 7871
rect 36461 7837 36495 7871
rect 36495 7837 36504 7871
rect 36452 7828 36504 7837
rect 37004 7871 37056 7880
rect 37004 7837 37013 7871
rect 37013 7837 37047 7871
rect 37047 7837 37056 7871
rect 37004 7828 37056 7837
rect 37372 7828 37424 7880
rect 37556 7760 37608 7812
rect 37740 7760 37792 7812
rect 39304 7828 39356 7880
rect 31944 7692 31996 7744
rect 32128 7692 32180 7744
rect 33600 7735 33652 7744
rect 33600 7701 33609 7735
rect 33609 7701 33643 7735
rect 33643 7701 33652 7735
rect 33600 7692 33652 7701
rect 38936 7692 38988 7744
rect 39396 7735 39448 7744
rect 39396 7701 39405 7735
rect 39405 7701 39439 7735
rect 39439 7701 39448 7735
rect 39396 7692 39448 7701
rect 3010 7590 3062 7642
rect 3074 7590 3126 7642
rect 3138 7590 3190 7642
rect 3202 7590 3254 7642
rect 3266 7590 3318 7642
rect 9010 7590 9062 7642
rect 9074 7590 9126 7642
rect 9138 7590 9190 7642
rect 9202 7590 9254 7642
rect 9266 7590 9318 7642
rect 15010 7590 15062 7642
rect 15074 7590 15126 7642
rect 15138 7590 15190 7642
rect 15202 7590 15254 7642
rect 15266 7590 15318 7642
rect 21010 7590 21062 7642
rect 21074 7590 21126 7642
rect 21138 7590 21190 7642
rect 21202 7590 21254 7642
rect 21266 7590 21318 7642
rect 27010 7590 27062 7642
rect 27074 7590 27126 7642
rect 27138 7590 27190 7642
rect 27202 7590 27254 7642
rect 27266 7590 27318 7642
rect 33010 7590 33062 7642
rect 33074 7590 33126 7642
rect 33138 7590 33190 7642
rect 33202 7590 33254 7642
rect 33266 7590 33318 7642
rect 39010 7590 39062 7642
rect 39074 7590 39126 7642
rect 39138 7590 39190 7642
rect 39202 7590 39254 7642
rect 39266 7590 39318 7642
rect 2504 7531 2556 7540
rect 2504 7497 2513 7531
rect 2513 7497 2547 7531
rect 2547 7497 2556 7531
rect 2504 7488 2556 7497
rect 2688 7531 2740 7540
rect 2688 7497 2697 7531
rect 2697 7497 2731 7531
rect 2731 7497 2740 7531
rect 2688 7488 2740 7497
rect 3424 7488 3476 7540
rect 4988 7531 5040 7540
rect 4988 7497 4997 7531
rect 4997 7497 5031 7531
rect 5031 7497 5040 7531
rect 4988 7488 5040 7497
rect 5172 7531 5224 7540
rect 5172 7497 5181 7531
rect 5181 7497 5215 7531
rect 5215 7497 5224 7531
rect 5172 7488 5224 7497
rect 8852 7488 8904 7540
rect 9496 7488 9548 7540
rect 10600 7488 10652 7540
rect 10876 7488 10928 7540
rect 15936 7488 15988 7540
rect 16580 7488 16632 7540
rect 17868 7488 17920 7540
rect 18512 7531 18564 7540
rect 18512 7497 18521 7531
rect 18521 7497 18555 7531
rect 18555 7497 18564 7531
rect 18512 7488 18564 7497
rect 18604 7488 18656 7540
rect 19616 7488 19668 7540
rect 756 7352 808 7404
rect 4896 7420 4948 7472
rect 7012 7463 7064 7472
rect 7012 7429 7021 7463
rect 7021 7429 7055 7463
rect 7055 7429 7064 7463
rect 7012 7420 7064 7429
rect 1584 7284 1636 7336
rect 2780 7284 2832 7336
rect 3148 7352 3200 7404
rect 4068 7352 4120 7404
rect 5908 7395 5960 7404
rect 3332 7327 3384 7336
rect 3332 7293 3341 7327
rect 3341 7293 3375 7327
rect 3375 7293 3384 7327
rect 3332 7284 3384 7293
rect 3976 7284 4028 7336
rect 5908 7361 5917 7395
rect 5917 7361 5951 7395
rect 5951 7361 5960 7395
rect 5908 7352 5960 7361
rect 6644 7352 6696 7404
rect 6828 7395 6880 7404
rect 6828 7361 6837 7395
rect 6837 7361 6871 7395
rect 6871 7361 6880 7395
rect 6828 7352 6880 7361
rect 8392 7420 8444 7472
rect 9680 7420 9732 7472
rect 7656 7352 7708 7404
rect 6368 7284 6420 7336
rect 3240 7216 3292 7268
rect 7472 7284 7524 7336
rect 7932 7216 7984 7268
rect 4344 7191 4396 7200
rect 4344 7157 4353 7191
rect 4353 7157 4387 7191
rect 4387 7157 4396 7191
rect 4344 7148 4396 7157
rect 7196 7148 7248 7200
rect 8300 7395 8352 7404
rect 8300 7361 8309 7395
rect 8309 7361 8343 7395
rect 8343 7361 8352 7395
rect 8300 7352 8352 7361
rect 8852 7352 8904 7404
rect 10508 7420 10560 7472
rect 12992 7420 13044 7472
rect 11704 7395 11756 7404
rect 11704 7361 11713 7395
rect 11713 7361 11747 7395
rect 11747 7361 11756 7395
rect 11704 7352 11756 7361
rect 12716 7352 12768 7404
rect 14648 7420 14700 7472
rect 16212 7420 16264 7472
rect 13544 7352 13596 7404
rect 9680 7284 9732 7336
rect 11520 7327 11572 7336
rect 11520 7293 11529 7327
rect 11529 7293 11563 7327
rect 11563 7293 11572 7327
rect 11520 7284 11572 7293
rect 13360 7327 13412 7336
rect 13360 7293 13369 7327
rect 13369 7293 13403 7327
rect 13403 7293 13412 7327
rect 13360 7284 13412 7293
rect 15292 7352 15344 7404
rect 15384 7395 15436 7404
rect 15384 7361 15393 7395
rect 15393 7361 15427 7395
rect 15427 7361 15436 7395
rect 15384 7352 15436 7361
rect 15568 7352 15620 7404
rect 15844 7395 15896 7404
rect 15844 7361 15853 7395
rect 15853 7361 15887 7395
rect 15887 7361 15896 7395
rect 15844 7352 15896 7361
rect 16028 7352 16080 7404
rect 16672 7463 16724 7472
rect 16672 7429 16681 7463
rect 16681 7429 16715 7463
rect 16715 7429 16724 7463
rect 16672 7420 16724 7429
rect 17040 7420 17092 7472
rect 18052 7420 18104 7472
rect 8668 7148 8720 7200
rect 9496 7148 9548 7200
rect 9956 7148 10008 7200
rect 10324 7148 10376 7200
rect 11428 7148 11480 7200
rect 11888 7191 11940 7200
rect 11888 7157 11897 7191
rect 11897 7157 11931 7191
rect 11931 7157 11940 7191
rect 11888 7148 11940 7157
rect 11980 7191 12032 7200
rect 11980 7157 11989 7191
rect 11989 7157 12023 7191
rect 12023 7157 12032 7191
rect 11980 7148 12032 7157
rect 13820 7191 13872 7200
rect 13820 7157 13829 7191
rect 13829 7157 13863 7191
rect 13863 7157 13872 7191
rect 13820 7148 13872 7157
rect 14280 7148 14332 7200
rect 14556 7148 14608 7200
rect 15936 7216 15988 7268
rect 16028 7191 16080 7200
rect 16028 7157 16037 7191
rect 16037 7157 16071 7191
rect 16071 7157 16080 7191
rect 16028 7148 16080 7157
rect 16672 7148 16724 7200
rect 16856 7191 16908 7200
rect 16856 7157 16865 7191
rect 16865 7157 16899 7191
rect 16899 7157 16908 7191
rect 16856 7148 16908 7157
rect 19064 7395 19116 7404
rect 19064 7361 19098 7395
rect 19098 7361 19116 7395
rect 19064 7352 19116 7361
rect 20352 7352 20404 7404
rect 21640 7531 21692 7540
rect 21640 7497 21649 7531
rect 21649 7497 21683 7531
rect 21683 7497 21692 7531
rect 21640 7488 21692 7497
rect 22100 7488 22152 7540
rect 23296 7488 23348 7540
rect 23480 7488 23532 7540
rect 22928 7420 22980 7472
rect 23204 7420 23256 7472
rect 21364 7352 21416 7404
rect 22652 7352 22704 7404
rect 23388 7352 23440 7404
rect 24124 7395 24176 7404
rect 24124 7361 24133 7395
rect 24133 7361 24167 7395
rect 24167 7361 24176 7395
rect 24124 7352 24176 7361
rect 24952 7531 25004 7540
rect 24952 7497 24961 7531
rect 24961 7497 24995 7531
rect 24995 7497 25004 7531
rect 24952 7488 25004 7497
rect 26516 7488 26568 7540
rect 29000 7488 29052 7540
rect 26240 7463 26292 7472
rect 26240 7429 26249 7463
rect 26249 7429 26283 7463
rect 26283 7429 26292 7463
rect 26240 7420 26292 7429
rect 27528 7420 27580 7472
rect 25688 7352 25740 7404
rect 26424 7284 26476 7336
rect 26792 7352 26844 7404
rect 29552 7420 29604 7472
rect 30012 7531 30064 7540
rect 30012 7497 30021 7531
rect 30021 7497 30055 7531
rect 30055 7497 30064 7531
rect 30012 7488 30064 7497
rect 31484 7488 31536 7540
rect 32956 7531 33008 7540
rect 32956 7497 32965 7531
rect 32965 7497 32999 7531
rect 32999 7497 33008 7531
rect 32956 7488 33008 7497
rect 33048 7488 33100 7540
rect 29828 7420 29880 7472
rect 32128 7420 32180 7472
rect 32220 7420 32272 7472
rect 28540 7352 28592 7404
rect 29368 7352 29420 7404
rect 29644 7395 29696 7404
rect 29644 7361 29653 7395
rect 29653 7361 29687 7395
rect 29687 7361 29696 7395
rect 29644 7352 29696 7361
rect 30104 7395 30156 7404
rect 30104 7361 30113 7395
rect 30113 7361 30147 7395
rect 30147 7361 30156 7395
rect 30104 7352 30156 7361
rect 30472 7352 30524 7404
rect 18788 7216 18840 7268
rect 22376 7216 22428 7268
rect 18604 7148 18656 7200
rect 20168 7148 20220 7200
rect 22192 7148 22244 7200
rect 22652 7148 22704 7200
rect 24124 7216 24176 7268
rect 25780 7148 25832 7200
rect 27068 7148 27120 7200
rect 29736 7327 29788 7336
rect 29736 7293 29745 7327
rect 29745 7293 29779 7327
rect 29779 7293 29788 7327
rect 29736 7284 29788 7293
rect 31944 7284 31996 7336
rect 32588 7395 32640 7404
rect 32588 7361 32597 7395
rect 32597 7361 32631 7395
rect 32631 7361 32640 7395
rect 32588 7352 32640 7361
rect 32772 7352 32824 7404
rect 34428 7488 34480 7540
rect 36452 7488 36504 7540
rect 34152 7420 34204 7472
rect 34612 7420 34664 7472
rect 38844 7488 38896 7540
rect 39580 7488 39632 7540
rect 33968 7395 34020 7404
rect 33968 7361 33977 7395
rect 33977 7361 34011 7395
rect 34011 7361 34020 7395
rect 33968 7352 34020 7361
rect 34244 7395 34296 7404
rect 34244 7361 34253 7395
rect 34253 7361 34287 7395
rect 34287 7361 34296 7395
rect 34244 7352 34296 7361
rect 34520 7395 34572 7404
rect 34520 7361 34529 7395
rect 34529 7361 34563 7395
rect 34563 7361 34572 7395
rect 34520 7352 34572 7361
rect 39764 7420 39816 7472
rect 32220 7259 32272 7268
rect 32220 7225 32229 7259
rect 32229 7225 32263 7259
rect 32263 7225 32272 7259
rect 32220 7216 32272 7225
rect 31944 7148 31996 7200
rect 32496 7148 32548 7200
rect 33232 7259 33284 7268
rect 33232 7225 33241 7259
rect 33241 7225 33275 7259
rect 33275 7225 33284 7259
rect 33232 7216 33284 7225
rect 33784 7284 33836 7336
rect 38292 7352 38344 7404
rect 38568 7216 38620 7268
rect 33784 7191 33836 7200
rect 33784 7157 33793 7191
rect 33793 7157 33827 7191
rect 33827 7157 33836 7191
rect 33784 7148 33836 7157
rect 34796 7148 34848 7200
rect 35992 7148 36044 7200
rect 39212 7395 39264 7404
rect 39212 7361 39221 7395
rect 39221 7361 39255 7395
rect 39255 7361 39264 7395
rect 39212 7352 39264 7361
rect 39396 7191 39448 7200
rect 39396 7157 39405 7191
rect 39405 7157 39439 7191
rect 39439 7157 39448 7191
rect 39396 7148 39448 7157
rect 1950 7046 2002 7098
rect 2014 7046 2066 7098
rect 2078 7046 2130 7098
rect 2142 7046 2194 7098
rect 2206 7046 2258 7098
rect 7950 7046 8002 7098
rect 8014 7046 8066 7098
rect 8078 7046 8130 7098
rect 8142 7046 8194 7098
rect 8206 7046 8258 7098
rect 13950 7046 14002 7098
rect 14014 7046 14066 7098
rect 14078 7046 14130 7098
rect 14142 7046 14194 7098
rect 14206 7046 14258 7098
rect 19950 7046 20002 7098
rect 20014 7046 20066 7098
rect 20078 7046 20130 7098
rect 20142 7046 20194 7098
rect 20206 7046 20258 7098
rect 25950 7046 26002 7098
rect 26014 7046 26066 7098
rect 26078 7046 26130 7098
rect 26142 7046 26194 7098
rect 26206 7046 26258 7098
rect 31950 7046 32002 7098
rect 32014 7046 32066 7098
rect 32078 7046 32130 7098
rect 32142 7046 32194 7098
rect 32206 7046 32258 7098
rect 37950 7046 38002 7098
rect 38014 7046 38066 7098
rect 38078 7046 38130 7098
rect 38142 7046 38194 7098
rect 38206 7046 38258 7098
rect 3608 6944 3660 6996
rect 3884 6944 3936 6996
rect 5448 6944 5500 6996
rect 1400 6808 1452 6860
rect 3240 6876 3292 6928
rect 1676 6672 1728 6724
rect 3148 6808 3200 6860
rect 3240 6783 3292 6792
rect 3240 6749 3249 6783
rect 3249 6749 3283 6783
rect 3283 6749 3292 6783
rect 3240 6740 3292 6749
rect 4068 6876 4120 6928
rect 4252 6876 4304 6928
rect 4344 6876 4396 6928
rect 7748 6944 7800 6996
rect 3516 6808 3568 6860
rect 4252 6783 4304 6792
rect 4252 6749 4261 6783
rect 4261 6749 4295 6783
rect 4295 6749 4304 6783
rect 4252 6740 4304 6749
rect 5172 6808 5224 6860
rect 6552 6808 6604 6860
rect 8852 6876 8904 6928
rect 4988 6783 5040 6792
rect 4988 6749 4997 6783
rect 4997 6749 5031 6783
rect 5031 6749 5040 6783
rect 4988 6740 5040 6749
rect 5448 6783 5500 6792
rect 5448 6749 5457 6783
rect 5457 6749 5491 6783
rect 5491 6749 5500 6783
rect 5448 6740 5500 6749
rect 5816 6740 5868 6792
rect 6920 6783 6972 6792
rect 6920 6749 6929 6783
rect 6929 6749 6963 6783
rect 6963 6749 6972 6783
rect 6920 6740 6972 6749
rect 1768 6647 1820 6656
rect 1768 6613 1777 6647
rect 1777 6613 1811 6647
rect 1811 6613 1820 6647
rect 1768 6604 1820 6613
rect 2228 6647 2280 6656
rect 2228 6613 2237 6647
rect 2237 6613 2271 6647
rect 2271 6613 2280 6647
rect 2228 6604 2280 6613
rect 3332 6604 3384 6656
rect 3792 6604 3844 6656
rect 3884 6647 3936 6656
rect 3884 6613 3893 6647
rect 3893 6613 3927 6647
rect 3927 6613 3936 6647
rect 3884 6604 3936 6613
rect 6828 6672 6880 6724
rect 4712 6604 4764 6656
rect 5172 6647 5224 6656
rect 5172 6613 5181 6647
rect 5181 6613 5215 6647
rect 5215 6613 5224 6647
rect 5172 6604 5224 6613
rect 5264 6604 5316 6656
rect 6920 6604 6972 6656
rect 8852 6740 8904 6792
rect 9588 6740 9640 6792
rect 9680 6740 9732 6792
rect 10876 6876 10928 6928
rect 11060 6987 11112 6996
rect 11060 6953 11069 6987
rect 11069 6953 11103 6987
rect 11103 6953 11112 6987
rect 11060 6944 11112 6953
rect 11704 6944 11756 6996
rect 12440 6944 12492 6996
rect 13360 6944 13412 6996
rect 7748 6672 7800 6724
rect 8116 6672 8168 6724
rect 8668 6672 8720 6724
rect 10600 6783 10652 6792
rect 10600 6749 10609 6783
rect 10609 6749 10643 6783
rect 10643 6749 10652 6783
rect 10600 6740 10652 6749
rect 10692 6783 10744 6792
rect 10692 6749 10701 6783
rect 10701 6749 10735 6783
rect 10735 6749 10744 6783
rect 10692 6740 10744 6749
rect 11152 6740 11204 6792
rect 11336 6808 11388 6860
rect 11980 6808 12032 6860
rect 12808 6876 12860 6928
rect 13636 6876 13688 6928
rect 12348 6740 12400 6792
rect 12808 6740 12860 6792
rect 14556 6808 14608 6860
rect 18236 6944 18288 6996
rect 15660 6851 15712 6860
rect 15660 6817 15669 6851
rect 15669 6817 15703 6851
rect 15703 6817 15712 6851
rect 15660 6808 15712 6817
rect 17316 6808 17368 6860
rect 17592 6808 17644 6860
rect 13912 6783 13964 6792
rect 13912 6749 13921 6783
rect 13921 6749 13955 6783
rect 13955 6749 13964 6783
rect 13912 6740 13964 6749
rect 7656 6604 7708 6656
rect 10876 6672 10928 6724
rect 12164 6672 12216 6724
rect 13636 6715 13688 6724
rect 13636 6681 13645 6715
rect 13645 6681 13679 6715
rect 13679 6681 13688 6715
rect 13636 6672 13688 6681
rect 15476 6672 15528 6724
rect 16672 6783 16724 6792
rect 16672 6749 16681 6783
rect 16681 6749 16715 6783
rect 16715 6749 16724 6783
rect 16672 6740 16724 6749
rect 17224 6783 17276 6792
rect 17224 6749 17233 6783
rect 17233 6749 17267 6783
rect 17267 6749 17276 6783
rect 17224 6740 17276 6749
rect 17500 6740 17552 6792
rect 18144 6919 18196 6928
rect 18144 6885 18153 6919
rect 18153 6885 18187 6919
rect 18187 6885 18196 6919
rect 18144 6876 18196 6885
rect 18512 6876 18564 6928
rect 22284 6944 22336 6996
rect 23572 6944 23624 6996
rect 25412 6944 25464 6996
rect 26700 6944 26752 6996
rect 18236 6851 18288 6860
rect 18236 6817 18245 6851
rect 18245 6817 18279 6851
rect 18279 6817 18288 6851
rect 18236 6808 18288 6817
rect 18604 6808 18656 6860
rect 19064 6876 19116 6928
rect 22008 6876 22060 6928
rect 17960 6740 18012 6792
rect 10140 6604 10192 6656
rect 10600 6604 10652 6656
rect 11244 6604 11296 6656
rect 13544 6604 13596 6656
rect 14188 6647 14240 6656
rect 14188 6613 14197 6647
rect 14197 6613 14231 6647
rect 14231 6613 14240 6647
rect 14188 6604 14240 6613
rect 14280 6604 14332 6656
rect 15660 6604 15712 6656
rect 16028 6604 16080 6656
rect 16764 6604 16816 6656
rect 17132 6604 17184 6656
rect 17224 6604 17276 6656
rect 17684 6647 17736 6656
rect 17684 6613 17693 6647
rect 17693 6613 17727 6647
rect 17727 6613 17736 6647
rect 17684 6604 17736 6613
rect 17868 6672 17920 6724
rect 19156 6740 19208 6792
rect 20352 6808 20404 6860
rect 22284 6808 22336 6860
rect 23848 6876 23900 6928
rect 26884 6919 26936 6928
rect 26884 6885 26893 6919
rect 26893 6885 26927 6919
rect 26927 6885 26936 6919
rect 26884 6876 26936 6885
rect 19432 6672 19484 6724
rect 19616 6783 19668 6792
rect 19616 6749 19625 6783
rect 19625 6749 19659 6783
rect 19659 6749 19668 6783
rect 19616 6740 19668 6749
rect 21364 6740 21416 6792
rect 22744 6740 22796 6792
rect 22928 6740 22980 6792
rect 23480 6783 23532 6792
rect 23480 6749 23489 6783
rect 23489 6749 23523 6783
rect 23523 6749 23532 6783
rect 23480 6740 23532 6749
rect 23572 6740 23624 6792
rect 20260 6672 20312 6724
rect 22284 6672 22336 6724
rect 21732 6604 21784 6656
rect 22008 6604 22060 6656
rect 22652 6647 22704 6656
rect 22652 6613 22661 6647
rect 22661 6613 22695 6647
rect 22695 6613 22704 6647
rect 22652 6604 22704 6613
rect 22928 6604 22980 6656
rect 23112 6647 23164 6656
rect 23112 6613 23121 6647
rect 23121 6613 23155 6647
rect 23155 6613 23164 6647
rect 23112 6604 23164 6613
rect 23940 6647 23992 6656
rect 23940 6613 23949 6647
rect 23949 6613 23983 6647
rect 23983 6613 23992 6647
rect 23940 6604 23992 6613
rect 24124 6672 24176 6724
rect 24676 6783 24728 6792
rect 24676 6749 24685 6783
rect 24685 6749 24719 6783
rect 24719 6749 24728 6783
rect 24676 6740 24728 6749
rect 24768 6740 24820 6792
rect 27528 6808 27580 6860
rect 25136 6740 25188 6792
rect 26240 6740 26292 6792
rect 24768 6604 24820 6656
rect 24860 6604 24912 6656
rect 25504 6647 25556 6656
rect 25504 6613 25513 6647
rect 25513 6613 25547 6647
rect 25547 6613 25556 6647
rect 25504 6604 25556 6613
rect 25964 6672 26016 6724
rect 26700 6672 26752 6724
rect 27068 6783 27120 6792
rect 27068 6749 27077 6783
rect 27077 6749 27111 6783
rect 27111 6749 27120 6783
rect 27068 6740 27120 6749
rect 27344 6783 27396 6792
rect 27344 6749 27353 6783
rect 27353 6749 27387 6783
rect 27387 6749 27396 6783
rect 27344 6740 27396 6749
rect 27620 6783 27672 6792
rect 27620 6749 27629 6783
rect 27629 6749 27663 6783
rect 27663 6749 27672 6783
rect 27620 6740 27672 6749
rect 28264 6740 28316 6792
rect 30104 6944 30156 6996
rect 31116 6944 31168 6996
rect 32312 6944 32364 6996
rect 34520 6987 34572 6996
rect 34520 6953 34529 6987
rect 34529 6953 34563 6987
rect 34563 6953 34572 6987
rect 34520 6944 34572 6953
rect 35808 6944 35860 6996
rect 39212 6944 39264 6996
rect 29092 6808 29144 6860
rect 31024 6919 31076 6928
rect 31024 6885 31033 6919
rect 31033 6885 31067 6919
rect 31067 6885 31076 6919
rect 31024 6876 31076 6885
rect 30472 6808 30524 6860
rect 31208 6808 31260 6860
rect 31392 6851 31444 6860
rect 31392 6817 31401 6851
rect 31401 6817 31435 6851
rect 31435 6817 31444 6851
rect 31392 6808 31444 6817
rect 31668 6808 31720 6860
rect 35716 6876 35768 6928
rect 37280 6876 37332 6928
rect 29460 6740 29512 6792
rect 29828 6783 29880 6792
rect 29828 6749 29837 6783
rect 29837 6749 29871 6783
rect 29871 6749 29880 6783
rect 29828 6740 29880 6749
rect 30196 6740 30248 6792
rect 27712 6672 27764 6724
rect 28632 6672 28684 6724
rect 30564 6740 30616 6792
rect 31484 6783 31536 6792
rect 31484 6749 31493 6783
rect 31493 6749 31527 6783
rect 31527 6749 31536 6783
rect 31484 6740 31536 6749
rect 35900 6808 35952 6860
rect 32036 6740 32088 6792
rect 32404 6740 32456 6792
rect 30840 6672 30892 6724
rect 31668 6672 31720 6724
rect 32956 6783 33008 6792
rect 32956 6749 32965 6783
rect 32965 6749 32999 6783
rect 32999 6749 33008 6783
rect 32956 6740 33008 6749
rect 35440 6740 35492 6792
rect 36084 6740 36136 6792
rect 36176 6740 36228 6792
rect 38476 6783 38528 6792
rect 38476 6749 38485 6783
rect 38485 6749 38519 6783
rect 38519 6749 38528 6783
rect 38476 6740 38528 6749
rect 38844 6783 38896 6792
rect 38844 6749 38853 6783
rect 38853 6749 38887 6783
rect 38887 6749 38896 6783
rect 38844 6740 38896 6749
rect 32772 6672 32824 6724
rect 34796 6672 34848 6724
rect 26884 6604 26936 6656
rect 27344 6604 27396 6656
rect 29000 6604 29052 6656
rect 29644 6604 29696 6656
rect 29920 6604 29972 6656
rect 30656 6604 30708 6656
rect 31852 6604 31904 6656
rect 32036 6647 32088 6656
rect 32036 6613 32045 6647
rect 32045 6613 32079 6647
rect 32079 6613 32088 6647
rect 32036 6604 32088 6613
rect 32312 6647 32364 6656
rect 32312 6613 32321 6647
rect 32321 6613 32355 6647
rect 32355 6613 32364 6647
rect 32312 6604 32364 6613
rect 34060 6647 34112 6656
rect 34060 6613 34069 6647
rect 34069 6613 34103 6647
rect 34103 6613 34112 6647
rect 34060 6604 34112 6613
rect 34152 6647 34204 6656
rect 34152 6613 34161 6647
rect 34161 6613 34195 6647
rect 34195 6613 34204 6647
rect 34152 6604 34204 6613
rect 35624 6604 35676 6656
rect 36728 6604 36780 6656
rect 38016 6647 38068 6656
rect 38016 6613 38025 6647
rect 38025 6613 38059 6647
rect 38059 6613 38068 6647
rect 38016 6604 38068 6613
rect 38660 6647 38712 6656
rect 38660 6613 38669 6647
rect 38669 6613 38703 6647
rect 38703 6613 38712 6647
rect 38660 6604 38712 6613
rect 39672 6672 39724 6724
rect 39488 6604 39540 6656
rect 3010 6502 3062 6554
rect 3074 6502 3126 6554
rect 3138 6502 3190 6554
rect 3202 6502 3254 6554
rect 3266 6502 3318 6554
rect 9010 6502 9062 6554
rect 9074 6502 9126 6554
rect 9138 6502 9190 6554
rect 9202 6502 9254 6554
rect 9266 6502 9318 6554
rect 15010 6502 15062 6554
rect 15074 6502 15126 6554
rect 15138 6502 15190 6554
rect 15202 6502 15254 6554
rect 15266 6502 15318 6554
rect 21010 6502 21062 6554
rect 21074 6502 21126 6554
rect 21138 6502 21190 6554
rect 21202 6502 21254 6554
rect 21266 6502 21318 6554
rect 27010 6502 27062 6554
rect 27074 6502 27126 6554
rect 27138 6502 27190 6554
rect 27202 6502 27254 6554
rect 27266 6502 27318 6554
rect 33010 6502 33062 6554
rect 33074 6502 33126 6554
rect 33138 6502 33190 6554
rect 33202 6502 33254 6554
rect 33266 6502 33318 6554
rect 39010 6502 39062 6554
rect 39074 6502 39126 6554
rect 39138 6502 39190 6554
rect 39202 6502 39254 6554
rect 39266 6502 39318 6554
rect 1492 6400 1544 6452
rect 2872 6400 2924 6452
rect 3424 6400 3476 6452
rect 5356 6400 5408 6452
rect 6184 6400 6236 6452
rect 6460 6443 6512 6452
rect 6460 6409 6469 6443
rect 6469 6409 6503 6443
rect 6503 6409 6512 6443
rect 6460 6400 6512 6409
rect 7012 6400 7064 6452
rect 7104 6400 7156 6452
rect 7564 6443 7616 6452
rect 7564 6409 7573 6443
rect 7573 6409 7607 6443
rect 7607 6409 7616 6443
rect 7564 6400 7616 6409
rect 7748 6400 7800 6452
rect 1308 6332 1360 6384
rect 2412 6332 2464 6384
rect 3976 6332 4028 6384
rect 1860 6264 1912 6316
rect 4344 6332 4396 6384
rect 7472 6332 7524 6384
rect 4436 6264 4488 6316
rect 4620 6307 4672 6316
rect 4620 6273 4629 6307
rect 4629 6273 4663 6307
rect 4663 6273 4672 6307
rect 4620 6264 4672 6273
rect 5448 6264 5500 6316
rect 5908 6264 5960 6316
rect 2136 6239 2188 6248
rect 2136 6205 2145 6239
rect 2145 6205 2179 6239
rect 2179 6205 2188 6239
rect 2136 6196 2188 6205
rect 3148 6128 3200 6180
rect 2872 6060 2924 6112
rect 3332 6239 3384 6248
rect 3332 6205 3341 6239
rect 3341 6205 3375 6239
rect 3375 6205 3384 6239
rect 3332 6196 3384 6205
rect 6644 6307 6696 6316
rect 6644 6273 6653 6307
rect 6653 6273 6687 6307
rect 6687 6273 6696 6307
rect 6644 6264 6696 6273
rect 7104 6264 7156 6316
rect 7288 6264 7340 6316
rect 7564 6264 7616 6316
rect 8116 6332 8168 6384
rect 8760 6400 8812 6452
rect 9036 6332 9088 6384
rect 3976 6128 4028 6180
rect 4528 6128 4580 6180
rect 4620 6128 4672 6180
rect 7656 6196 7708 6248
rect 8116 6196 8168 6248
rect 8668 6307 8720 6316
rect 8668 6273 8677 6307
rect 8677 6273 8711 6307
rect 8711 6273 8720 6307
rect 8668 6264 8720 6273
rect 8760 6307 8812 6316
rect 8760 6273 8769 6307
rect 8769 6273 8803 6307
rect 8803 6273 8812 6307
rect 8760 6264 8812 6273
rect 3608 6060 3660 6112
rect 3700 6060 3752 6112
rect 4712 6060 4764 6112
rect 5540 6060 5592 6112
rect 6460 6128 6512 6180
rect 7748 6128 7800 6180
rect 8024 6128 8076 6180
rect 9128 6264 9180 6316
rect 10508 6400 10560 6452
rect 10692 6400 10744 6452
rect 10876 6400 10928 6452
rect 9496 6375 9548 6384
rect 9496 6341 9505 6375
rect 9505 6341 9539 6375
rect 9539 6341 9548 6375
rect 9496 6332 9548 6341
rect 10416 6332 10468 6384
rect 9588 6264 9640 6316
rect 10140 6307 10192 6316
rect 10140 6273 10149 6307
rect 10149 6273 10183 6307
rect 10183 6273 10192 6307
rect 12164 6400 12216 6452
rect 18236 6400 18288 6452
rect 18328 6400 18380 6452
rect 25964 6400 26016 6452
rect 26424 6400 26476 6452
rect 26792 6443 26844 6452
rect 26792 6409 26801 6443
rect 26801 6409 26835 6443
rect 26835 6409 26844 6443
rect 26792 6400 26844 6409
rect 26976 6400 27028 6452
rect 27528 6400 27580 6452
rect 10140 6264 10192 6273
rect 9404 6196 9456 6248
rect 11244 6264 11296 6316
rect 11888 6307 11940 6316
rect 11888 6273 11922 6307
rect 11922 6273 11940 6307
rect 11888 6264 11940 6273
rect 12716 6332 12768 6384
rect 13544 6332 13596 6384
rect 13820 6332 13872 6384
rect 13912 6332 13964 6384
rect 15476 6332 15528 6384
rect 11428 6196 11480 6248
rect 14464 6264 14516 6316
rect 15108 6264 15160 6316
rect 15568 6264 15620 6316
rect 16396 6375 16448 6384
rect 16396 6341 16405 6375
rect 16405 6341 16439 6375
rect 16439 6341 16448 6375
rect 16396 6332 16448 6341
rect 17224 6332 17276 6384
rect 17408 6332 17460 6384
rect 17868 6332 17920 6384
rect 21364 6332 21416 6384
rect 22192 6375 22244 6384
rect 22192 6341 22201 6375
rect 22201 6341 22235 6375
rect 22235 6341 22244 6375
rect 22192 6332 22244 6341
rect 10692 6128 10744 6180
rect 10232 6060 10284 6112
rect 10324 6103 10376 6112
rect 10324 6069 10333 6103
rect 10333 6069 10367 6103
rect 10367 6069 10376 6103
rect 10324 6060 10376 6069
rect 10876 6103 10928 6112
rect 10876 6069 10885 6103
rect 10885 6069 10919 6103
rect 10919 6069 10928 6103
rect 10876 6060 10928 6069
rect 11336 6103 11388 6112
rect 11336 6069 11345 6103
rect 11345 6069 11379 6103
rect 11379 6069 11388 6103
rect 11336 6060 11388 6069
rect 14188 6196 14240 6248
rect 13820 6128 13872 6180
rect 14924 6128 14976 6180
rect 11980 6060 12032 6112
rect 12716 6060 12768 6112
rect 13084 6103 13136 6112
rect 13084 6069 13093 6103
rect 13093 6069 13127 6103
rect 13127 6069 13136 6103
rect 13084 6060 13136 6069
rect 13544 6060 13596 6112
rect 14556 6060 14608 6112
rect 16580 6264 16632 6316
rect 16856 6307 16908 6316
rect 16856 6273 16865 6307
rect 16865 6273 16899 6307
rect 16899 6273 16908 6307
rect 16856 6264 16908 6273
rect 16948 6264 17000 6316
rect 18604 6307 18656 6316
rect 18604 6273 18613 6307
rect 18613 6273 18647 6307
rect 18647 6273 18656 6307
rect 18604 6264 18656 6273
rect 16396 6196 16448 6248
rect 17040 6239 17092 6248
rect 17040 6205 17049 6239
rect 17049 6205 17083 6239
rect 17083 6205 17092 6239
rect 17040 6196 17092 6205
rect 17408 6239 17460 6248
rect 17408 6205 17417 6239
rect 17417 6205 17451 6239
rect 17451 6205 17460 6239
rect 17408 6196 17460 6205
rect 18144 6196 18196 6248
rect 18420 6196 18472 6248
rect 19248 6264 19300 6316
rect 20628 6264 20680 6316
rect 21548 6307 21600 6316
rect 21548 6273 21557 6307
rect 21557 6273 21591 6307
rect 21591 6273 21600 6307
rect 21548 6264 21600 6273
rect 22100 6264 22152 6316
rect 22652 6332 22704 6384
rect 25504 6332 25556 6384
rect 25780 6332 25832 6384
rect 22468 6264 22520 6316
rect 23112 6264 23164 6316
rect 23480 6264 23532 6316
rect 24676 6264 24728 6316
rect 25228 6307 25280 6316
rect 25228 6273 25237 6307
rect 25237 6273 25271 6307
rect 25271 6273 25280 6307
rect 25228 6264 25280 6273
rect 25688 6307 25740 6316
rect 25688 6273 25697 6307
rect 25697 6273 25731 6307
rect 25731 6273 25740 6307
rect 25688 6264 25740 6273
rect 25872 6264 25924 6316
rect 26240 6264 26292 6316
rect 26608 6307 26660 6316
rect 26608 6273 26617 6307
rect 26617 6273 26651 6307
rect 26651 6273 26660 6307
rect 26608 6264 26660 6273
rect 23388 6196 23440 6248
rect 23572 6196 23624 6248
rect 27620 6307 27672 6316
rect 27620 6273 27629 6307
rect 27629 6273 27663 6307
rect 27663 6273 27672 6307
rect 27620 6264 27672 6273
rect 27528 6196 27580 6248
rect 29736 6400 29788 6452
rect 31392 6443 31444 6452
rect 31392 6409 31401 6443
rect 31401 6409 31435 6443
rect 31435 6409 31444 6443
rect 31392 6400 31444 6409
rect 31576 6400 31628 6452
rect 31944 6400 31996 6452
rect 34060 6400 34112 6452
rect 34888 6400 34940 6452
rect 35532 6400 35584 6452
rect 36084 6443 36136 6452
rect 36084 6409 36093 6443
rect 36093 6409 36127 6443
rect 36127 6409 36136 6443
rect 36084 6400 36136 6409
rect 36912 6400 36964 6452
rect 38476 6400 38528 6452
rect 39396 6443 39448 6452
rect 39396 6409 39405 6443
rect 39405 6409 39439 6443
rect 39439 6409 39448 6443
rect 39396 6400 39448 6409
rect 28724 6264 28776 6316
rect 31116 6332 31168 6384
rect 36636 6332 36688 6384
rect 38844 6332 38896 6384
rect 30104 6264 30156 6316
rect 30288 6307 30340 6316
rect 30288 6273 30297 6307
rect 30297 6273 30331 6307
rect 30331 6273 30340 6307
rect 30288 6264 30340 6273
rect 30656 6307 30708 6316
rect 30656 6273 30665 6307
rect 30665 6273 30699 6307
rect 30699 6273 30708 6307
rect 30656 6264 30708 6273
rect 30012 6196 30064 6248
rect 31024 6264 31076 6316
rect 31760 6264 31812 6316
rect 34520 6264 34572 6316
rect 35348 6264 35400 6316
rect 35624 6264 35676 6316
rect 36176 6264 36228 6316
rect 37096 6264 37148 6316
rect 32312 6239 32364 6248
rect 32312 6205 32321 6239
rect 32321 6205 32355 6239
rect 32355 6205 32364 6239
rect 32312 6196 32364 6205
rect 16948 6128 17000 6180
rect 16304 6060 16356 6112
rect 17500 6060 17552 6112
rect 17684 6060 17736 6112
rect 18420 6103 18472 6112
rect 18420 6069 18429 6103
rect 18429 6069 18463 6103
rect 18463 6069 18472 6103
rect 18420 6060 18472 6069
rect 18512 6060 18564 6112
rect 19064 6128 19116 6180
rect 22284 6128 22336 6180
rect 22560 6171 22612 6180
rect 22560 6137 22569 6171
rect 22569 6137 22603 6171
rect 22603 6137 22612 6171
rect 22560 6128 22612 6137
rect 19248 6103 19300 6112
rect 19248 6069 19257 6103
rect 19257 6069 19291 6103
rect 19291 6069 19300 6103
rect 19248 6060 19300 6069
rect 19432 6060 19484 6112
rect 21456 6060 21508 6112
rect 23480 6128 23532 6180
rect 23756 6128 23808 6180
rect 22928 6103 22980 6112
rect 22928 6069 22937 6103
rect 22937 6069 22971 6103
rect 22971 6069 22980 6103
rect 22928 6060 22980 6069
rect 23020 6060 23072 6112
rect 24952 6060 25004 6112
rect 25044 6103 25096 6112
rect 25044 6069 25053 6103
rect 25053 6069 25087 6103
rect 25087 6069 25096 6103
rect 25044 6060 25096 6069
rect 25504 6103 25556 6112
rect 25504 6069 25513 6103
rect 25513 6069 25547 6103
rect 25547 6069 25556 6103
rect 25504 6060 25556 6069
rect 25688 6060 25740 6112
rect 25872 6060 25924 6112
rect 26976 6060 27028 6112
rect 27160 6103 27212 6112
rect 27160 6069 27169 6103
rect 27169 6069 27203 6103
rect 27203 6069 27212 6103
rect 27160 6060 27212 6069
rect 28632 6060 28684 6112
rect 29552 6060 29604 6112
rect 31300 6060 31352 6112
rect 32036 6060 32088 6112
rect 32312 6060 32364 6112
rect 34888 6196 34940 6248
rect 36268 6196 36320 6248
rect 38476 6196 38528 6248
rect 37556 6128 37608 6180
rect 33416 6103 33468 6112
rect 33416 6069 33425 6103
rect 33425 6069 33459 6103
rect 33459 6069 33468 6103
rect 33416 6060 33468 6069
rect 35256 6060 35308 6112
rect 38844 6103 38896 6112
rect 38844 6069 38853 6103
rect 38853 6069 38887 6103
rect 38887 6069 38896 6103
rect 38844 6060 38896 6069
rect 1950 5958 2002 6010
rect 2014 5958 2066 6010
rect 2078 5958 2130 6010
rect 2142 5958 2194 6010
rect 2206 5958 2258 6010
rect 7950 5958 8002 6010
rect 8014 5958 8066 6010
rect 8078 5958 8130 6010
rect 8142 5958 8194 6010
rect 8206 5958 8258 6010
rect 13950 5958 14002 6010
rect 14014 5958 14066 6010
rect 14078 5958 14130 6010
rect 14142 5958 14194 6010
rect 14206 5958 14258 6010
rect 19950 5958 20002 6010
rect 20014 5958 20066 6010
rect 20078 5958 20130 6010
rect 20142 5958 20194 6010
rect 20206 5958 20258 6010
rect 25950 5958 26002 6010
rect 26014 5958 26066 6010
rect 26078 5958 26130 6010
rect 26142 5958 26194 6010
rect 26206 5958 26258 6010
rect 31950 5958 32002 6010
rect 32014 5958 32066 6010
rect 32078 5958 32130 6010
rect 32142 5958 32194 6010
rect 32206 5958 32258 6010
rect 37950 5958 38002 6010
rect 38014 5958 38066 6010
rect 38078 5958 38130 6010
rect 38142 5958 38194 6010
rect 38206 5958 38258 6010
rect 2504 5856 2556 5908
rect 3332 5856 3384 5908
rect 4160 5856 4212 5908
rect 4620 5856 4672 5908
rect 2688 5788 2740 5840
rect 5080 5788 5132 5840
rect 6736 5856 6788 5908
rect 7380 5856 7432 5908
rect 7840 5856 7892 5908
rect 8392 5856 8444 5908
rect 4712 5720 4764 5772
rect 5448 5720 5500 5772
rect 5540 5763 5592 5772
rect 5540 5729 5549 5763
rect 5549 5729 5583 5763
rect 5583 5729 5592 5763
rect 5540 5720 5592 5729
rect 7196 5788 7248 5840
rect 1032 5652 1084 5704
rect 2320 5695 2372 5704
rect 2320 5661 2329 5695
rect 2329 5661 2363 5695
rect 2363 5661 2372 5695
rect 2320 5652 2372 5661
rect 2504 5695 2556 5704
rect 2504 5661 2513 5695
rect 2513 5661 2547 5695
rect 2547 5661 2556 5695
rect 2504 5652 2556 5661
rect 388 5584 440 5636
rect 3516 5584 3568 5636
rect 3976 5652 4028 5704
rect 4528 5652 4580 5704
rect 5356 5652 5408 5704
rect 5908 5652 5960 5704
rect 7288 5652 7340 5704
rect 4620 5584 4672 5636
rect 2504 5516 2556 5568
rect 5816 5584 5868 5636
rect 7472 5584 7524 5636
rect 9312 5856 9364 5908
rect 10416 5899 10468 5908
rect 10416 5865 10425 5899
rect 10425 5865 10459 5899
rect 10459 5865 10468 5899
rect 10416 5856 10468 5865
rect 10692 5856 10744 5908
rect 13820 5856 13872 5908
rect 14280 5856 14332 5908
rect 15108 5856 15160 5908
rect 8852 5720 8904 5772
rect 10876 5788 10928 5840
rect 14464 5788 14516 5840
rect 15568 5899 15620 5908
rect 15568 5865 15577 5899
rect 15577 5865 15611 5899
rect 15611 5865 15620 5899
rect 15568 5856 15620 5865
rect 15936 5856 15988 5908
rect 16212 5788 16264 5840
rect 16304 5788 16356 5840
rect 17316 5899 17368 5908
rect 17316 5865 17325 5899
rect 17325 5865 17359 5899
rect 17359 5865 17368 5899
rect 17316 5856 17368 5865
rect 17592 5856 17644 5908
rect 9680 5652 9732 5704
rect 13084 5720 13136 5772
rect 11428 5695 11480 5704
rect 11428 5661 11437 5695
rect 11437 5661 11471 5695
rect 11471 5661 11480 5695
rect 11428 5652 11480 5661
rect 11612 5695 11664 5704
rect 11612 5661 11621 5695
rect 11621 5661 11655 5695
rect 11655 5661 11664 5695
rect 11612 5652 11664 5661
rect 8668 5584 8720 5636
rect 10324 5584 10376 5636
rect 11336 5584 11388 5636
rect 12256 5652 12308 5704
rect 13636 5652 13688 5704
rect 15476 5695 15528 5704
rect 15476 5661 15485 5695
rect 15485 5661 15519 5695
rect 15519 5661 15528 5695
rect 15476 5652 15528 5661
rect 15660 5652 15712 5704
rect 12072 5627 12124 5636
rect 12072 5593 12081 5627
rect 12081 5593 12115 5627
rect 12115 5593 12124 5627
rect 12072 5584 12124 5593
rect 12164 5627 12216 5636
rect 12164 5593 12173 5627
rect 12173 5593 12207 5627
rect 12207 5593 12216 5627
rect 12164 5584 12216 5593
rect 5172 5516 5224 5568
rect 5356 5559 5408 5568
rect 5356 5525 5365 5559
rect 5365 5525 5399 5559
rect 5399 5525 5408 5559
rect 5356 5516 5408 5525
rect 6552 5516 6604 5568
rect 8300 5516 8352 5568
rect 11428 5516 11480 5568
rect 15108 5584 15160 5636
rect 16028 5695 16080 5704
rect 16028 5661 16037 5695
rect 16037 5661 16071 5695
rect 16071 5661 16080 5695
rect 16028 5652 16080 5661
rect 16212 5695 16264 5704
rect 16212 5661 16221 5695
rect 16221 5661 16255 5695
rect 16255 5661 16264 5695
rect 16212 5652 16264 5661
rect 16580 5695 16632 5704
rect 16580 5661 16589 5695
rect 16589 5661 16623 5695
rect 16623 5661 16632 5695
rect 16580 5652 16632 5661
rect 17776 5652 17828 5704
rect 16672 5584 16724 5636
rect 18512 5788 18564 5840
rect 18420 5720 18472 5772
rect 18880 5720 18932 5772
rect 20720 5856 20772 5908
rect 24492 5856 24544 5908
rect 26516 5856 26568 5908
rect 27160 5856 27212 5908
rect 27896 5856 27948 5908
rect 28264 5856 28316 5908
rect 29552 5856 29604 5908
rect 23112 5831 23164 5840
rect 23112 5797 23121 5831
rect 23121 5797 23155 5831
rect 23155 5797 23164 5831
rect 23112 5788 23164 5797
rect 24032 5831 24084 5840
rect 24032 5797 24041 5831
rect 24041 5797 24075 5831
rect 24075 5797 24084 5831
rect 24032 5788 24084 5797
rect 24216 5788 24268 5840
rect 28080 5788 28132 5840
rect 29184 5788 29236 5840
rect 30196 5788 30248 5840
rect 31208 5899 31260 5908
rect 31208 5865 31217 5899
rect 31217 5865 31251 5899
rect 31251 5865 31260 5899
rect 31208 5856 31260 5865
rect 36636 5856 36688 5908
rect 36820 5856 36872 5908
rect 37832 5856 37884 5908
rect 34152 5788 34204 5840
rect 36360 5788 36412 5840
rect 39396 5831 39448 5840
rect 39396 5797 39405 5831
rect 39405 5797 39439 5831
rect 39439 5797 39448 5831
rect 39396 5788 39448 5797
rect 18328 5652 18380 5704
rect 18788 5695 18840 5704
rect 18788 5661 18797 5695
rect 18797 5661 18831 5695
rect 18831 5661 18840 5695
rect 18788 5652 18840 5661
rect 19340 5652 19392 5704
rect 22008 5720 22060 5772
rect 22284 5763 22336 5772
rect 22284 5729 22318 5763
rect 22318 5729 22336 5763
rect 22284 5720 22336 5729
rect 12348 5516 12400 5568
rect 16948 5516 17000 5568
rect 17132 5516 17184 5568
rect 17776 5516 17828 5568
rect 18328 5516 18380 5568
rect 18512 5559 18564 5568
rect 18512 5525 18521 5559
rect 18521 5525 18555 5559
rect 18555 5525 18564 5559
rect 18512 5516 18564 5525
rect 19708 5584 19760 5636
rect 21640 5652 21692 5704
rect 22652 5720 22704 5772
rect 24584 5720 24636 5772
rect 24952 5763 25004 5772
rect 24952 5729 24961 5763
rect 24961 5729 24995 5763
rect 24995 5729 25004 5763
rect 24952 5720 25004 5729
rect 27436 5720 27488 5772
rect 29276 5720 29328 5772
rect 22468 5695 22520 5704
rect 22468 5661 22477 5695
rect 22477 5661 22511 5695
rect 22511 5661 22520 5695
rect 22468 5652 22520 5661
rect 23112 5652 23164 5704
rect 24400 5652 24452 5704
rect 24768 5695 24820 5704
rect 24768 5661 24777 5695
rect 24777 5661 24811 5695
rect 24811 5661 24820 5695
rect 24768 5652 24820 5661
rect 25872 5652 25924 5704
rect 26332 5652 26384 5704
rect 21364 5584 21416 5636
rect 18788 5516 18840 5568
rect 19064 5516 19116 5568
rect 21456 5516 21508 5568
rect 22008 5516 22060 5568
rect 23756 5584 23808 5636
rect 23940 5584 23992 5636
rect 23204 5559 23256 5568
rect 23204 5525 23213 5559
rect 23213 5525 23247 5559
rect 23247 5525 23256 5559
rect 23204 5516 23256 5525
rect 23572 5516 23624 5568
rect 24216 5516 24268 5568
rect 24400 5559 24452 5568
rect 24400 5525 24409 5559
rect 24409 5525 24443 5559
rect 24443 5525 24452 5559
rect 24400 5516 24452 5525
rect 24860 5516 24912 5568
rect 26424 5516 26476 5568
rect 28264 5584 28316 5636
rect 27344 5516 27396 5568
rect 27620 5559 27672 5568
rect 27620 5525 27629 5559
rect 27629 5525 27663 5559
rect 27663 5525 27672 5559
rect 27620 5516 27672 5525
rect 28632 5652 28684 5704
rect 28724 5695 28776 5704
rect 28724 5661 28733 5695
rect 28733 5661 28767 5695
rect 28767 5661 28776 5695
rect 28724 5652 28776 5661
rect 29000 5695 29052 5704
rect 29000 5661 29009 5695
rect 29009 5661 29043 5695
rect 29043 5661 29052 5695
rect 29000 5652 29052 5661
rect 29092 5652 29144 5704
rect 32956 5720 33008 5772
rect 34612 5720 34664 5772
rect 34796 5763 34848 5772
rect 34796 5729 34805 5763
rect 34805 5729 34839 5763
rect 34839 5729 34848 5763
rect 34796 5720 34848 5729
rect 37280 5720 37332 5772
rect 30012 5652 30064 5704
rect 30380 5652 30432 5704
rect 30748 5652 30800 5704
rect 29644 5584 29696 5636
rect 30656 5584 30708 5636
rect 32036 5695 32088 5704
rect 32036 5661 32045 5695
rect 32045 5661 32079 5695
rect 32079 5661 32088 5695
rect 32036 5652 32088 5661
rect 32220 5652 32272 5704
rect 33416 5695 33468 5704
rect 33416 5661 33425 5695
rect 33425 5661 33459 5695
rect 33459 5661 33468 5695
rect 33416 5652 33468 5661
rect 34520 5652 34572 5704
rect 35532 5652 35584 5704
rect 29000 5516 29052 5568
rect 29552 5559 29604 5568
rect 29552 5525 29561 5559
rect 29561 5525 29595 5559
rect 29595 5525 29604 5559
rect 29552 5516 29604 5525
rect 32956 5516 33008 5568
rect 33232 5559 33284 5568
rect 33232 5525 33241 5559
rect 33241 5525 33275 5559
rect 33275 5525 33284 5559
rect 33232 5516 33284 5525
rect 34796 5516 34848 5568
rect 35532 5516 35584 5568
rect 37280 5584 37332 5636
rect 37556 5584 37608 5636
rect 38568 5652 38620 5704
rect 39212 5695 39264 5704
rect 39212 5661 39221 5695
rect 39221 5661 39255 5695
rect 39255 5661 39264 5695
rect 39212 5652 39264 5661
rect 39764 5584 39816 5636
rect 39948 5516 40000 5568
rect 3010 5414 3062 5466
rect 3074 5414 3126 5466
rect 3138 5414 3190 5466
rect 3202 5414 3254 5466
rect 3266 5414 3318 5466
rect 9010 5414 9062 5466
rect 9074 5414 9126 5466
rect 9138 5414 9190 5466
rect 9202 5414 9254 5466
rect 9266 5414 9318 5466
rect 15010 5414 15062 5466
rect 15074 5414 15126 5466
rect 15138 5414 15190 5466
rect 15202 5414 15254 5466
rect 15266 5414 15318 5466
rect 21010 5414 21062 5466
rect 21074 5414 21126 5466
rect 21138 5414 21190 5466
rect 21202 5414 21254 5466
rect 21266 5414 21318 5466
rect 27010 5414 27062 5466
rect 27074 5414 27126 5466
rect 27138 5414 27190 5466
rect 27202 5414 27254 5466
rect 27266 5414 27318 5466
rect 33010 5414 33062 5466
rect 33074 5414 33126 5466
rect 33138 5414 33190 5466
rect 33202 5414 33254 5466
rect 33266 5414 33318 5466
rect 39010 5414 39062 5466
rect 39074 5414 39126 5466
rect 39138 5414 39190 5466
rect 39202 5414 39254 5466
rect 39266 5414 39318 5466
rect 1492 5312 1544 5364
rect 1768 5312 1820 5364
rect 1216 5244 1268 5296
rect 2780 5312 2832 5364
rect 5908 5312 5960 5364
rect 6276 5312 6328 5364
rect 848 5176 900 5228
rect 3884 5244 3936 5296
rect 5356 5244 5408 5296
rect 6828 5312 6880 5364
rect 7012 5312 7064 5364
rect 8944 5312 8996 5364
rect 9680 5312 9732 5364
rect 940 5108 992 5160
rect 1768 5083 1820 5092
rect 1768 5049 1777 5083
rect 1777 5049 1811 5083
rect 1811 5049 1820 5083
rect 1768 5040 1820 5049
rect 3516 5176 3568 5228
rect 3608 5219 3660 5228
rect 3608 5185 3617 5219
rect 3617 5185 3651 5219
rect 3651 5185 3660 5219
rect 3608 5176 3660 5185
rect 6184 5219 6236 5228
rect 6184 5185 6193 5219
rect 6193 5185 6227 5219
rect 6227 5185 6236 5219
rect 6184 5176 6236 5185
rect 6276 5176 6328 5228
rect 7012 5176 7064 5228
rect 7840 5176 7892 5228
rect 9036 5176 9088 5228
rect 9128 5176 9180 5228
rect 9864 5176 9916 5228
rect 8484 5151 8536 5160
rect 112 4972 164 5024
rect 2780 5083 2832 5092
rect 2780 5049 2789 5083
rect 2789 5049 2823 5083
rect 2823 5049 2832 5083
rect 2780 5040 2832 5049
rect 8484 5117 8493 5151
rect 8493 5117 8527 5151
rect 8527 5117 8536 5151
rect 8484 5108 8536 5117
rect 10692 5244 10744 5296
rect 11244 5244 11296 5296
rect 10324 5219 10376 5228
rect 10324 5185 10333 5219
rect 10333 5185 10367 5219
rect 10367 5185 10376 5219
rect 10324 5176 10376 5185
rect 10416 5219 10468 5228
rect 10416 5185 10425 5219
rect 10425 5185 10459 5219
rect 10459 5185 10468 5219
rect 10416 5176 10468 5185
rect 11428 5176 11480 5228
rect 11796 5219 11848 5228
rect 11796 5185 11805 5219
rect 11805 5185 11839 5219
rect 11839 5185 11848 5219
rect 11796 5176 11848 5185
rect 13360 5244 13412 5296
rect 11980 5176 12032 5228
rect 14740 5176 14792 5228
rect 15476 5244 15528 5296
rect 15660 5287 15712 5296
rect 15660 5253 15678 5287
rect 15678 5253 15712 5287
rect 15660 5244 15712 5253
rect 16212 5355 16264 5364
rect 16212 5321 16221 5355
rect 16221 5321 16255 5355
rect 16255 5321 16264 5355
rect 16212 5312 16264 5321
rect 17408 5244 17460 5296
rect 17592 5244 17644 5296
rect 18328 5312 18380 5364
rect 18696 5312 18748 5364
rect 19432 5312 19484 5364
rect 21180 5244 21232 5296
rect 5356 5040 5408 5092
rect 6368 5040 6420 5092
rect 3424 4972 3476 5024
rect 4620 5015 4672 5024
rect 4620 4981 4629 5015
rect 4629 4981 4663 5015
rect 4663 4981 4672 5015
rect 4620 4972 4672 4981
rect 5540 4972 5592 5024
rect 5816 4972 5868 5024
rect 6092 4972 6144 5024
rect 6736 5040 6788 5092
rect 7472 4972 7524 5024
rect 10232 5040 10284 5092
rect 9864 5015 9916 5024
rect 9864 4981 9873 5015
rect 9873 4981 9907 5015
rect 9907 4981 9916 5015
rect 9864 4972 9916 4981
rect 9956 5015 10008 5024
rect 9956 4981 9965 5015
rect 9965 4981 9999 5015
rect 9999 4981 10008 5015
rect 9956 4972 10008 4981
rect 11060 4972 11112 5024
rect 12900 5108 12952 5160
rect 14188 5108 14240 5160
rect 14832 5108 14884 5160
rect 12164 5083 12216 5092
rect 12164 5049 12173 5083
rect 12173 5049 12207 5083
rect 12207 5049 12216 5083
rect 12164 5040 12216 5049
rect 12624 5040 12676 5092
rect 14188 4972 14240 5024
rect 14464 4972 14516 5024
rect 16948 5219 17000 5228
rect 16948 5185 16957 5219
rect 16957 5185 16991 5219
rect 16991 5185 17000 5219
rect 16948 5176 17000 5185
rect 18972 5176 19024 5228
rect 19156 5219 19208 5228
rect 19156 5185 19165 5219
rect 19165 5185 19199 5219
rect 19199 5185 19208 5219
rect 19156 5176 19208 5185
rect 19616 5176 19668 5228
rect 20444 5176 20496 5228
rect 19432 5151 19484 5160
rect 19432 5117 19441 5151
rect 19441 5117 19475 5151
rect 19475 5117 19484 5151
rect 19432 5108 19484 5117
rect 20352 5108 20404 5160
rect 21548 5312 21600 5364
rect 23480 5355 23532 5364
rect 23480 5321 23489 5355
rect 23489 5321 23523 5355
rect 23523 5321 23532 5355
rect 23480 5312 23532 5321
rect 25320 5312 25372 5364
rect 26700 5312 26752 5364
rect 27160 5312 27212 5364
rect 27436 5312 27488 5364
rect 29092 5355 29144 5364
rect 29092 5321 29101 5355
rect 29101 5321 29135 5355
rect 29135 5321 29144 5355
rect 29092 5312 29144 5321
rect 29184 5355 29236 5364
rect 29184 5321 29193 5355
rect 29193 5321 29227 5355
rect 29227 5321 29236 5355
rect 29184 5312 29236 5321
rect 29644 5312 29696 5364
rect 30288 5312 30340 5364
rect 32404 5312 32456 5364
rect 36544 5312 36596 5364
rect 38384 5312 38436 5364
rect 38752 5312 38804 5364
rect 39396 5355 39448 5364
rect 39396 5321 39405 5355
rect 39405 5321 39439 5355
rect 39439 5321 39448 5355
rect 39396 5312 39448 5321
rect 21456 5244 21508 5296
rect 16212 4972 16264 5024
rect 19156 5040 19208 5092
rect 19340 5083 19392 5092
rect 19340 5049 19349 5083
rect 19349 5049 19383 5083
rect 19383 5049 19392 5083
rect 19340 5040 19392 5049
rect 22100 5108 22152 5160
rect 22376 5151 22428 5160
rect 22376 5117 22385 5151
rect 22385 5117 22419 5151
rect 22419 5117 22428 5151
rect 22376 5108 22428 5117
rect 23204 5244 23256 5296
rect 25504 5244 25556 5296
rect 23020 5219 23072 5228
rect 23020 5185 23029 5219
rect 23029 5185 23063 5219
rect 23063 5185 23072 5219
rect 23020 5176 23072 5185
rect 23388 5176 23440 5228
rect 23572 5219 23624 5228
rect 23572 5185 23581 5219
rect 23581 5185 23615 5219
rect 23615 5185 23624 5219
rect 23572 5176 23624 5185
rect 23756 5219 23808 5228
rect 23756 5185 23765 5219
rect 23765 5185 23799 5219
rect 23799 5185 23808 5219
rect 23756 5176 23808 5185
rect 25596 5176 25648 5228
rect 26332 5244 26384 5296
rect 26424 5244 26476 5296
rect 25964 5176 26016 5228
rect 27344 5176 27396 5228
rect 29460 5244 29512 5296
rect 27620 5176 27672 5228
rect 28356 5176 28408 5228
rect 30656 5176 30708 5228
rect 32036 5244 32088 5296
rect 37740 5176 37792 5228
rect 38200 5176 38252 5228
rect 38660 5176 38712 5228
rect 25688 5108 25740 5160
rect 26792 5108 26844 5160
rect 27068 5108 27120 5160
rect 28448 5151 28500 5160
rect 28448 5117 28457 5151
rect 28457 5117 28491 5151
rect 28491 5117 28500 5151
rect 28448 5108 28500 5117
rect 27896 5083 27948 5092
rect 27896 5049 27905 5083
rect 27905 5049 27939 5083
rect 27939 5049 27948 5083
rect 27896 5040 27948 5049
rect 19064 4972 19116 5024
rect 21272 4972 21324 5024
rect 21548 5015 21600 5024
rect 21548 4981 21557 5015
rect 21557 4981 21591 5015
rect 21591 4981 21600 5015
rect 21548 4972 21600 4981
rect 21640 4972 21692 5024
rect 21732 4972 21784 5024
rect 22284 4972 22336 5024
rect 23296 4972 23348 5024
rect 25228 4972 25280 5024
rect 26700 4972 26752 5024
rect 26792 5015 26844 5024
rect 26792 4981 26801 5015
rect 26801 4981 26835 5015
rect 26835 4981 26844 5015
rect 26792 4972 26844 4981
rect 27436 4972 27488 5024
rect 27528 4972 27580 5024
rect 28908 5040 28960 5092
rect 31208 5151 31260 5160
rect 31208 5117 31217 5151
rect 31217 5117 31251 5151
rect 31251 5117 31260 5151
rect 31208 5108 31260 5117
rect 33876 5108 33928 5160
rect 29828 4972 29880 5024
rect 33508 4972 33560 5024
rect 38200 4972 38252 5024
rect 38476 4972 38528 5024
rect 39028 5015 39080 5024
rect 39028 4981 39037 5015
rect 39037 4981 39071 5015
rect 39071 4981 39080 5015
rect 39028 4972 39080 4981
rect 1950 4870 2002 4922
rect 2014 4870 2066 4922
rect 2078 4870 2130 4922
rect 2142 4870 2194 4922
rect 2206 4870 2258 4922
rect 7950 4870 8002 4922
rect 8014 4870 8066 4922
rect 8078 4870 8130 4922
rect 8142 4870 8194 4922
rect 8206 4870 8258 4922
rect 13950 4870 14002 4922
rect 14014 4870 14066 4922
rect 14078 4870 14130 4922
rect 14142 4870 14194 4922
rect 14206 4870 14258 4922
rect 19950 4870 20002 4922
rect 20014 4870 20066 4922
rect 20078 4870 20130 4922
rect 20142 4870 20194 4922
rect 20206 4870 20258 4922
rect 25950 4870 26002 4922
rect 26014 4870 26066 4922
rect 26078 4870 26130 4922
rect 26142 4870 26194 4922
rect 26206 4870 26258 4922
rect 31950 4870 32002 4922
rect 32014 4870 32066 4922
rect 32078 4870 32130 4922
rect 32142 4870 32194 4922
rect 32206 4870 32258 4922
rect 37950 4870 38002 4922
rect 38014 4870 38066 4922
rect 38078 4870 38130 4922
rect 38142 4870 38194 4922
rect 38206 4870 38258 4922
rect 1492 4768 1544 4820
rect 2412 4811 2464 4820
rect 2412 4777 2421 4811
rect 2421 4777 2455 4811
rect 2455 4777 2464 4811
rect 2412 4768 2464 4777
rect 4804 4768 4856 4820
rect 1124 4700 1176 4752
rect 756 4632 808 4684
rect 2596 4564 2648 4616
rect 2872 4607 2924 4616
rect 2872 4573 2881 4607
rect 2881 4573 2915 4607
rect 2915 4573 2924 4607
rect 2872 4564 2924 4573
rect 3884 4632 3936 4684
rect 204 4428 256 4480
rect 2044 4539 2096 4548
rect 2044 4505 2053 4539
rect 2053 4505 2087 4539
rect 2087 4505 2096 4539
rect 2044 4496 2096 4505
rect 6460 4700 6512 4752
rect 6092 4632 6144 4684
rect 6368 4632 6420 4684
rect 7840 4768 7892 4820
rect 9404 4768 9456 4820
rect 9496 4768 9548 4820
rect 11888 4768 11940 4820
rect 13084 4768 13136 4820
rect 7748 4743 7800 4752
rect 7748 4709 7757 4743
rect 7757 4709 7791 4743
rect 7791 4709 7800 4743
rect 7748 4700 7800 4709
rect 8392 4700 8444 4752
rect 9036 4675 9088 4684
rect 5448 4607 5500 4616
rect 5448 4573 5457 4607
rect 5457 4573 5491 4607
rect 5491 4573 5500 4607
rect 5448 4564 5500 4573
rect 5724 4607 5776 4616
rect 5724 4573 5733 4607
rect 5733 4573 5767 4607
rect 5767 4573 5776 4607
rect 5724 4564 5776 4573
rect 6276 4564 6328 4616
rect 6644 4496 6696 4548
rect 2688 4471 2740 4480
rect 2688 4437 2697 4471
rect 2697 4437 2731 4471
rect 2731 4437 2740 4471
rect 2688 4428 2740 4437
rect 4068 4428 4120 4480
rect 5356 4428 5408 4480
rect 6828 4428 6880 4480
rect 8116 4564 8168 4616
rect 9036 4641 9045 4675
rect 9045 4641 9079 4675
rect 9079 4641 9088 4675
rect 9036 4632 9088 4641
rect 9312 4632 9364 4684
rect 9496 4675 9548 4684
rect 9496 4641 9505 4675
rect 9505 4641 9539 4675
rect 9539 4641 9548 4675
rect 9496 4632 9548 4641
rect 10784 4632 10836 4684
rect 11336 4743 11388 4752
rect 11336 4709 11345 4743
rect 11345 4709 11379 4743
rect 11379 4709 11388 4743
rect 11336 4700 11388 4709
rect 11520 4700 11572 4752
rect 12624 4700 12676 4752
rect 13360 4700 13412 4752
rect 13268 4675 13320 4684
rect 13268 4641 13277 4675
rect 13277 4641 13311 4675
rect 13311 4641 13320 4675
rect 13268 4632 13320 4641
rect 8576 4428 8628 4480
rect 11520 4564 11572 4616
rect 12440 4564 12492 4616
rect 14464 4700 14516 4752
rect 14924 4768 14976 4820
rect 15476 4768 15528 4820
rect 16672 4768 16724 4820
rect 17132 4811 17184 4820
rect 17132 4777 17141 4811
rect 17141 4777 17175 4811
rect 17175 4777 17184 4811
rect 17132 4768 17184 4777
rect 14188 4564 14240 4616
rect 14372 4564 14424 4616
rect 14740 4675 14792 4684
rect 14740 4641 14749 4675
rect 14749 4641 14783 4675
rect 14783 4641 14792 4675
rect 14740 4632 14792 4641
rect 15752 4632 15804 4684
rect 9956 4496 10008 4548
rect 11060 4496 11112 4548
rect 12164 4496 12216 4548
rect 13360 4496 13412 4548
rect 16396 4564 16448 4616
rect 16948 4632 17000 4684
rect 18052 4700 18104 4752
rect 19248 4700 19300 4752
rect 20904 4700 20956 4752
rect 16672 4607 16724 4616
rect 16672 4573 16681 4607
rect 16681 4573 16715 4607
rect 16715 4573 16724 4607
rect 16672 4564 16724 4573
rect 17040 4607 17092 4616
rect 17040 4573 17049 4607
rect 17049 4573 17083 4607
rect 17083 4573 17092 4607
rect 17040 4564 17092 4573
rect 19432 4632 19484 4684
rect 20628 4632 20680 4684
rect 21456 4768 21508 4820
rect 23112 4768 23164 4820
rect 23572 4768 23624 4820
rect 22928 4700 22980 4752
rect 23756 4700 23808 4752
rect 27160 4768 27212 4820
rect 18236 4564 18288 4616
rect 18696 4564 18748 4616
rect 20444 4564 20496 4616
rect 20812 4607 20864 4616
rect 20812 4573 20821 4607
rect 20821 4573 20855 4607
rect 20855 4573 20864 4607
rect 20812 4564 20864 4573
rect 21548 4675 21600 4684
rect 21548 4641 21557 4675
rect 21557 4641 21591 4675
rect 21591 4641 21600 4675
rect 21548 4632 21600 4641
rect 21640 4632 21692 4684
rect 21916 4632 21968 4684
rect 22284 4632 22336 4684
rect 23940 4632 23992 4684
rect 23572 4564 23624 4616
rect 24768 4564 24820 4616
rect 24860 4607 24912 4616
rect 24860 4573 24869 4607
rect 24869 4573 24903 4607
rect 24903 4573 24912 4607
rect 24860 4564 24912 4573
rect 27068 4700 27120 4752
rect 27620 4700 27672 4752
rect 25228 4632 25280 4684
rect 10692 4428 10744 4480
rect 12532 4428 12584 4480
rect 14832 4428 14884 4480
rect 15384 4428 15436 4480
rect 15568 4428 15620 4480
rect 16304 4428 16356 4480
rect 16396 4428 16448 4480
rect 23296 4496 23348 4548
rect 25504 4496 25556 4548
rect 18328 4471 18380 4480
rect 18328 4437 18337 4471
rect 18337 4437 18371 4471
rect 18371 4437 18380 4471
rect 18328 4428 18380 4437
rect 20444 4428 20496 4480
rect 20536 4428 20588 4480
rect 20996 4428 21048 4480
rect 21548 4428 21600 4480
rect 24400 4471 24452 4480
rect 24400 4437 24409 4471
rect 24409 4437 24443 4471
rect 24443 4437 24452 4471
rect 24400 4428 24452 4437
rect 25320 4428 25372 4480
rect 26976 4632 27028 4684
rect 29000 4768 29052 4820
rect 30656 4768 30708 4820
rect 28908 4632 28960 4684
rect 26240 4607 26292 4616
rect 26240 4573 26249 4607
rect 26249 4573 26283 4607
rect 26283 4573 26292 4607
rect 26240 4564 26292 4573
rect 26608 4564 26660 4616
rect 27436 4564 27488 4616
rect 28264 4607 28316 4616
rect 28264 4573 28273 4607
rect 28273 4573 28307 4607
rect 28307 4573 28316 4607
rect 28264 4564 28316 4573
rect 28356 4607 28408 4616
rect 28356 4573 28390 4607
rect 28390 4573 28408 4607
rect 28356 4564 28408 4573
rect 28540 4607 28592 4616
rect 28540 4573 28549 4607
rect 28549 4573 28583 4607
rect 28583 4573 28592 4607
rect 28540 4564 28592 4573
rect 30380 4564 30432 4616
rect 26976 4496 27028 4548
rect 29736 4496 29788 4548
rect 31116 4564 31168 4616
rect 30656 4496 30708 4548
rect 31668 4632 31720 4684
rect 33600 4700 33652 4752
rect 35992 4811 36044 4820
rect 35992 4777 36001 4811
rect 36001 4777 36035 4811
rect 36035 4777 36044 4811
rect 35992 4768 36044 4777
rect 37004 4768 37056 4820
rect 37648 4768 37700 4820
rect 39396 4743 39448 4752
rect 39396 4709 39405 4743
rect 39405 4709 39439 4743
rect 39439 4709 39448 4743
rect 39396 4700 39448 4709
rect 32220 4564 32272 4616
rect 32404 4564 32456 4616
rect 32496 4607 32548 4616
rect 32496 4573 32505 4607
rect 32505 4573 32539 4607
rect 32539 4573 32548 4607
rect 32496 4564 32548 4573
rect 33508 4675 33560 4684
rect 33508 4641 33517 4675
rect 33517 4641 33551 4675
rect 33551 4641 33560 4675
rect 33508 4632 33560 4641
rect 35440 4607 35492 4616
rect 35440 4573 35449 4607
rect 35449 4573 35483 4607
rect 35483 4573 35492 4607
rect 35440 4564 35492 4573
rect 35532 4564 35584 4616
rect 32588 4496 32640 4548
rect 32404 4428 32456 4480
rect 32864 4428 32916 4480
rect 35348 4428 35400 4480
rect 36452 4496 36504 4548
rect 39856 4496 39908 4548
rect 39672 4428 39724 4480
rect 3010 4326 3062 4378
rect 3074 4326 3126 4378
rect 3138 4326 3190 4378
rect 3202 4326 3254 4378
rect 3266 4326 3318 4378
rect 9010 4326 9062 4378
rect 9074 4326 9126 4378
rect 9138 4326 9190 4378
rect 9202 4326 9254 4378
rect 9266 4326 9318 4378
rect 15010 4326 15062 4378
rect 15074 4326 15126 4378
rect 15138 4326 15190 4378
rect 15202 4326 15254 4378
rect 15266 4326 15318 4378
rect 21010 4326 21062 4378
rect 21074 4326 21126 4378
rect 21138 4326 21190 4378
rect 21202 4326 21254 4378
rect 21266 4326 21318 4378
rect 27010 4326 27062 4378
rect 27074 4326 27126 4378
rect 27138 4326 27190 4378
rect 27202 4326 27254 4378
rect 27266 4326 27318 4378
rect 33010 4326 33062 4378
rect 33074 4326 33126 4378
rect 33138 4326 33190 4378
rect 33202 4326 33254 4378
rect 33266 4326 33318 4378
rect 39010 4326 39062 4378
rect 39074 4326 39126 4378
rect 39138 4326 39190 4378
rect 39202 4326 39254 4378
rect 39266 4326 39318 4378
rect 2688 4156 2740 4208
rect 2872 4156 2924 4208
rect 3884 4224 3936 4276
rect 4344 4224 4396 4276
rect 6368 4224 6420 4276
rect 6920 4224 6972 4276
rect 7012 4224 7064 4276
rect 8576 4224 8628 4276
rect 7472 4156 7524 4208
rect 8300 4156 8352 4208
rect 296 4088 348 4140
rect 5172 4131 5224 4140
rect 5172 4097 5181 4131
rect 5181 4097 5215 4131
rect 5215 4097 5224 4131
rect 5172 4088 5224 4097
rect 5264 4131 5316 4140
rect 5264 4097 5273 4131
rect 5273 4097 5307 4131
rect 5307 4097 5316 4131
rect 5264 4088 5316 4097
rect 5356 4088 5408 4140
rect 5816 4131 5868 4140
rect 5816 4097 5825 4131
rect 5825 4097 5859 4131
rect 5859 4097 5868 4131
rect 5816 4088 5868 4097
rect 7012 4088 7064 4140
rect 8116 4088 8168 4140
rect 8944 4129 8996 4138
rect 756 4020 808 4072
rect 2688 4020 2740 4072
rect 3792 4020 3844 4072
rect 6092 4020 6144 4072
rect 6552 4063 6604 4072
rect 6552 4029 6561 4063
rect 6561 4029 6595 4063
rect 6595 4029 6604 4063
rect 6552 4020 6604 4029
rect 8392 4020 8444 4072
rect 8944 4095 8978 4129
rect 8978 4095 8996 4129
rect 8944 4086 8996 4095
rect 9956 4224 10008 4276
rect 10048 4224 10100 4276
rect 10416 4224 10468 4276
rect 12624 4224 12676 4276
rect 12900 4267 12952 4276
rect 12900 4233 12909 4267
rect 12909 4233 12943 4267
rect 12943 4233 12952 4267
rect 12900 4224 12952 4233
rect 13360 4224 13412 4276
rect 13452 4267 13504 4276
rect 13452 4233 13461 4267
rect 13461 4233 13495 4267
rect 13495 4233 13504 4267
rect 13452 4224 13504 4233
rect 14648 4224 14700 4276
rect 15384 4224 15436 4276
rect 9220 4131 9272 4140
rect 9220 4097 9229 4131
rect 9229 4097 9263 4131
rect 9263 4097 9272 4131
rect 9220 4088 9272 4097
rect 9772 4156 9824 4208
rect 9496 4129 9548 4140
rect 9496 4095 9505 4129
rect 9505 4095 9539 4129
rect 9539 4095 9548 4129
rect 9496 4088 9548 4095
rect 10048 4088 10100 4140
rect 10600 4088 10652 4140
rect 10784 4156 10836 4208
rect 11336 4156 11388 4208
rect 11428 4088 11480 4140
rect 11520 4131 11572 4140
rect 11520 4097 11529 4131
rect 11529 4097 11563 4131
rect 11563 4097 11572 4131
rect 11520 4088 11572 4097
rect 572 3884 624 3936
rect 2320 3884 2372 3936
rect 2504 3884 2556 3936
rect 4988 3995 5040 4004
rect 4988 3961 4997 3995
rect 4997 3961 5031 3995
rect 5031 3961 5040 3995
rect 4988 3952 5040 3961
rect 5172 3884 5224 3936
rect 5908 3952 5960 4004
rect 7656 3952 7708 4004
rect 8576 3995 8628 4004
rect 8576 3961 8585 3995
rect 8585 3961 8619 3995
rect 8619 3961 8628 3995
rect 8576 3952 8628 3961
rect 9036 3952 9088 4004
rect 9864 4020 9916 4072
rect 9220 3952 9272 4004
rect 9772 3952 9824 4004
rect 10784 4063 10836 4072
rect 10784 4029 10793 4063
rect 10793 4029 10827 4063
rect 10827 4029 10836 4063
rect 10784 4020 10836 4029
rect 13084 4131 13136 4140
rect 13084 4097 13093 4131
rect 13093 4097 13127 4131
rect 13127 4097 13136 4131
rect 13084 4088 13136 4097
rect 13268 4131 13320 4140
rect 13268 4097 13277 4131
rect 13277 4097 13311 4131
rect 13311 4097 13320 4131
rect 13268 4088 13320 4097
rect 13544 4131 13596 4140
rect 13544 4097 13553 4131
rect 13553 4097 13587 4131
rect 13587 4097 13596 4131
rect 13544 4088 13596 4097
rect 14372 4156 14424 4208
rect 14464 4199 14516 4208
rect 14464 4165 14473 4199
rect 14473 4165 14507 4199
rect 14507 4165 14516 4199
rect 14464 4156 14516 4165
rect 14832 4156 14884 4208
rect 15752 4224 15804 4276
rect 16396 4224 16448 4276
rect 16672 4224 16724 4276
rect 18236 4224 18288 4276
rect 22192 4267 22244 4276
rect 22192 4233 22201 4267
rect 22201 4233 22235 4267
rect 22235 4233 22244 4267
rect 22192 4224 22244 4233
rect 14096 4088 14148 4140
rect 13820 4063 13872 4072
rect 13820 4029 13829 4063
rect 13829 4029 13863 4063
rect 13863 4029 13872 4063
rect 13820 4020 13872 4029
rect 14832 4020 14884 4072
rect 16028 4131 16080 4140
rect 16028 4097 16037 4131
rect 16037 4097 16071 4131
rect 16071 4097 16080 4131
rect 16028 4088 16080 4097
rect 16764 4156 16816 4208
rect 17684 4156 17736 4208
rect 20720 4156 20772 4208
rect 23112 4224 23164 4276
rect 24584 4224 24636 4276
rect 25412 4267 25464 4276
rect 25412 4233 25421 4267
rect 25421 4233 25455 4267
rect 25455 4233 25464 4267
rect 25412 4224 25464 4233
rect 25504 4224 25556 4276
rect 29920 4224 29972 4276
rect 35808 4224 35860 4276
rect 23020 4156 23072 4208
rect 26240 4156 26292 4208
rect 26792 4156 26844 4208
rect 8944 3884 8996 3936
rect 9588 3927 9640 3936
rect 9588 3893 9597 3927
rect 9597 3893 9631 3927
rect 9631 3893 9640 3927
rect 9588 3884 9640 3893
rect 10968 3884 11020 3936
rect 11704 3884 11756 3936
rect 16120 4063 16172 4072
rect 16120 4029 16129 4063
rect 16129 4029 16163 4063
rect 16163 4029 16172 4063
rect 16120 4020 16172 4029
rect 16028 3952 16080 4004
rect 16488 4088 16540 4140
rect 18328 4088 18380 4140
rect 17960 4020 18012 4072
rect 18236 4020 18288 4072
rect 18880 4020 18932 4072
rect 18972 4063 19024 4072
rect 18972 4029 18981 4063
rect 18981 4029 19015 4063
rect 19015 4029 19024 4063
rect 18972 4020 19024 4029
rect 19524 4088 19576 4140
rect 20720 4020 20772 4072
rect 17868 3952 17920 4004
rect 20812 3952 20864 4004
rect 20996 4063 21048 4072
rect 20996 4029 21005 4063
rect 21005 4029 21039 4063
rect 21039 4029 21048 4063
rect 20996 4020 21048 4029
rect 22376 4020 22428 4072
rect 22468 4063 22520 4072
rect 22468 4029 22477 4063
rect 22477 4029 22511 4063
rect 22511 4029 22520 4063
rect 22468 4020 22520 4029
rect 23112 4063 23164 4072
rect 23112 4029 23121 4063
rect 23121 4029 23155 4063
rect 23155 4029 23164 4063
rect 23112 4020 23164 4029
rect 23296 4131 23348 4140
rect 23296 4097 23305 4131
rect 23305 4097 23339 4131
rect 23339 4097 23348 4131
rect 23296 4088 23348 4097
rect 23756 4088 23808 4140
rect 24400 4131 24452 4140
rect 24400 4097 24409 4131
rect 24409 4097 24443 4131
rect 24443 4097 24452 4131
rect 24400 4088 24452 4097
rect 24676 4088 24728 4140
rect 27896 4156 27948 4208
rect 27988 4199 28040 4208
rect 27988 4165 27997 4199
rect 27997 4165 28031 4199
rect 28031 4165 28040 4199
rect 27988 4156 28040 4165
rect 28356 4156 28408 4208
rect 28908 4199 28960 4208
rect 28908 4165 28917 4199
rect 28917 4165 28951 4199
rect 28951 4165 28960 4199
rect 28908 4156 28960 4165
rect 21364 3952 21416 4004
rect 16488 3927 16540 3936
rect 16488 3893 16497 3927
rect 16497 3893 16531 3927
rect 16531 3893 16540 3927
rect 16488 3884 16540 3893
rect 18328 3884 18380 3936
rect 18788 3884 18840 3936
rect 18880 3884 18932 3936
rect 22928 3884 22980 3936
rect 23664 3927 23716 3936
rect 23664 3893 23673 3927
rect 23673 3893 23707 3927
rect 23707 3893 23716 3927
rect 23664 3884 23716 3893
rect 25228 4063 25280 4072
rect 25228 4029 25237 4063
rect 25237 4029 25271 4063
rect 25271 4029 25280 4063
rect 25228 4020 25280 4029
rect 25320 4063 25372 4072
rect 25320 4029 25329 4063
rect 25329 4029 25363 4063
rect 25363 4029 25372 4063
rect 25320 4020 25372 4029
rect 26332 4020 26384 4072
rect 27344 4020 27396 4072
rect 27620 4088 27672 4140
rect 31668 4156 31720 4208
rect 34980 4156 35032 4208
rect 29920 4131 29972 4140
rect 29920 4097 29929 4131
rect 29929 4097 29963 4131
rect 29963 4097 29972 4131
rect 29920 4088 29972 4097
rect 30656 4131 30708 4140
rect 30656 4097 30665 4131
rect 30665 4097 30699 4131
rect 30699 4097 30708 4131
rect 30656 4088 30708 4097
rect 32404 4131 32456 4140
rect 32404 4097 32413 4131
rect 32413 4097 32447 4131
rect 32447 4097 32456 4131
rect 32404 4088 32456 4097
rect 32864 4088 32916 4140
rect 33416 4088 33468 4140
rect 34888 4131 34940 4140
rect 34888 4097 34897 4131
rect 34897 4097 34931 4131
rect 34931 4097 34940 4131
rect 34888 4088 34940 4097
rect 35440 4088 35492 4140
rect 36268 4088 36320 4140
rect 36636 4088 36688 4140
rect 38844 4131 38896 4140
rect 38844 4097 38853 4131
rect 38853 4097 38887 4131
rect 38887 4097 38896 4131
rect 38844 4088 38896 4097
rect 39580 4088 39632 4140
rect 26700 3952 26752 4004
rect 28264 4063 28316 4072
rect 28264 4029 28273 4063
rect 28273 4029 28307 4063
rect 28307 4029 28316 4063
rect 28264 4020 28316 4029
rect 28724 4020 28776 4072
rect 30104 4020 30156 4072
rect 31300 4020 31352 4072
rect 32588 4020 32640 4072
rect 33784 4020 33836 4072
rect 23940 3884 23992 3936
rect 25504 3884 25556 3936
rect 27344 3927 27396 3936
rect 27344 3893 27353 3927
rect 27353 3893 27387 3927
rect 27387 3893 27396 3927
rect 27344 3884 27396 3893
rect 28908 3952 28960 4004
rect 30656 3952 30708 4004
rect 31760 3952 31812 4004
rect 37464 3952 37516 4004
rect 39396 3995 39448 4004
rect 39396 3961 39405 3995
rect 39405 3961 39439 3995
rect 39439 3961 39448 3995
rect 39396 3952 39448 3961
rect 29736 3927 29788 3936
rect 29736 3893 29745 3927
rect 29745 3893 29779 3927
rect 29779 3893 29788 3927
rect 29736 3884 29788 3893
rect 30380 3884 30432 3936
rect 31116 3884 31168 3936
rect 32772 3927 32824 3936
rect 32772 3893 32781 3927
rect 32781 3893 32815 3927
rect 32815 3893 32824 3927
rect 32772 3884 32824 3893
rect 35992 3927 36044 3936
rect 35992 3893 36001 3927
rect 36001 3893 36035 3927
rect 36035 3893 36044 3927
rect 35992 3884 36044 3893
rect 39028 3927 39080 3936
rect 39028 3893 39037 3927
rect 39037 3893 39071 3927
rect 39071 3893 39080 3927
rect 39028 3884 39080 3893
rect 1950 3782 2002 3834
rect 2014 3782 2066 3834
rect 2078 3782 2130 3834
rect 2142 3782 2194 3834
rect 2206 3782 2258 3834
rect 7950 3782 8002 3834
rect 8014 3782 8066 3834
rect 8078 3782 8130 3834
rect 8142 3782 8194 3834
rect 8206 3782 8258 3834
rect 13950 3782 14002 3834
rect 14014 3782 14066 3834
rect 14078 3782 14130 3834
rect 14142 3782 14194 3834
rect 14206 3782 14258 3834
rect 19950 3782 20002 3834
rect 20014 3782 20066 3834
rect 20078 3782 20130 3834
rect 20142 3782 20194 3834
rect 20206 3782 20258 3834
rect 25950 3782 26002 3834
rect 26014 3782 26066 3834
rect 26078 3782 26130 3834
rect 26142 3782 26194 3834
rect 26206 3782 26258 3834
rect 31950 3782 32002 3834
rect 32014 3782 32066 3834
rect 32078 3782 32130 3834
rect 32142 3782 32194 3834
rect 32206 3782 32258 3834
rect 37950 3782 38002 3834
rect 38014 3782 38066 3834
rect 38078 3782 38130 3834
rect 38142 3782 38194 3834
rect 38206 3782 38258 3834
rect 1308 3680 1360 3732
rect 1124 3612 1176 3664
rect 388 3544 440 3596
rect 756 3476 808 3528
rect 1952 3655 2004 3664
rect 1952 3621 1961 3655
rect 1961 3621 1995 3655
rect 1995 3621 2004 3655
rect 1952 3612 2004 3621
rect 2320 3519 2372 3528
rect 2320 3485 2329 3519
rect 2329 3485 2363 3519
rect 2363 3485 2372 3519
rect 2320 3476 2372 3485
rect 2688 3612 2740 3664
rect 3792 3612 3844 3664
rect 4344 3612 4396 3664
rect 2688 3476 2740 3528
rect 5448 3723 5500 3732
rect 5448 3689 5457 3723
rect 5457 3689 5491 3723
rect 5491 3689 5500 3723
rect 5448 3680 5500 3689
rect 5816 3680 5868 3732
rect 5908 3680 5960 3732
rect 7196 3680 7248 3732
rect 6644 3612 6696 3664
rect 2780 3408 2832 3460
rect 1768 3340 1820 3392
rect 2872 3340 2924 3392
rect 3056 3383 3108 3392
rect 3056 3349 3065 3383
rect 3065 3349 3099 3383
rect 3099 3349 3108 3383
rect 3056 3340 3108 3349
rect 3700 3340 3752 3392
rect 3976 3383 4028 3392
rect 3976 3349 3985 3383
rect 3985 3349 4019 3383
rect 4019 3349 4028 3383
rect 3976 3340 4028 3349
rect 4712 3519 4764 3528
rect 4712 3485 4721 3519
rect 4721 3485 4755 3519
rect 4755 3485 4764 3519
rect 4712 3476 4764 3485
rect 5540 3519 5592 3528
rect 5540 3485 5549 3519
rect 5549 3485 5583 3519
rect 5583 3485 5592 3519
rect 5540 3476 5592 3485
rect 7196 3408 7248 3460
rect 7472 3544 7524 3596
rect 7656 3587 7708 3596
rect 7656 3553 7665 3587
rect 7665 3553 7699 3587
rect 7699 3553 7708 3587
rect 7656 3544 7708 3553
rect 8392 3680 8444 3732
rect 9036 3680 9088 3732
rect 10140 3680 10192 3732
rect 10784 3680 10836 3732
rect 11612 3723 11664 3732
rect 11612 3689 11621 3723
rect 11621 3689 11655 3723
rect 11655 3689 11664 3723
rect 11612 3680 11664 3689
rect 13176 3680 13228 3732
rect 13728 3680 13780 3732
rect 13268 3612 13320 3664
rect 14464 3723 14516 3732
rect 14464 3689 14473 3723
rect 14473 3689 14507 3723
rect 14507 3689 14516 3723
rect 14464 3680 14516 3689
rect 14740 3680 14792 3732
rect 20720 3680 20772 3732
rect 20996 3723 21048 3732
rect 20996 3689 21005 3723
rect 21005 3689 21039 3723
rect 21039 3689 21048 3723
rect 20996 3680 21048 3689
rect 16028 3612 16080 3664
rect 18236 3612 18288 3664
rect 19156 3612 19208 3664
rect 20352 3612 20404 3664
rect 23020 3680 23072 3732
rect 23112 3723 23164 3732
rect 23112 3689 23121 3723
rect 23121 3689 23155 3723
rect 23155 3689 23164 3723
rect 23112 3680 23164 3689
rect 24492 3655 24544 3664
rect 24492 3621 24501 3655
rect 24501 3621 24535 3655
rect 24535 3621 24544 3655
rect 24492 3612 24544 3621
rect 7380 3519 7432 3528
rect 7380 3485 7389 3519
rect 7389 3485 7423 3519
rect 7423 3485 7432 3519
rect 7380 3476 7432 3485
rect 8300 3476 8352 3528
rect 9220 3476 9272 3528
rect 9312 3519 9364 3528
rect 9312 3485 9321 3519
rect 9321 3485 9355 3519
rect 9355 3485 9364 3519
rect 9312 3476 9364 3485
rect 9680 3544 9732 3596
rect 11428 3544 11480 3596
rect 10600 3476 10652 3528
rect 11060 3476 11112 3528
rect 11888 3587 11940 3596
rect 11888 3553 11897 3587
rect 11897 3553 11931 3587
rect 11931 3553 11940 3587
rect 11888 3544 11940 3553
rect 13728 3544 13780 3596
rect 13084 3476 13136 3528
rect 13452 3476 13504 3528
rect 14464 3544 14516 3596
rect 14280 3476 14332 3528
rect 14740 3476 14792 3528
rect 14832 3519 14884 3528
rect 14832 3485 14841 3519
rect 14841 3485 14875 3519
rect 14875 3485 14884 3519
rect 14832 3476 14884 3485
rect 5356 3340 5408 3392
rect 7748 3340 7800 3392
rect 9312 3340 9364 3392
rect 9496 3340 9548 3392
rect 10232 3383 10284 3392
rect 10232 3349 10241 3383
rect 10241 3349 10275 3383
rect 10275 3349 10284 3383
rect 10232 3340 10284 3349
rect 10324 3340 10376 3392
rect 10784 3340 10836 3392
rect 11980 3340 12032 3392
rect 12164 3451 12216 3460
rect 12164 3417 12198 3451
rect 12198 3417 12216 3451
rect 12164 3408 12216 3417
rect 12348 3408 12400 3460
rect 12256 3340 12308 3392
rect 13636 3340 13688 3392
rect 14096 3408 14148 3460
rect 15384 3544 15436 3596
rect 17592 3544 17644 3596
rect 18972 3544 19024 3596
rect 19708 3544 19760 3596
rect 15108 3476 15160 3528
rect 15844 3519 15896 3528
rect 15844 3485 15853 3519
rect 15853 3485 15887 3519
rect 15887 3485 15896 3519
rect 15844 3476 15896 3485
rect 16948 3519 17000 3528
rect 16948 3485 16957 3519
rect 16957 3485 16991 3519
rect 16991 3485 17000 3519
rect 16948 3476 17000 3485
rect 17960 3519 18012 3528
rect 17960 3485 17969 3519
rect 17969 3485 18003 3519
rect 18003 3485 18012 3519
rect 17960 3476 18012 3485
rect 18236 3519 18288 3528
rect 18236 3485 18245 3519
rect 18245 3485 18279 3519
rect 18279 3485 18288 3519
rect 18236 3476 18288 3485
rect 18512 3519 18564 3528
rect 18512 3485 18521 3519
rect 18521 3485 18555 3519
rect 18555 3485 18564 3519
rect 18512 3476 18564 3485
rect 18788 3519 18840 3528
rect 18788 3485 18797 3519
rect 18797 3485 18831 3519
rect 18831 3485 18840 3519
rect 18788 3476 18840 3485
rect 19064 3519 19116 3528
rect 19064 3485 19073 3519
rect 19073 3485 19107 3519
rect 19107 3485 19116 3519
rect 19064 3476 19116 3485
rect 21364 3476 21416 3528
rect 21456 3519 21508 3528
rect 21456 3485 21465 3519
rect 21465 3485 21499 3519
rect 21499 3485 21508 3519
rect 21456 3476 21508 3485
rect 22100 3519 22152 3528
rect 22100 3485 22109 3519
rect 22109 3485 22143 3519
rect 22143 3485 22152 3519
rect 22100 3476 22152 3485
rect 23480 3519 23532 3528
rect 23480 3485 23489 3519
rect 23489 3485 23523 3519
rect 23523 3485 23532 3519
rect 23480 3476 23532 3485
rect 27528 3680 27580 3732
rect 28264 3680 28316 3732
rect 25412 3612 25464 3664
rect 25964 3612 26016 3664
rect 30656 3612 30708 3664
rect 38384 3680 38436 3732
rect 32864 3612 32916 3664
rect 38844 3612 38896 3664
rect 39396 3655 39448 3664
rect 39396 3621 39405 3655
rect 39405 3621 39439 3655
rect 39439 3621 39448 3655
rect 39396 3612 39448 3621
rect 25780 3587 25832 3596
rect 25780 3553 25789 3587
rect 25789 3553 25823 3587
rect 25823 3553 25832 3587
rect 25780 3544 25832 3553
rect 26516 3544 26568 3596
rect 26792 3587 26844 3596
rect 26792 3553 26801 3587
rect 26801 3553 26835 3587
rect 26835 3553 26844 3587
rect 26792 3544 26844 3553
rect 27712 3544 27764 3596
rect 31116 3544 31168 3596
rect 35256 3544 35308 3596
rect 25964 3519 26016 3528
rect 25964 3485 25973 3519
rect 25973 3485 26007 3519
rect 26007 3485 26016 3519
rect 25964 3476 26016 3485
rect 14004 3340 14056 3392
rect 15384 3340 15436 3392
rect 15476 3383 15528 3392
rect 15476 3349 15485 3383
rect 15485 3349 15519 3383
rect 15519 3349 15528 3383
rect 15476 3340 15528 3349
rect 15660 3383 15712 3392
rect 15660 3349 15669 3383
rect 15669 3349 15703 3383
rect 15703 3349 15712 3383
rect 15660 3340 15712 3349
rect 17132 3383 17184 3392
rect 17132 3349 17141 3383
rect 17141 3349 17175 3383
rect 17175 3349 17184 3383
rect 17132 3340 17184 3349
rect 17224 3383 17276 3392
rect 17224 3349 17233 3383
rect 17233 3349 17267 3383
rect 17267 3349 17276 3383
rect 17224 3340 17276 3349
rect 18236 3340 18288 3392
rect 18512 3340 18564 3392
rect 18696 3340 18748 3392
rect 19340 3340 19392 3392
rect 21640 3383 21692 3392
rect 21640 3349 21649 3383
rect 21649 3349 21683 3383
rect 21683 3349 21692 3383
rect 21640 3340 21692 3349
rect 22100 3340 22152 3392
rect 24216 3408 24268 3460
rect 25320 3408 25372 3460
rect 25412 3408 25464 3460
rect 26148 3408 26200 3460
rect 28172 3519 28224 3528
rect 28172 3485 28181 3519
rect 28181 3485 28215 3519
rect 28215 3485 28224 3519
rect 28172 3476 28224 3485
rect 31576 3476 31628 3528
rect 31944 3519 31996 3528
rect 31944 3485 31953 3519
rect 31953 3485 31987 3519
rect 31987 3485 31996 3519
rect 31944 3476 31996 3485
rect 32312 3476 32364 3528
rect 35992 3476 36044 3528
rect 37280 3544 37332 3596
rect 38476 3408 38528 3460
rect 28448 3340 28500 3392
rect 29644 3340 29696 3392
rect 30196 3340 30248 3392
rect 32220 3340 32272 3392
rect 32956 3340 33008 3392
rect 33968 3340 34020 3392
rect 34428 3340 34480 3392
rect 35808 3383 35860 3392
rect 35808 3349 35817 3383
rect 35817 3349 35851 3383
rect 35851 3349 35860 3383
rect 35808 3340 35860 3349
rect 39948 3340 40000 3392
rect 3010 3238 3062 3290
rect 3074 3238 3126 3290
rect 3138 3238 3190 3290
rect 3202 3238 3254 3290
rect 3266 3238 3318 3290
rect 9010 3238 9062 3290
rect 9074 3238 9126 3290
rect 9138 3238 9190 3290
rect 9202 3238 9254 3290
rect 9266 3238 9318 3290
rect 15010 3238 15062 3290
rect 15074 3238 15126 3290
rect 15138 3238 15190 3290
rect 15202 3238 15254 3290
rect 15266 3238 15318 3290
rect 21010 3238 21062 3290
rect 21074 3238 21126 3290
rect 21138 3238 21190 3290
rect 21202 3238 21254 3290
rect 21266 3238 21318 3290
rect 27010 3238 27062 3290
rect 27074 3238 27126 3290
rect 27138 3238 27190 3290
rect 27202 3238 27254 3290
rect 27266 3238 27318 3290
rect 33010 3238 33062 3290
rect 33074 3238 33126 3290
rect 33138 3238 33190 3290
rect 33202 3238 33254 3290
rect 33266 3238 33318 3290
rect 39010 3238 39062 3290
rect 39074 3238 39126 3290
rect 39138 3238 39190 3290
rect 39202 3238 39254 3290
rect 39266 3238 39318 3290
rect 1032 3068 1084 3120
rect 1952 3136 2004 3188
rect 4712 3111 4764 3120
rect 572 3000 624 3052
rect 4712 3077 4721 3111
rect 4721 3077 4755 3111
rect 4755 3077 4764 3111
rect 4712 3068 4764 3077
rect 6828 3136 6880 3188
rect 7196 3136 7248 3188
rect 7932 3136 7984 3188
rect 8484 3136 8536 3188
rect 9956 3179 10008 3188
rect 9956 3145 9965 3179
rect 9965 3145 9999 3179
rect 9999 3145 10008 3179
rect 9956 3136 10008 3145
rect 10140 3136 10192 3188
rect 10784 3136 10836 3188
rect 11796 3136 11848 3188
rect 11888 3136 11940 3188
rect 13636 3136 13688 3188
rect 13820 3136 13872 3188
rect 14004 3136 14056 3188
rect 14556 3136 14608 3188
rect 16028 3136 16080 3188
rect 23848 3136 23900 3188
rect 24124 3179 24176 3188
rect 24124 3145 24133 3179
rect 24133 3145 24167 3179
rect 24167 3145 24176 3179
rect 24124 3136 24176 3145
rect 25228 3179 25280 3188
rect 25228 3145 25237 3179
rect 25237 3145 25271 3179
rect 25271 3145 25280 3179
rect 25228 3136 25280 3145
rect 480 2932 532 2984
rect 2320 3043 2372 3052
rect 2320 3009 2329 3043
rect 2329 3009 2363 3043
rect 2363 3009 2372 3043
rect 2320 3000 2372 3009
rect 2596 3043 2648 3052
rect 2596 3009 2605 3043
rect 2605 3009 2639 3043
rect 2639 3009 2648 3043
rect 2596 3000 2648 3009
rect 2688 3000 2740 3052
rect 7472 3000 7524 3052
rect 7748 3000 7800 3052
rect 7932 3000 7984 3052
rect 8576 3000 8628 3052
rect 3608 2932 3660 2984
rect 3700 2932 3752 2984
rect 2412 2864 2464 2916
rect 4068 2864 4120 2916
rect 4896 2907 4948 2916
rect 4896 2873 4905 2907
rect 4905 2873 4939 2907
rect 4939 2873 4948 2907
rect 4896 2864 4948 2873
rect 6920 2975 6972 2984
rect 6920 2941 6929 2975
rect 6929 2941 6963 2975
rect 6963 2941 6972 2975
rect 6920 2932 6972 2941
rect 8484 2932 8536 2984
rect 9772 3043 9824 3052
rect 9772 3009 9781 3043
rect 9781 3009 9815 3043
rect 9815 3009 9824 3043
rect 9772 3000 9824 3009
rect 10508 3000 10560 3052
rect 10600 3043 10652 3052
rect 10600 3009 10609 3043
rect 10609 3009 10643 3043
rect 10643 3009 10652 3043
rect 10600 3000 10652 3009
rect 11612 3000 11664 3052
rect 11704 3043 11756 3052
rect 11704 3009 11713 3043
rect 11713 3009 11747 3043
rect 11747 3009 11756 3043
rect 11704 3000 11756 3009
rect 11796 3043 11848 3052
rect 11796 3009 11805 3043
rect 11805 3009 11839 3043
rect 11839 3009 11848 3043
rect 11796 3000 11848 3009
rect 11980 3000 12032 3052
rect 12900 3043 12952 3052
rect 12900 3009 12909 3043
rect 12909 3009 12943 3043
rect 12943 3009 12952 3043
rect 12900 3000 12952 3009
rect 13176 3043 13228 3052
rect 13176 3009 13185 3043
rect 13185 3009 13219 3043
rect 13219 3009 13228 3043
rect 13176 3000 13228 3009
rect 14648 3068 14700 3120
rect 16120 3068 16172 3120
rect 14832 3000 14884 3052
rect 17224 3068 17276 3120
rect 19432 3068 19484 3120
rect 10140 2932 10192 2984
rect 13544 2932 13596 2984
rect 13912 2932 13964 2984
rect 14004 2975 14056 2984
rect 14004 2941 14013 2975
rect 14013 2941 14047 2975
rect 14047 2941 14056 2975
rect 14004 2932 14056 2941
rect 14924 2932 14976 2984
rect 17500 2932 17552 2984
rect 17592 2975 17644 2984
rect 17592 2941 17601 2975
rect 17601 2941 17635 2975
rect 17635 2941 17644 2975
rect 17592 2932 17644 2941
rect 2872 2796 2924 2848
rect 3792 2796 3844 2848
rect 5908 2796 5960 2848
rect 6184 2796 6236 2848
rect 13636 2864 13688 2916
rect 6920 2796 6972 2848
rect 9036 2796 9088 2848
rect 11060 2796 11112 2848
rect 11336 2839 11388 2848
rect 11336 2805 11345 2839
rect 11345 2805 11379 2839
rect 11379 2805 11388 2839
rect 11336 2796 11388 2805
rect 13728 2796 13780 2848
rect 14740 2796 14792 2848
rect 15016 2839 15068 2848
rect 15016 2805 15025 2839
rect 15025 2805 15059 2839
rect 15059 2805 15068 2839
rect 15016 2796 15068 2805
rect 17500 2839 17552 2848
rect 17500 2805 17509 2839
rect 17509 2805 17543 2839
rect 17543 2805 17552 2839
rect 17500 2796 17552 2805
rect 17776 3043 17828 3052
rect 17776 3009 17785 3043
rect 17785 3009 17819 3043
rect 17819 3009 17828 3043
rect 17776 3000 17828 3009
rect 18788 3043 18840 3052
rect 18788 3009 18797 3043
rect 18797 3009 18831 3043
rect 18831 3009 18840 3043
rect 18788 3000 18840 3009
rect 19708 3000 19760 3052
rect 20352 3000 20404 3052
rect 20720 3043 20772 3052
rect 20720 3009 20729 3043
rect 20729 3009 20763 3043
rect 20763 3009 20772 3043
rect 20720 3000 20772 3009
rect 20904 3068 20956 3120
rect 21824 3068 21876 3120
rect 21456 3000 21508 3052
rect 23388 3000 23440 3052
rect 25136 3068 25188 3120
rect 25780 3136 25832 3188
rect 28540 3136 28592 3188
rect 30104 3136 30156 3188
rect 26148 3068 26200 3120
rect 25504 3043 25556 3052
rect 25504 3009 25513 3043
rect 25513 3009 25547 3043
rect 25547 3009 25556 3043
rect 25504 3000 25556 3009
rect 25780 3043 25832 3052
rect 25780 3009 25789 3043
rect 25789 3009 25823 3043
rect 25823 3009 25832 3043
rect 25780 3000 25832 3009
rect 26332 3000 26384 3052
rect 26792 3043 26844 3052
rect 26792 3009 26801 3043
rect 26801 3009 26835 3043
rect 26835 3009 26844 3043
rect 26792 3000 26844 3009
rect 28632 3068 28684 3120
rect 28540 3000 28592 3052
rect 30564 3136 30616 3188
rect 30748 3136 30800 3188
rect 32864 3136 32916 3188
rect 31208 3068 31260 3120
rect 31484 3068 31536 3120
rect 31944 3068 31996 3120
rect 32220 3068 32272 3120
rect 18328 2932 18380 2984
rect 18236 2907 18288 2916
rect 18236 2873 18245 2907
rect 18245 2873 18279 2907
rect 18279 2873 18288 2907
rect 18236 2864 18288 2873
rect 19248 2864 19300 2916
rect 22008 2975 22060 2984
rect 22008 2941 22017 2975
rect 22017 2941 22051 2975
rect 22051 2941 22060 2975
rect 22008 2932 22060 2941
rect 23572 2975 23624 2984
rect 23572 2941 23581 2975
rect 23581 2941 23615 2975
rect 23615 2941 23624 2975
rect 23572 2932 23624 2941
rect 20352 2864 20404 2916
rect 24216 2975 24268 2984
rect 24216 2941 24225 2975
rect 24225 2941 24259 2975
rect 24259 2941 24268 2975
rect 24216 2932 24268 2941
rect 19432 2839 19484 2848
rect 19432 2805 19441 2839
rect 19441 2805 19475 2839
rect 19475 2805 19484 2839
rect 19432 2796 19484 2805
rect 21456 2839 21508 2848
rect 21456 2805 21465 2839
rect 21465 2805 21499 2839
rect 21499 2805 21508 2839
rect 21456 2796 21508 2805
rect 23204 2796 23256 2848
rect 25964 2839 26016 2848
rect 25964 2805 25973 2839
rect 25973 2805 26007 2839
rect 26007 2805 26016 2839
rect 25964 2796 26016 2805
rect 26608 2839 26660 2848
rect 26608 2805 26617 2839
rect 26617 2805 26651 2839
rect 26651 2805 26660 2839
rect 26608 2796 26660 2805
rect 27252 2796 27304 2848
rect 29644 2975 29696 2984
rect 29644 2941 29653 2975
rect 29653 2941 29687 2975
rect 29687 2941 29696 2975
rect 29644 2932 29696 2941
rect 31576 3043 31628 3052
rect 31576 3009 31585 3043
rect 31585 3009 31619 3043
rect 31619 3009 31628 3043
rect 31576 3000 31628 3009
rect 31668 3000 31720 3052
rect 32864 3000 32916 3052
rect 30748 2864 30800 2916
rect 31944 2932 31996 2984
rect 32128 2975 32180 2984
rect 32128 2941 32137 2975
rect 32137 2941 32171 2975
rect 32171 2941 32180 2975
rect 32128 2932 32180 2941
rect 36268 3136 36320 3188
rect 37372 3136 37424 3188
rect 39396 3179 39448 3188
rect 39396 3145 39405 3179
rect 39405 3145 39439 3179
rect 39439 3145 39448 3179
rect 39396 3136 39448 3145
rect 33048 3068 33100 3120
rect 33416 3043 33468 3052
rect 33416 3009 33425 3043
rect 33425 3009 33459 3043
rect 33459 3009 33468 3043
rect 33416 3000 33468 3009
rect 33692 3043 33744 3052
rect 33692 3009 33701 3043
rect 33701 3009 33735 3043
rect 33735 3009 33744 3043
rect 33692 3000 33744 3009
rect 34244 3068 34296 3120
rect 30380 2796 30432 2848
rect 30472 2796 30524 2848
rect 32864 2864 32916 2916
rect 33048 2796 33100 2848
rect 34336 2864 34388 2916
rect 35716 2864 35768 2916
rect 38844 3043 38896 3052
rect 38844 3009 38853 3043
rect 38853 3009 38887 3043
rect 38887 3009 38896 3043
rect 38844 3000 38896 3009
rect 39488 2932 39540 2984
rect 39764 2864 39816 2916
rect 34704 2796 34756 2848
rect 39028 2839 39080 2848
rect 39028 2805 39037 2839
rect 39037 2805 39071 2839
rect 39071 2805 39080 2839
rect 39028 2796 39080 2805
rect 1950 2694 2002 2746
rect 2014 2694 2066 2746
rect 2078 2694 2130 2746
rect 2142 2694 2194 2746
rect 2206 2694 2258 2746
rect 7950 2694 8002 2746
rect 8014 2694 8066 2746
rect 8078 2694 8130 2746
rect 8142 2694 8194 2746
rect 8206 2694 8258 2746
rect 13950 2694 14002 2746
rect 14014 2694 14066 2746
rect 14078 2694 14130 2746
rect 14142 2694 14194 2746
rect 14206 2694 14258 2746
rect 19950 2694 20002 2746
rect 20014 2694 20066 2746
rect 20078 2694 20130 2746
rect 20142 2694 20194 2746
rect 20206 2694 20258 2746
rect 25950 2694 26002 2746
rect 26014 2694 26066 2746
rect 26078 2694 26130 2746
rect 26142 2694 26194 2746
rect 26206 2694 26258 2746
rect 31950 2694 32002 2746
rect 32014 2694 32066 2746
rect 32078 2694 32130 2746
rect 32142 2694 32194 2746
rect 32206 2694 32258 2746
rect 37950 2694 38002 2746
rect 38014 2694 38066 2746
rect 38078 2694 38130 2746
rect 38142 2694 38194 2746
rect 38206 2694 38258 2746
rect 1584 2592 1636 2644
rect 1768 2592 1820 2644
rect 4712 2592 4764 2644
rect 6000 2635 6052 2644
rect 6000 2601 6009 2635
rect 6009 2601 6043 2635
rect 6043 2601 6052 2635
rect 6000 2592 6052 2601
rect 1124 2524 1176 2576
rect 1308 2456 1360 2508
rect 940 2388 992 2440
rect 2596 2431 2648 2440
rect 2596 2397 2605 2431
rect 2605 2397 2639 2431
rect 2639 2397 2648 2431
rect 2596 2388 2648 2397
rect 3884 2524 3936 2576
rect 11060 2592 11112 2644
rect 13452 2592 13504 2644
rect 14556 2635 14608 2644
rect 4528 2456 4580 2508
rect 4712 2456 4764 2508
rect 4068 2431 4120 2440
rect 4068 2397 4077 2431
rect 4077 2397 4111 2431
rect 4111 2397 4120 2431
rect 4068 2388 4120 2397
rect 4804 2431 4856 2440
rect 4804 2397 4813 2431
rect 4813 2397 4847 2431
rect 4847 2397 4856 2431
rect 4804 2388 4856 2397
rect 5908 2431 5960 2440
rect 5908 2397 5917 2431
rect 5917 2397 5951 2431
rect 5951 2397 5960 2431
rect 5908 2388 5960 2397
rect 6184 2431 6236 2440
rect 6184 2397 6193 2431
rect 6193 2397 6227 2431
rect 6227 2397 6236 2431
rect 6184 2388 6236 2397
rect 7012 2431 7064 2440
rect 7012 2397 7021 2431
rect 7021 2397 7055 2431
rect 7055 2397 7064 2431
rect 7012 2388 7064 2397
rect 7472 2388 7524 2440
rect 10324 2524 10376 2576
rect 10968 2567 11020 2576
rect 10968 2533 10977 2567
rect 10977 2533 11011 2567
rect 11011 2533 11020 2567
rect 10968 2524 11020 2533
rect 11612 2524 11664 2576
rect 14556 2601 14565 2635
rect 14565 2601 14599 2635
rect 14599 2601 14608 2635
rect 14556 2592 14608 2601
rect 14648 2592 14700 2644
rect 15476 2592 15528 2644
rect 15844 2592 15896 2644
rect 18236 2592 18288 2644
rect 21364 2592 21416 2644
rect 22928 2635 22980 2644
rect 22928 2601 22937 2635
rect 22937 2601 22971 2635
rect 22971 2601 22980 2635
rect 22928 2592 22980 2601
rect 26792 2592 26844 2644
rect 388 2320 440 2372
rect 1584 2295 1636 2304
rect 1584 2261 1593 2295
rect 1593 2261 1627 2295
rect 1627 2261 1636 2295
rect 1584 2252 1636 2261
rect 2228 2252 2280 2304
rect 2872 2295 2924 2304
rect 2872 2261 2881 2295
rect 2881 2261 2915 2295
rect 2915 2261 2924 2295
rect 2872 2252 2924 2261
rect 7656 2320 7708 2372
rect 8576 2431 8628 2440
rect 8576 2397 8585 2431
rect 8585 2397 8619 2431
rect 8619 2397 8628 2431
rect 8576 2388 8628 2397
rect 9036 2499 9088 2508
rect 9036 2465 9045 2499
rect 9045 2465 9079 2499
rect 9079 2465 9088 2499
rect 9036 2456 9088 2465
rect 9496 2456 9548 2508
rect 10140 2388 10192 2440
rect 10324 2431 10376 2440
rect 10324 2397 10333 2431
rect 10333 2397 10367 2431
rect 10367 2397 10376 2431
rect 10324 2388 10376 2397
rect 3424 2252 3476 2304
rect 4436 2252 4488 2304
rect 5540 2252 5592 2304
rect 6644 2252 6696 2304
rect 7748 2252 7800 2304
rect 8576 2252 8628 2304
rect 8760 2363 8812 2372
rect 8760 2329 8769 2363
rect 8769 2329 8803 2363
rect 8803 2329 8812 2363
rect 8760 2320 8812 2329
rect 9496 2320 9548 2372
rect 11336 2456 11388 2508
rect 12348 2456 12400 2508
rect 10600 2388 10652 2440
rect 10784 2431 10836 2440
rect 10784 2397 10793 2431
rect 10793 2397 10827 2431
rect 10827 2397 10836 2431
rect 10784 2388 10836 2397
rect 11888 2431 11940 2440
rect 11888 2397 11897 2431
rect 11897 2397 11931 2431
rect 11931 2397 11940 2431
rect 11888 2388 11940 2397
rect 13176 2456 13228 2508
rect 13728 2499 13780 2508
rect 13728 2465 13737 2499
rect 13737 2465 13771 2499
rect 13771 2465 13780 2499
rect 13728 2456 13780 2465
rect 17040 2524 17092 2576
rect 29460 2592 29512 2644
rect 30932 2592 30984 2644
rect 31392 2592 31444 2644
rect 30380 2524 30432 2576
rect 15016 2456 15068 2508
rect 15568 2456 15620 2508
rect 11980 2363 12032 2372
rect 11980 2329 11989 2363
rect 11989 2329 12023 2363
rect 12023 2329 12032 2363
rect 11980 2320 12032 2329
rect 12072 2320 12124 2372
rect 14556 2388 14608 2440
rect 14740 2431 14792 2440
rect 14740 2397 14749 2431
rect 14749 2397 14783 2431
rect 14783 2397 14792 2431
rect 14740 2388 14792 2397
rect 15844 2388 15896 2440
rect 15936 2388 15988 2440
rect 18328 2456 18380 2508
rect 18972 2499 19024 2508
rect 18972 2465 18981 2499
rect 18981 2465 19015 2499
rect 19015 2465 19024 2499
rect 18972 2456 19024 2465
rect 21456 2456 21508 2508
rect 21640 2456 21692 2508
rect 17500 2388 17552 2440
rect 18696 2431 18748 2440
rect 18696 2397 18705 2431
rect 18705 2397 18739 2431
rect 18739 2397 18748 2431
rect 18696 2388 18748 2397
rect 19432 2431 19484 2440
rect 19432 2397 19441 2431
rect 19441 2397 19475 2431
rect 19475 2397 19484 2431
rect 19432 2388 19484 2397
rect 19892 2388 19944 2440
rect 20904 2388 20956 2440
rect 23204 2388 23256 2440
rect 9588 2252 9640 2304
rect 9772 2252 9824 2304
rect 9956 2252 10008 2304
rect 11060 2252 11112 2304
rect 11704 2252 11756 2304
rect 12348 2252 12400 2304
rect 12440 2295 12492 2304
rect 12440 2261 12449 2295
rect 12449 2261 12483 2295
rect 12483 2261 12492 2295
rect 12440 2252 12492 2261
rect 13084 2295 13136 2304
rect 13084 2261 13093 2295
rect 13093 2261 13127 2295
rect 13127 2261 13136 2295
rect 13084 2252 13136 2261
rect 14372 2252 14424 2304
rect 15476 2252 15528 2304
rect 16580 2252 16632 2304
rect 17500 2295 17552 2304
rect 17500 2261 17509 2295
rect 17509 2261 17543 2295
rect 17543 2261 17552 2295
rect 17500 2252 17552 2261
rect 19248 2295 19300 2304
rect 19248 2261 19257 2295
rect 19257 2261 19291 2295
rect 19291 2261 19300 2295
rect 19248 2252 19300 2261
rect 20812 2252 20864 2304
rect 21088 2295 21140 2304
rect 21088 2261 21097 2295
rect 21097 2261 21131 2295
rect 21131 2261 21140 2295
rect 21088 2252 21140 2261
rect 21548 2252 21600 2304
rect 25872 2252 25924 2304
rect 26884 2456 26936 2508
rect 27528 2499 27580 2508
rect 27528 2465 27537 2499
rect 27537 2465 27571 2499
rect 27571 2465 27580 2499
rect 27528 2456 27580 2465
rect 27804 2388 27856 2440
rect 31484 2524 31536 2576
rect 32312 2592 32364 2644
rect 38292 2592 38344 2644
rect 31576 2456 31628 2508
rect 31668 2388 31720 2440
rect 31392 2320 31444 2372
rect 32680 2388 32732 2440
rect 32772 2388 32824 2440
rect 33048 2499 33100 2508
rect 33048 2465 33057 2499
rect 33057 2465 33091 2499
rect 33091 2465 33100 2499
rect 33048 2456 33100 2465
rect 33692 2388 33744 2440
rect 37832 2456 37884 2508
rect 34520 2388 34572 2440
rect 34612 2388 34664 2440
rect 38108 2431 38160 2440
rect 38108 2397 38117 2431
rect 38117 2397 38151 2431
rect 38151 2397 38160 2431
rect 38108 2388 38160 2397
rect 39396 2567 39448 2576
rect 39396 2533 39405 2567
rect 39405 2533 39439 2567
rect 39439 2533 39448 2567
rect 39396 2524 39448 2533
rect 38844 2431 38896 2440
rect 38844 2397 38853 2431
rect 38853 2397 38887 2431
rect 38887 2397 38896 2431
rect 38844 2388 38896 2397
rect 37464 2320 37516 2372
rect 32864 2252 32916 2304
rect 33416 2252 33468 2304
rect 37924 2295 37976 2304
rect 37924 2261 37933 2295
rect 37933 2261 37967 2295
rect 37967 2261 37976 2295
rect 37924 2252 37976 2261
rect 38292 2295 38344 2304
rect 38292 2261 38301 2295
rect 38301 2261 38335 2295
rect 38335 2261 38344 2295
rect 38292 2252 38344 2261
rect 38936 2252 38988 2304
rect 39948 2252 40000 2304
rect 3010 2150 3062 2202
rect 3074 2150 3126 2202
rect 3138 2150 3190 2202
rect 3202 2150 3254 2202
rect 3266 2150 3318 2202
rect 9010 2150 9062 2202
rect 9074 2150 9126 2202
rect 9138 2150 9190 2202
rect 9202 2150 9254 2202
rect 9266 2150 9318 2202
rect 15010 2150 15062 2202
rect 15074 2150 15126 2202
rect 15138 2150 15190 2202
rect 15202 2150 15254 2202
rect 15266 2150 15318 2202
rect 21010 2150 21062 2202
rect 21074 2150 21126 2202
rect 21138 2150 21190 2202
rect 21202 2150 21254 2202
rect 21266 2150 21318 2202
rect 27010 2150 27062 2202
rect 27074 2150 27126 2202
rect 27138 2150 27190 2202
rect 27202 2150 27254 2202
rect 27266 2150 27318 2202
rect 33010 2150 33062 2202
rect 33074 2150 33126 2202
rect 33138 2150 33190 2202
rect 33202 2150 33254 2202
rect 33266 2150 33318 2202
rect 39010 2150 39062 2202
rect 39074 2150 39126 2202
rect 39138 2150 39190 2202
rect 39202 2150 39254 2202
rect 39266 2150 39318 2202
rect 1584 2048 1636 2100
rect 7564 2048 7616 2100
rect 9496 2048 9548 2100
rect 10692 2048 10744 2100
rect 12072 2048 12124 2100
rect 12164 2048 12216 2100
rect 17868 2048 17920 2100
rect 18328 2048 18380 2100
rect 26792 2048 26844 2100
rect 27712 2048 27764 2100
rect 37464 2048 37516 2100
rect 2872 1980 2924 2032
rect 11704 1980 11756 2032
rect 3792 1912 3844 1964
rect 15752 1980 15804 2032
rect 26884 1980 26936 2032
rect 34612 1980 34664 2032
rect 11980 1912 12032 1964
rect 5908 1844 5960 1896
rect 13820 1844 13872 1896
rect 20444 1912 20496 1964
rect 32588 1912 32640 1964
rect 20812 1844 20864 1896
rect 28080 1844 28132 1896
rect 38108 1844 38160 1896
rect 4804 1776 4856 1828
rect 16304 1776 16356 1828
rect 17132 1776 17184 1828
rect 36912 1776 36964 1828
rect 11152 1708 11204 1760
rect 33416 1708 33468 1760
rect 10140 1640 10192 1692
rect 11244 1640 11296 1692
rect 11980 1640 12032 1692
rect 12532 1640 12584 1692
rect 31576 1640 31628 1692
rect 1768 1572 1820 1624
rect 17960 1572 18012 1624
rect 25872 1572 25924 1624
rect 30012 1572 30064 1624
rect 7656 1504 7708 1556
rect 12808 1504 12860 1556
rect 11152 1436 11204 1488
rect 32496 1436 32548 1488
rect 6736 1300 6788 1352
rect 35072 1300 35124 1352
rect 10968 1232 11020 1284
rect 39580 1232 39632 1284
rect 13084 1164 13136 1216
rect 38844 1164 38896 1216
rect 7564 1096 7616 1148
rect 17316 1096 17368 1148
rect 3516 1028 3568 1080
rect 28172 1028 28224 1080
rect 10232 960 10284 1012
rect 33876 960 33928 1012
rect 8760 892 8812 944
rect 29828 892 29880 944
rect 7380 824 7432 876
rect 23480 824 23532 876
rect 4528 756 4580 808
rect 18420 756 18472 808
rect 7472 688 7524 740
rect 27528 688 27580 740
rect 1492 620 1544 672
rect 18052 620 18104 672
rect 7288 552 7340 604
rect 23940 552 23992 604
rect 4712 484 4764 536
rect 29552 484 29604 536
rect 2504 416 2556 468
rect 16948 416 17000 468
rect 23204 144 23256 196
rect 24308 144 24360 196
rect 38568 144 38620 196
rect 37740 76 37792 128
rect 22192 8 22244 60
rect 39488 8 39540 60
<< metal2 >>
rect 2884 11206 3188 11234
rect 1492 10464 1544 10470
rect 1492 10406 1544 10412
rect 1306 9616 1362 9625
rect 1306 9551 1362 9560
rect 110 9344 166 9353
rect 110 9279 166 9288
rect 124 5030 152 9279
rect 386 9072 442 9081
rect 386 9007 442 9016
rect 202 8800 258 8809
rect 202 8735 258 8744
rect 112 5024 164 5030
rect 112 4966 164 4972
rect 216 4486 244 8735
rect 294 6352 350 6361
rect 294 6287 350 6296
rect 204 4480 256 4486
rect 204 4422 256 4428
rect 308 4146 336 6287
rect 400 5642 428 9007
rect 846 8528 902 8537
rect 846 8463 902 8472
rect 756 7880 808 7886
rect 756 7822 808 7828
rect 768 7721 796 7822
rect 754 7712 810 7721
rect 754 7647 810 7656
rect 754 7440 810 7449
rect 754 7375 756 7384
rect 808 7375 810 7384
rect 756 7346 808 7352
rect 754 7168 810 7177
rect 754 7103 810 7112
rect 478 5808 534 5817
rect 478 5743 534 5752
rect 388 5636 440 5642
rect 388 5578 440 5584
rect 386 4176 442 4185
rect 296 4140 348 4146
rect 386 4111 442 4120
rect 296 4082 348 4088
rect 400 3602 428 4111
rect 388 3596 440 3602
rect 388 3538 440 3544
rect 492 2990 520 5743
rect 570 5264 626 5273
rect 570 5199 626 5208
rect 584 3942 612 5199
rect 768 4690 796 7103
rect 860 5234 888 8463
rect 1124 8424 1176 8430
rect 1124 8366 1176 8372
rect 1136 8265 1164 8366
rect 1122 8256 1178 8265
rect 1122 8191 1178 8200
rect 1214 7984 1270 7993
rect 1214 7919 1216 7928
rect 1268 7919 1270 7928
rect 1216 7890 1268 7896
rect 1030 6896 1086 6905
rect 1030 6831 1086 6840
rect 938 6624 994 6633
rect 938 6559 994 6568
rect 848 5228 900 5234
rect 848 5170 900 5176
rect 952 5166 980 6559
rect 1044 5710 1072 6831
rect 1320 6390 1348 9551
rect 1400 8968 1452 8974
rect 1400 8910 1452 8916
rect 1412 8498 1440 8910
rect 1400 8492 1452 8498
rect 1400 8434 1452 8440
rect 1400 6860 1452 6866
rect 1400 6802 1452 6808
rect 1308 6384 1360 6390
rect 1308 6326 1360 6332
rect 1214 6080 1270 6089
rect 1214 6015 1270 6024
rect 1032 5704 1084 5710
rect 1032 5646 1084 5652
rect 1030 5536 1086 5545
rect 1030 5471 1086 5480
rect 940 5160 992 5166
rect 940 5102 992 5108
rect 756 4684 808 4690
rect 756 4626 808 4632
rect 756 4072 808 4078
rect 756 4014 808 4020
rect 572 3936 624 3942
rect 768 3913 796 4014
rect 572 3878 624 3884
rect 754 3904 810 3913
rect 754 3839 810 3848
rect 754 3632 810 3641
rect 754 3567 810 3576
rect 768 3534 796 3567
rect 756 3528 808 3534
rect 756 3470 808 3476
rect 1044 3126 1072 5471
rect 1228 5302 1256 6015
rect 1216 5296 1268 5302
rect 1216 5238 1268 5244
rect 1306 4992 1362 5001
rect 1306 4927 1362 4936
rect 1124 4752 1176 4758
rect 1122 4720 1124 4729
rect 1176 4720 1178 4729
rect 1122 4655 1178 4664
rect 1122 4448 1178 4457
rect 1122 4383 1178 4392
rect 1136 3670 1164 4383
rect 1320 3738 1348 4927
rect 1308 3732 1360 3738
rect 1308 3674 1360 3680
rect 1124 3664 1176 3670
rect 1124 3606 1176 3612
rect 1032 3120 1084 3126
rect 1032 3062 1084 3068
rect 572 3052 624 3058
rect 572 2994 624 3000
rect 480 2984 532 2990
rect 480 2926 532 2932
rect 584 2825 612 2994
rect 570 2816 626 2825
rect 570 2751 626 2760
rect 1412 2774 1440 6802
rect 1504 6458 1532 10406
rect 2044 10260 2096 10266
rect 2044 10202 2096 10208
rect 1768 9784 1820 9790
rect 1768 9726 1820 9732
rect 1676 9512 1728 9518
rect 1676 9454 1728 9460
rect 1584 8900 1636 8906
rect 1584 8842 1636 8848
rect 1596 8634 1624 8842
rect 1584 8628 1636 8634
rect 1584 8570 1636 8576
rect 1688 8498 1716 9454
rect 1676 8492 1728 8498
rect 1676 8434 1728 8440
rect 1584 7336 1636 7342
rect 1584 7278 1636 7284
rect 1492 6452 1544 6458
rect 1492 6394 1544 6400
rect 1492 5364 1544 5370
rect 1492 5306 1544 5312
rect 1504 4826 1532 5306
rect 1492 4820 1544 4826
rect 1492 4762 1544 4768
rect 1412 2746 1532 2774
rect 1124 2576 1176 2582
rect 1124 2518 1176 2524
rect 940 2440 992 2446
rect 940 2382 992 2388
rect 388 2372 440 2378
rect 388 2314 440 2320
rect 400 1737 428 2314
rect 386 1728 442 1737
rect 386 1663 442 1672
rect 952 1465 980 2382
rect 938 1456 994 1465
rect 938 1391 994 1400
rect 1136 56 1164 2518
rect 1308 2508 1360 2514
rect 1308 2450 1360 2456
rect 1320 2281 1348 2450
rect 1306 2272 1362 2281
rect 1306 2207 1362 2216
rect 1504 678 1532 2746
rect 1596 2650 1624 7278
rect 1676 6724 1728 6730
rect 1676 6666 1728 6672
rect 1688 3380 1716 6666
rect 1780 6662 1808 9726
rect 1860 9172 1912 9178
rect 1860 9114 1912 9120
rect 1872 8498 1900 9114
rect 1860 8492 1912 8498
rect 1860 8434 1912 8440
rect 2056 8378 2084 10202
rect 2318 9888 2374 9897
rect 2318 9823 2374 9832
rect 2136 9240 2188 9246
rect 2136 9182 2188 9188
rect 2148 8498 2176 9182
rect 2136 8492 2188 8498
rect 2136 8434 2188 8440
rect 1872 8350 2084 8378
rect 1768 6656 1820 6662
rect 1768 6598 1820 6604
rect 1872 6440 1900 8350
rect 1950 8188 2258 8197
rect 1950 8186 1956 8188
rect 2012 8186 2036 8188
rect 2092 8186 2116 8188
rect 2172 8186 2196 8188
rect 2252 8186 2258 8188
rect 2012 8134 2014 8186
rect 2194 8134 2196 8186
rect 1950 8132 1956 8134
rect 2012 8132 2036 8134
rect 2092 8132 2116 8134
rect 2172 8132 2196 8134
rect 2252 8132 2258 8134
rect 1950 8123 2258 8132
rect 1950 7100 2258 7109
rect 1950 7098 1956 7100
rect 2012 7098 2036 7100
rect 2092 7098 2116 7100
rect 2172 7098 2196 7100
rect 2252 7098 2258 7100
rect 2012 7046 2014 7098
rect 2194 7046 2196 7098
rect 1950 7044 1956 7046
rect 2012 7044 2036 7046
rect 2092 7044 2116 7046
rect 2172 7044 2196 7046
rect 2252 7044 2258 7046
rect 1950 7035 2258 7044
rect 2228 6656 2280 6662
rect 2228 6598 2280 6604
rect 1780 6412 1900 6440
rect 1780 5370 1808 6412
rect 2240 6361 2268 6598
rect 2226 6352 2282 6361
rect 1860 6316 1912 6322
rect 2226 6287 2282 6296
rect 1860 6258 1912 6264
rect 1768 5364 1820 5370
rect 1768 5306 1820 5312
rect 1766 5128 1822 5137
rect 1766 5063 1768 5072
rect 1820 5063 1822 5072
rect 1768 5034 1820 5040
rect 1768 3392 1820 3398
rect 1688 3352 1768 3380
rect 1768 3334 1820 3340
rect 1872 2774 1900 6258
rect 2136 6248 2188 6254
rect 2134 6216 2136 6225
rect 2188 6216 2190 6225
rect 2134 6151 2190 6160
rect 1950 6012 2258 6021
rect 1950 6010 1956 6012
rect 2012 6010 2036 6012
rect 2092 6010 2116 6012
rect 2172 6010 2196 6012
rect 2252 6010 2258 6012
rect 2012 5958 2014 6010
rect 2194 5958 2196 6010
rect 1950 5956 1956 5958
rect 2012 5956 2036 5958
rect 2092 5956 2116 5958
rect 2172 5956 2196 5958
rect 2252 5956 2258 5958
rect 1950 5947 2258 5956
rect 2332 5710 2360 9823
rect 2502 9208 2558 9217
rect 2502 9143 2558 9152
rect 2516 8498 2544 9143
rect 2504 8492 2556 8498
rect 2504 8434 2556 8440
rect 2596 8288 2648 8294
rect 2596 8230 2648 8236
rect 2688 8288 2740 8294
rect 2688 8230 2740 8236
rect 2608 8129 2636 8230
rect 2594 8120 2650 8129
rect 2594 8055 2650 8064
rect 2412 7880 2464 7886
rect 2596 7880 2648 7886
rect 2412 7822 2464 7828
rect 2594 7848 2596 7857
rect 2648 7848 2650 7857
rect 2424 6474 2452 7822
rect 2504 7812 2556 7818
rect 2594 7783 2650 7792
rect 2504 7754 2556 7760
rect 2516 7546 2544 7754
rect 2700 7732 2728 8230
rect 2608 7704 2728 7732
rect 2780 7744 2832 7750
rect 2504 7540 2556 7546
rect 2504 7482 2556 7488
rect 2424 6446 2544 6474
rect 2412 6384 2464 6390
rect 2412 6326 2464 6332
rect 2320 5704 2372 5710
rect 2320 5646 2372 5652
rect 1950 4924 2258 4933
rect 1950 4922 1956 4924
rect 2012 4922 2036 4924
rect 2092 4922 2116 4924
rect 2172 4922 2196 4924
rect 2252 4922 2258 4924
rect 2012 4870 2014 4922
rect 2194 4870 2196 4922
rect 1950 4868 1956 4870
rect 2012 4868 2036 4870
rect 2092 4868 2116 4870
rect 2172 4868 2196 4870
rect 2252 4868 2258 4870
rect 1950 4859 2258 4868
rect 2424 4826 2452 6326
rect 2516 6089 2544 6446
rect 2502 6080 2558 6089
rect 2502 6015 2558 6024
rect 2502 5944 2558 5953
rect 2502 5879 2504 5888
rect 2556 5879 2558 5888
rect 2504 5850 2556 5856
rect 2504 5704 2556 5710
rect 2502 5672 2504 5681
rect 2556 5672 2558 5681
rect 2502 5607 2558 5616
rect 2504 5568 2556 5574
rect 2504 5510 2556 5516
rect 2412 4820 2464 4826
rect 2412 4762 2464 4768
rect 2042 4584 2098 4593
rect 2042 4519 2044 4528
rect 2096 4519 2098 4528
rect 2044 4490 2096 4496
rect 2516 4026 2544 5510
rect 2608 4622 2636 7704
rect 2780 7686 2832 7692
rect 2688 7540 2740 7546
rect 2688 7482 2740 7488
rect 2700 7426 2728 7482
rect 2792 7426 2820 7686
rect 2700 7398 2820 7426
rect 2780 7336 2832 7342
rect 2780 7278 2832 7284
rect 2686 6352 2742 6361
rect 2686 6287 2742 6296
rect 2700 5846 2728 6287
rect 2688 5840 2740 5846
rect 2688 5782 2740 5788
rect 2792 5370 2820 7278
rect 2884 6458 2912 11206
rect 3160 11098 3188 11206
rect 3238 11194 3294 11250
rect 3514 11194 3570 11250
rect 3790 11194 3846 11250
rect 4066 11194 4122 11250
rect 4342 11194 4398 11250
rect 4618 11194 4674 11250
rect 4894 11194 4950 11250
rect 5170 11194 5226 11250
rect 5446 11194 5502 11250
rect 5722 11194 5778 11250
rect 5998 11194 6054 11250
rect 6274 11194 6330 11250
rect 6550 11194 6606 11250
rect 6644 11212 6696 11218
rect 3252 11098 3280 11194
rect 3160 11070 3280 11098
rect 3528 10470 3556 11194
rect 3516 10464 3568 10470
rect 3516 10406 3568 10412
rect 3700 9988 3752 9994
rect 3700 9930 3752 9936
rect 3424 9716 3476 9722
rect 3424 9658 3476 9664
rect 3010 8732 3318 8741
rect 3010 8730 3016 8732
rect 3072 8730 3096 8732
rect 3152 8730 3176 8732
rect 3232 8730 3256 8732
rect 3312 8730 3318 8732
rect 3072 8678 3074 8730
rect 3254 8678 3256 8730
rect 3010 8676 3016 8678
rect 3072 8676 3096 8678
rect 3152 8676 3176 8678
rect 3232 8676 3256 8678
rect 3312 8676 3318 8678
rect 3010 8667 3318 8676
rect 3010 7644 3318 7653
rect 3010 7642 3016 7644
rect 3072 7642 3096 7644
rect 3152 7642 3176 7644
rect 3232 7642 3256 7644
rect 3312 7642 3318 7644
rect 3072 7590 3074 7642
rect 3254 7590 3256 7642
rect 3010 7588 3016 7590
rect 3072 7588 3096 7590
rect 3152 7588 3176 7590
rect 3232 7588 3256 7590
rect 3312 7588 3318 7590
rect 3010 7579 3318 7588
rect 3436 7546 3464 9658
rect 3514 9072 3570 9081
rect 3514 9007 3570 9016
rect 3608 9036 3660 9042
rect 3528 8634 3556 9007
rect 3608 8978 3660 8984
rect 3516 8628 3568 8634
rect 3516 8570 3568 8576
rect 3424 7540 3476 7546
rect 3424 7482 3476 7488
rect 3148 7404 3200 7410
rect 3148 7346 3200 7352
rect 3160 6866 3188 7346
rect 3332 7336 3384 7342
rect 3332 7278 3384 7284
rect 3240 7268 3292 7274
rect 3240 7210 3292 7216
rect 3252 7041 3280 7210
rect 3238 7032 3294 7041
rect 3238 6967 3294 6976
rect 3240 6928 3292 6934
rect 3238 6896 3240 6905
rect 3292 6896 3294 6905
rect 3148 6860 3200 6866
rect 3238 6831 3294 6840
rect 3148 6802 3200 6808
rect 3240 6792 3292 6798
rect 3238 6760 3240 6769
rect 3292 6760 3294 6769
rect 3344 6746 3372 7278
rect 3620 7002 3648 8978
rect 3608 6996 3660 7002
rect 3608 6938 3660 6944
rect 3516 6860 3568 6866
rect 3568 6820 3648 6848
rect 3516 6802 3568 6808
rect 3344 6718 3556 6746
rect 3238 6695 3294 6704
rect 3332 6656 3384 6662
rect 3384 6604 3464 6610
rect 3332 6598 3464 6604
rect 3344 6582 3464 6598
rect 3010 6556 3318 6565
rect 3010 6554 3016 6556
rect 3072 6554 3096 6556
rect 3152 6554 3176 6556
rect 3232 6554 3256 6556
rect 3312 6554 3318 6556
rect 3072 6502 3074 6554
rect 3254 6502 3256 6554
rect 3010 6500 3016 6502
rect 3072 6500 3096 6502
rect 3152 6500 3176 6502
rect 3232 6500 3256 6502
rect 3312 6500 3318 6502
rect 3010 6491 3318 6500
rect 3436 6458 3464 6582
rect 2872 6452 2924 6458
rect 2872 6394 2924 6400
rect 3424 6452 3476 6458
rect 3424 6394 3476 6400
rect 3528 6338 3556 6718
rect 3436 6310 3556 6338
rect 3332 6248 3384 6254
rect 3332 6190 3384 6196
rect 3148 6180 3200 6186
rect 3148 6122 3200 6128
rect 2872 6112 2924 6118
rect 2872 6054 2924 6060
rect 2780 5364 2832 5370
rect 2780 5306 2832 5312
rect 2780 5092 2832 5098
rect 2780 5034 2832 5040
rect 2596 4616 2648 4622
rect 2596 4558 2648 4564
rect 2688 4480 2740 4486
rect 2688 4422 2740 4428
rect 2700 4214 2728 4422
rect 2688 4208 2740 4214
rect 2792 4185 2820 5034
rect 2884 4622 2912 6054
rect 3160 5817 3188 6122
rect 3344 5914 3372 6190
rect 3332 5908 3384 5914
rect 3332 5850 3384 5856
rect 3146 5808 3202 5817
rect 3146 5743 3202 5752
rect 3436 5522 3464 6310
rect 3620 6118 3648 6820
rect 3712 6118 3740 9930
rect 3804 6662 3832 11194
rect 3884 8832 3936 8838
rect 3884 8774 3936 8780
rect 3896 8498 3924 8774
rect 3976 8560 4028 8566
rect 3976 8502 4028 8508
rect 3884 8492 3936 8498
rect 3884 8434 3936 8440
rect 3884 7812 3936 7818
rect 3884 7754 3936 7760
rect 3896 7002 3924 7754
rect 3988 7721 4016 8502
rect 4080 8378 4108 11194
rect 4356 9790 4384 11194
rect 4526 10296 4582 10305
rect 4526 10231 4582 10240
rect 4344 9784 4396 9790
rect 4344 9726 4396 9732
rect 4434 9616 4490 9625
rect 4434 9551 4490 9560
rect 4252 9376 4304 9382
rect 4252 9318 4304 9324
rect 4080 8350 4200 8378
rect 4068 7880 4120 7886
rect 4068 7822 4120 7828
rect 3974 7712 4030 7721
rect 3974 7647 4030 7656
rect 4080 7410 4108 7822
rect 4068 7404 4120 7410
rect 4068 7346 4120 7352
rect 3976 7336 4028 7342
rect 3976 7278 4028 7284
rect 3884 6996 3936 7002
rect 3884 6938 3936 6944
rect 3792 6656 3844 6662
rect 3792 6598 3844 6604
rect 3884 6656 3936 6662
rect 3884 6598 3936 6604
rect 3608 6112 3660 6118
rect 3608 6054 3660 6060
rect 3700 6112 3752 6118
rect 3700 6054 3752 6060
rect 3528 5642 3648 5658
rect 3516 5636 3648 5642
rect 3568 5630 3648 5636
rect 3516 5578 3568 5584
rect 3514 5536 3570 5545
rect 3436 5494 3514 5522
rect 3010 5468 3318 5477
rect 3514 5471 3570 5480
rect 3010 5466 3016 5468
rect 3072 5466 3096 5468
rect 3152 5466 3176 5468
rect 3232 5466 3256 5468
rect 3312 5466 3318 5468
rect 3072 5414 3074 5466
rect 3254 5414 3256 5466
rect 3010 5412 3016 5414
rect 3072 5412 3096 5414
rect 3152 5412 3176 5414
rect 3232 5412 3256 5414
rect 3312 5412 3318 5414
rect 3010 5403 3318 5412
rect 3528 5234 3556 5471
rect 3620 5234 3648 5630
rect 3896 5302 3924 6598
rect 3988 6390 4016 7278
rect 4068 6928 4120 6934
rect 4068 6870 4120 6876
rect 3976 6384 4028 6390
rect 3976 6326 4028 6332
rect 3976 6180 4028 6186
rect 3976 6122 4028 6128
rect 3988 5953 4016 6122
rect 3974 5944 4030 5953
rect 3974 5879 4030 5888
rect 3976 5704 4028 5710
rect 3976 5646 4028 5652
rect 3884 5296 3936 5302
rect 3884 5238 3936 5244
rect 3516 5228 3568 5234
rect 3516 5170 3568 5176
rect 3608 5228 3660 5234
rect 3608 5170 3660 5176
rect 3424 5024 3476 5030
rect 3424 4966 3476 4972
rect 2872 4616 2924 4622
rect 2872 4558 2924 4564
rect 3010 4380 3318 4389
rect 3010 4378 3016 4380
rect 3072 4378 3096 4380
rect 3152 4378 3176 4380
rect 3232 4378 3256 4380
rect 3312 4378 3318 4380
rect 3072 4326 3074 4378
rect 3254 4326 3256 4378
rect 3010 4324 3016 4326
rect 3072 4324 3096 4326
rect 3152 4324 3176 4326
rect 3232 4324 3256 4326
rect 3312 4324 3318 4326
rect 3010 4315 3318 4324
rect 2872 4208 2924 4214
rect 2688 4150 2740 4156
rect 2778 4176 2834 4185
rect 2872 4150 2924 4156
rect 2778 4111 2834 4120
rect 2424 3998 2544 4026
rect 2688 4072 2740 4078
rect 2688 4014 2740 4020
rect 2778 4040 2834 4049
rect 2320 3936 2372 3942
rect 2320 3878 2372 3884
rect 1950 3836 2258 3845
rect 1950 3834 1956 3836
rect 2012 3834 2036 3836
rect 2092 3834 2116 3836
rect 2172 3834 2196 3836
rect 2252 3834 2258 3836
rect 2012 3782 2014 3834
rect 2194 3782 2196 3834
rect 1950 3780 1956 3782
rect 2012 3780 2036 3782
rect 2092 3780 2116 3782
rect 2172 3780 2196 3782
rect 2252 3780 2258 3782
rect 1950 3771 2258 3780
rect 1952 3664 2004 3670
rect 1952 3606 2004 3612
rect 1964 3194 1992 3606
rect 2332 3534 2360 3878
rect 2320 3528 2372 3534
rect 2320 3470 2372 3476
rect 1952 3188 2004 3194
rect 1952 3130 2004 3136
rect 2320 3052 2372 3058
rect 2320 2994 2372 3000
rect 1688 2746 1900 2774
rect 1950 2748 2258 2757
rect 1950 2746 1956 2748
rect 2012 2746 2036 2748
rect 2092 2746 2116 2748
rect 2172 2746 2196 2748
rect 2252 2746 2258 2748
rect 1584 2644 1636 2650
rect 1584 2586 1636 2592
rect 1688 2417 1716 2746
rect 2012 2694 2014 2746
rect 2194 2694 2196 2746
rect 1950 2692 1956 2694
rect 2012 2692 2036 2694
rect 2092 2692 2116 2694
rect 2172 2692 2196 2694
rect 2252 2692 2258 2694
rect 1950 2683 2258 2692
rect 1768 2644 1820 2650
rect 1768 2586 1820 2592
rect 1674 2408 1730 2417
rect 1674 2343 1730 2352
rect 1584 2304 1636 2310
rect 1584 2246 1636 2252
rect 1596 2106 1624 2246
rect 1584 2100 1636 2106
rect 1584 2042 1636 2048
rect 1780 1630 1808 2586
rect 2228 2304 2280 2310
rect 2228 2246 2280 2252
rect 1768 1624 1820 1630
rect 1768 1566 1820 1572
rect 1492 672 1544 678
rect 1492 614 1544 620
rect 2240 56 2268 2246
rect 2332 2009 2360 2994
rect 2424 2922 2452 3998
rect 2504 3936 2556 3942
rect 2504 3878 2556 3884
rect 2412 2916 2464 2922
rect 2412 2858 2464 2864
rect 2318 2000 2374 2009
rect 2318 1935 2374 1944
rect 2516 474 2544 3878
rect 2700 3670 2728 4014
rect 2778 3975 2834 3984
rect 2688 3664 2740 3670
rect 2688 3606 2740 3612
rect 2688 3528 2740 3534
rect 2688 3470 2740 3476
rect 2700 3369 2728 3470
rect 2792 3466 2820 3975
rect 2780 3460 2832 3466
rect 2780 3402 2832 3408
rect 2884 3398 2912 4150
rect 3054 3496 3110 3505
rect 3054 3431 3110 3440
rect 3068 3398 3096 3431
rect 2872 3392 2924 3398
rect 2686 3360 2742 3369
rect 2872 3334 2924 3340
rect 3056 3392 3108 3398
rect 3056 3334 3108 3340
rect 2686 3295 2742 3304
rect 2686 3088 2742 3097
rect 2596 3052 2648 3058
rect 2686 3023 2688 3032
rect 2596 2994 2648 3000
rect 2740 3023 2742 3032
rect 2688 2994 2740 3000
rect 2608 2553 2636 2994
rect 2884 2854 2912 3334
rect 3010 3292 3318 3301
rect 3010 3290 3016 3292
rect 3072 3290 3096 3292
rect 3152 3290 3176 3292
rect 3232 3290 3256 3292
rect 3312 3290 3318 3292
rect 3072 3238 3074 3290
rect 3254 3238 3256 3290
rect 3010 3236 3016 3238
rect 3072 3236 3096 3238
rect 3152 3236 3176 3238
rect 3232 3236 3256 3238
rect 3312 3236 3318 3238
rect 3010 3227 3318 3236
rect 2872 2848 2924 2854
rect 2872 2790 2924 2796
rect 3436 2774 3464 4966
rect 3620 2990 3648 5170
rect 3884 4684 3936 4690
rect 3884 4626 3936 4632
rect 3896 4282 3924 4626
rect 3884 4276 3936 4282
rect 3884 4218 3936 4224
rect 3988 4162 4016 5646
rect 4080 4486 4108 6870
rect 4172 5914 4200 8350
rect 4264 6934 4292 9318
rect 4448 8634 4476 9551
rect 4436 8628 4488 8634
rect 4436 8570 4488 8576
rect 4344 7200 4396 7206
rect 4344 7142 4396 7148
rect 4434 7168 4490 7177
rect 4356 6934 4384 7142
rect 4434 7103 4490 7112
rect 4252 6928 4304 6934
rect 4252 6870 4304 6876
rect 4344 6928 4396 6934
rect 4344 6870 4396 6876
rect 4252 6792 4304 6798
rect 4250 6760 4252 6769
rect 4304 6760 4306 6769
rect 4250 6695 4306 6704
rect 4448 6474 4476 7103
rect 4356 6446 4476 6474
rect 4356 6390 4384 6446
rect 4344 6384 4396 6390
rect 4344 6326 4396 6332
rect 4436 6316 4488 6322
rect 4436 6258 4488 6264
rect 4160 5908 4212 5914
rect 4160 5850 4212 5856
rect 4342 5808 4398 5817
rect 4342 5743 4398 5752
rect 4068 4480 4120 4486
rect 4068 4422 4120 4428
rect 4356 4282 4384 5743
rect 4344 4276 4396 4282
rect 4344 4218 4396 4224
rect 3896 4134 4016 4162
rect 3792 4072 3844 4078
rect 3792 4014 3844 4020
rect 3804 3670 3832 4014
rect 3792 3664 3844 3670
rect 3792 3606 3844 3612
rect 3700 3392 3752 3398
rect 3700 3334 3752 3340
rect 3712 2990 3740 3334
rect 3608 2984 3660 2990
rect 3608 2926 3660 2932
rect 3700 2984 3752 2990
rect 3700 2926 3752 2932
rect 3792 2848 3844 2854
rect 3792 2790 3844 2796
rect 3436 2746 3556 2774
rect 2594 2544 2650 2553
rect 2594 2479 2650 2488
rect 2596 2440 2648 2446
rect 2596 2382 2648 2388
rect 2608 649 2636 2382
rect 2872 2304 2924 2310
rect 2872 2246 2924 2252
rect 3424 2304 3476 2310
rect 3424 2246 3476 2252
rect 2884 2038 2912 2246
rect 3010 2204 3318 2213
rect 3010 2202 3016 2204
rect 3072 2202 3096 2204
rect 3152 2202 3176 2204
rect 3232 2202 3256 2204
rect 3312 2202 3318 2204
rect 3072 2150 3074 2202
rect 3254 2150 3256 2202
rect 3010 2148 3016 2150
rect 3072 2148 3096 2150
rect 3152 2148 3176 2150
rect 3232 2148 3256 2150
rect 3312 2148 3318 2150
rect 3010 2139 3318 2148
rect 2872 2032 2924 2038
rect 2872 1974 2924 1980
rect 3436 1170 3464 2246
rect 3344 1142 3464 1170
rect 2594 640 2650 649
rect 2594 575 2650 584
rect 2504 468 2556 474
rect 2504 410 2556 416
rect 3344 56 3372 1142
rect 3528 1086 3556 2746
rect 3804 1970 3832 2790
rect 3896 2582 3924 4134
rect 4344 3664 4396 3670
rect 4342 3632 4344 3641
rect 4396 3632 4398 3641
rect 4342 3567 4398 3576
rect 3976 3392 4028 3398
rect 3976 3334 4028 3340
rect 3884 2576 3936 2582
rect 3884 2518 3936 2524
rect 3792 1964 3844 1970
rect 3792 1906 3844 1912
rect 3516 1080 3568 1086
rect 3516 1022 3568 1028
rect 3988 785 4016 3334
rect 4066 2952 4122 2961
rect 4066 2887 4068 2896
rect 4120 2887 4122 2896
rect 4068 2858 4120 2864
rect 4068 2440 4120 2446
rect 4068 2382 4120 2388
rect 4448 2394 4476 6258
rect 4540 6186 4568 10231
rect 4632 9722 4660 11194
rect 4710 10704 4766 10713
rect 4710 10639 4766 10648
rect 4620 9716 4672 9722
rect 4620 9658 4672 9664
rect 4724 9602 4752 10639
rect 4632 9574 4752 9602
rect 4632 6322 4660 9574
rect 4804 8492 4856 8498
rect 4804 8434 4856 8440
rect 4712 8424 4764 8430
rect 4712 8366 4764 8372
rect 4724 8090 4752 8366
rect 4712 8084 4764 8090
rect 4712 8026 4764 8032
rect 4712 6656 4764 6662
rect 4712 6598 4764 6604
rect 4620 6316 4672 6322
rect 4620 6258 4672 6264
rect 4528 6180 4580 6186
rect 4528 6122 4580 6128
rect 4620 6180 4672 6186
rect 4620 6122 4672 6128
rect 4632 5914 4660 6122
rect 4724 6118 4752 6598
rect 4712 6112 4764 6118
rect 4712 6054 4764 6060
rect 4620 5908 4672 5914
rect 4620 5850 4672 5856
rect 4528 5704 4580 5710
rect 4528 5646 4580 5652
rect 4540 2514 4568 5646
rect 4632 5642 4660 5850
rect 4712 5772 4764 5778
rect 4712 5714 4764 5720
rect 4620 5636 4672 5642
rect 4620 5578 4672 5584
rect 4620 5024 4672 5030
rect 4620 4966 4672 4972
rect 4528 2508 4580 2514
rect 4528 2450 4580 2456
rect 4080 1873 4108 2382
rect 4448 2366 4568 2394
rect 4436 2304 4488 2310
rect 4436 2246 4488 2252
rect 4066 1864 4122 1873
rect 4066 1799 4122 1808
rect 3974 776 4030 785
rect 3974 711 4030 720
rect 4448 56 4476 2246
rect 4540 814 4568 2366
rect 4632 1329 4660 4966
rect 4724 3618 4752 5714
rect 4816 4826 4844 8434
rect 4908 8022 4936 11194
rect 4986 10568 5042 10577
rect 4986 10503 5042 10512
rect 4896 8016 4948 8022
rect 4896 7958 4948 7964
rect 4896 7744 4948 7750
rect 4896 7686 4948 7692
rect 4908 7478 4936 7686
rect 5000 7546 5028 10503
rect 5184 8106 5212 11194
rect 5262 10432 5318 10441
rect 5262 10367 5318 10376
rect 5092 8078 5212 8106
rect 4988 7540 5040 7546
rect 4988 7482 5040 7488
rect 4896 7472 4948 7478
rect 4896 7414 4948 7420
rect 4988 6792 5040 6798
rect 4988 6734 5040 6740
rect 4894 6624 4950 6633
rect 4894 6559 4950 6568
rect 4804 4820 4856 4826
rect 4804 4762 4856 4768
rect 4724 3590 4844 3618
rect 4712 3528 4764 3534
rect 4712 3470 4764 3476
rect 4724 3126 4752 3470
rect 4712 3120 4764 3126
rect 4712 3062 4764 3068
rect 4816 2774 4844 3590
rect 4908 3097 4936 6559
rect 5000 4010 5028 6734
rect 5092 5846 5120 8078
rect 5172 7948 5224 7954
rect 5172 7890 5224 7896
rect 5184 7546 5212 7890
rect 5172 7540 5224 7546
rect 5172 7482 5224 7488
rect 5170 7440 5226 7449
rect 5170 7375 5226 7384
rect 5184 6866 5212 7375
rect 5172 6860 5224 6866
rect 5172 6802 5224 6808
rect 5276 6746 5304 10367
rect 5460 9194 5488 11194
rect 5632 9308 5684 9314
rect 5632 9250 5684 9256
rect 5184 6718 5304 6746
rect 5368 9166 5488 9194
rect 5540 9240 5592 9246
rect 5540 9182 5592 9188
rect 5184 6662 5212 6718
rect 5172 6656 5224 6662
rect 5172 6598 5224 6604
rect 5264 6656 5316 6662
rect 5264 6598 5316 6604
rect 5170 6488 5226 6497
rect 5170 6423 5226 6432
rect 5080 5840 5132 5846
rect 5080 5782 5132 5788
rect 5184 5658 5212 6423
rect 5092 5630 5212 5658
rect 4988 4004 5040 4010
rect 4988 3946 5040 3952
rect 5092 3924 5120 5630
rect 5172 5568 5224 5574
rect 5172 5510 5224 5516
rect 5184 4146 5212 5510
rect 5276 4146 5304 6598
rect 5368 6458 5396 9166
rect 5448 9104 5500 9110
rect 5448 9046 5500 9052
rect 5460 8634 5488 9046
rect 5448 8628 5500 8634
rect 5448 8570 5500 8576
rect 5448 6996 5500 7002
rect 5448 6938 5500 6944
rect 5460 6798 5488 6938
rect 5448 6792 5500 6798
rect 5448 6734 5500 6740
rect 5460 6633 5488 6734
rect 5446 6624 5502 6633
rect 5446 6559 5502 6568
rect 5446 6488 5502 6497
rect 5356 6452 5408 6458
rect 5552 6474 5580 9182
rect 5644 7886 5672 9250
rect 5632 7880 5684 7886
rect 5632 7822 5684 7828
rect 5630 6896 5686 6905
rect 5630 6831 5686 6840
rect 5502 6446 5580 6474
rect 5446 6423 5502 6432
rect 5356 6394 5408 6400
rect 5448 6316 5500 6322
rect 5448 6258 5500 6264
rect 5354 5808 5410 5817
rect 5460 5778 5488 6258
rect 5540 6112 5592 6118
rect 5540 6054 5592 6060
rect 5552 5778 5580 6054
rect 5354 5743 5410 5752
rect 5448 5772 5500 5778
rect 5368 5710 5396 5743
rect 5448 5714 5500 5720
rect 5540 5772 5592 5778
rect 5540 5714 5592 5720
rect 5356 5704 5408 5710
rect 5356 5646 5408 5652
rect 5356 5568 5408 5574
rect 5356 5510 5408 5516
rect 5368 5302 5396 5510
rect 5356 5296 5408 5302
rect 5356 5238 5408 5244
rect 5368 5098 5396 5238
rect 5356 5092 5408 5098
rect 5356 5034 5408 5040
rect 5540 5024 5592 5030
rect 5540 4966 5592 4972
rect 5448 4616 5500 4622
rect 5448 4558 5500 4564
rect 5356 4480 5408 4486
rect 5356 4422 5408 4428
rect 5368 4146 5396 4422
rect 5172 4140 5224 4146
rect 5172 4082 5224 4088
rect 5264 4140 5316 4146
rect 5264 4082 5316 4088
rect 5356 4140 5408 4146
rect 5356 4082 5408 4088
rect 5172 3936 5224 3942
rect 5092 3896 5172 3924
rect 5172 3878 5224 3884
rect 5354 3904 5410 3913
rect 5354 3839 5410 3848
rect 5368 3398 5396 3839
rect 5460 3738 5488 4558
rect 5448 3732 5500 3738
rect 5448 3674 5500 3680
rect 5552 3534 5580 4966
rect 5540 3528 5592 3534
rect 5540 3470 5592 3476
rect 5356 3392 5408 3398
rect 5356 3334 5408 3340
rect 4894 3088 4950 3097
rect 4894 3023 4950 3032
rect 4896 2916 4948 2922
rect 4896 2858 4948 2864
rect 4724 2746 4844 2774
rect 4724 2650 4752 2746
rect 4712 2644 4764 2650
rect 4712 2586 4764 2592
rect 4908 2553 4936 2858
rect 4894 2544 4950 2553
rect 4712 2508 4764 2514
rect 4894 2479 4950 2488
rect 4712 2450 4764 2456
rect 4618 1320 4674 1329
rect 4618 1255 4674 1264
rect 4528 808 4580 814
rect 4528 750 4580 756
rect 4724 542 4752 2450
rect 4804 2440 4856 2446
rect 4804 2382 4856 2388
rect 4816 1834 4844 2382
rect 5540 2304 5592 2310
rect 5540 2246 5592 2252
rect 4804 1828 4856 1834
rect 4804 1770 4856 1776
rect 4712 536 4764 542
rect 4712 478 4764 484
rect 5552 56 5580 2246
rect 5644 513 5672 6831
rect 5736 5250 5764 11194
rect 5908 9580 5960 9586
rect 5908 9522 5960 9528
rect 5814 8936 5870 8945
rect 5814 8871 5870 8880
rect 5828 8634 5856 8871
rect 5816 8628 5868 8634
rect 5816 8570 5868 8576
rect 5920 8106 5948 9522
rect 6012 9042 6040 11194
rect 6092 9920 6144 9926
rect 6092 9862 6144 9868
rect 6000 9036 6052 9042
rect 6000 8978 6052 8984
rect 6104 8634 6132 9862
rect 6184 9852 6236 9858
rect 6184 9794 6236 9800
rect 6092 8628 6144 8634
rect 6092 8570 6144 8576
rect 6000 8492 6052 8498
rect 6000 8434 6052 8440
rect 5828 8078 5948 8106
rect 5828 6882 5856 8078
rect 5908 7880 5960 7886
rect 5908 7822 5960 7828
rect 5920 7410 5948 7822
rect 5908 7404 5960 7410
rect 5908 7346 5960 7352
rect 5828 6854 5948 6882
rect 5816 6792 5868 6798
rect 5816 6734 5868 6740
rect 5828 6497 5856 6734
rect 5814 6488 5870 6497
rect 5814 6423 5870 6432
rect 5828 5642 5856 6423
rect 5920 6322 5948 6854
rect 5908 6316 5960 6322
rect 5908 6258 5960 6264
rect 5908 5704 5960 5710
rect 5908 5646 5960 5652
rect 5816 5636 5868 5642
rect 5816 5578 5868 5584
rect 5920 5370 5948 5646
rect 5908 5364 5960 5370
rect 5908 5306 5960 5312
rect 5736 5222 5948 5250
rect 5816 5024 5868 5030
rect 5816 4966 5868 4972
rect 5724 4616 5776 4622
rect 5828 4604 5856 4966
rect 5776 4576 5856 4604
rect 5724 4558 5776 4564
rect 5816 4140 5868 4146
rect 5816 4082 5868 4088
rect 5828 3738 5856 4082
rect 5920 4010 5948 5222
rect 5908 4004 5960 4010
rect 5908 3946 5960 3952
rect 5816 3732 5868 3738
rect 5816 3674 5868 3680
rect 5908 3732 5960 3738
rect 5908 3674 5960 3680
rect 5920 2854 5948 3674
rect 5908 2848 5960 2854
rect 5908 2790 5960 2796
rect 6012 2650 6040 8434
rect 6092 8356 6144 8362
rect 6092 8298 6144 8304
rect 6104 5030 6132 8298
rect 6196 6458 6224 9794
rect 6184 6452 6236 6458
rect 6184 6394 6236 6400
rect 6288 5370 6316 11194
rect 6460 10192 6512 10198
rect 6460 10134 6512 10140
rect 6368 9648 6420 9654
rect 6368 9590 6420 9596
rect 6380 7449 6408 9590
rect 6366 7440 6422 7449
rect 6366 7375 6422 7384
rect 6368 7336 6420 7342
rect 6368 7278 6420 7284
rect 6380 5545 6408 7278
rect 6472 6458 6500 10134
rect 6564 9994 6592 11194
rect 6826 11194 6882 11250
rect 7102 11194 7158 11250
rect 7378 11194 7434 11250
rect 7654 11194 7710 11250
rect 7930 11194 7986 11250
rect 8206 11194 8262 11250
rect 8482 11194 8538 11250
rect 8758 11194 8814 11250
rect 9034 11194 9090 11250
rect 9310 11194 9366 11250
rect 9586 11194 9642 11250
rect 9862 11194 9918 11250
rect 10138 11194 10194 11250
rect 10414 11194 10470 11250
rect 10690 11194 10746 11250
rect 10966 11194 11022 11250
rect 11242 11194 11298 11250
rect 11518 11194 11574 11250
rect 11794 11194 11850 11250
rect 12070 11194 12126 11250
rect 12346 11194 12402 11250
rect 12622 11194 12678 11250
rect 12898 11212 12954 11250
rect 12898 11194 12900 11212
rect 6644 11154 6696 11160
rect 6552 9988 6604 9994
rect 6552 9930 6604 9936
rect 6656 8634 6684 11154
rect 6734 8800 6790 8809
rect 6734 8735 6790 8744
rect 6644 8628 6696 8634
rect 6644 8570 6696 8576
rect 6644 8288 6696 8294
rect 6644 8230 6696 8236
rect 6656 7818 6684 8230
rect 6644 7812 6696 7818
rect 6644 7754 6696 7760
rect 6552 7744 6604 7750
rect 6748 7698 6776 8735
rect 6552 7686 6604 7692
rect 6564 6866 6592 7686
rect 6656 7670 6776 7698
rect 6656 7410 6684 7670
rect 6840 7528 6868 11194
rect 7012 10124 7064 10130
rect 7012 10066 7064 10072
rect 6920 8968 6972 8974
rect 6920 8910 6972 8916
rect 6932 8090 6960 8910
rect 7024 8634 7052 10066
rect 7012 8628 7064 8634
rect 7012 8570 7064 8576
rect 6920 8084 6972 8090
rect 6920 8026 6972 8032
rect 7010 7984 7066 7993
rect 7010 7919 7066 7928
rect 6918 7848 6974 7857
rect 6918 7783 6974 7792
rect 6748 7500 6868 7528
rect 6644 7404 6696 7410
rect 6644 7346 6696 7352
rect 6552 6860 6604 6866
rect 6552 6802 6604 6808
rect 6460 6452 6512 6458
rect 6460 6394 6512 6400
rect 6644 6316 6696 6322
rect 6644 6258 6696 6264
rect 6460 6180 6512 6186
rect 6460 6122 6512 6128
rect 6366 5536 6422 5545
rect 6366 5471 6422 5480
rect 6276 5364 6328 5370
rect 6276 5306 6328 5312
rect 6184 5228 6236 5234
rect 6184 5170 6236 5176
rect 6276 5228 6328 5234
rect 6276 5170 6328 5176
rect 6092 5024 6144 5030
rect 6092 4966 6144 4972
rect 6092 4684 6144 4690
rect 6092 4626 6144 4632
rect 6104 4078 6132 4626
rect 6196 4185 6224 5170
rect 6288 4622 6316 5170
rect 6368 5092 6420 5098
rect 6368 5034 6420 5040
rect 6380 4690 6408 5034
rect 6472 4758 6500 6122
rect 6552 5568 6604 5574
rect 6552 5510 6604 5516
rect 6460 4752 6512 4758
rect 6460 4694 6512 4700
rect 6368 4684 6420 4690
rect 6368 4626 6420 4632
rect 6276 4616 6328 4622
rect 6276 4558 6328 4564
rect 6380 4282 6408 4626
rect 6368 4276 6420 4282
rect 6368 4218 6420 4224
rect 6182 4176 6238 4185
rect 6182 4111 6238 4120
rect 6564 4078 6592 5510
rect 6656 5273 6684 6258
rect 6748 5914 6776 7500
rect 6828 7404 6880 7410
rect 6828 7346 6880 7352
rect 6840 7041 6868 7346
rect 6826 7032 6882 7041
rect 6826 6967 6882 6976
rect 6932 6798 6960 7783
rect 7024 7478 7052 7919
rect 7012 7472 7064 7478
rect 7012 7414 7064 7420
rect 7010 7304 7066 7313
rect 7010 7239 7066 7248
rect 6920 6792 6972 6798
rect 6920 6734 6972 6740
rect 6828 6724 6880 6730
rect 6828 6666 6880 6672
rect 6840 6361 6868 6666
rect 6920 6656 6972 6662
rect 6920 6598 6972 6604
rect 6826 6352 6882 6361
rect 6826 6287 6882 6296
rect 6736 5908 6788 5914
rect 6736 5850 6788 5856
rect 6828 5364 6880 5370
rect 6828 5306 6880 5312
rect 6642 5264 6698 5273
rect 6642 5199 6698 5208
rect 6736 5092 6788 5098
rect 6736 5034 6788 5040
rect 6644 4548 6696 4554
rect 6644 4490 6696 4496
rect 6092 4072 6144 4078
rect 6092 4014 6144 4020
rect 6552 4072 6604 4078
rect 6552 4014 6604 4020
rect 6656 3670 6684 4490
rect 6644 3664 6696 3670
rect 6642 3632 6644 3641
rect 6696 3632 6698 3641
rect 6642 3567 6698 3576
rect 6184 2848 6236 2854
rect 6184 2790 6236 2796
rect 6000 2644 6052 2650
rect 6000 2586 6052 2592
rect 6196 2446 6224 2790
rect 5908 2440 5960 2446
rect 5908 2382 5960 2388
rect 6184 2440 6236 2446
rect 6184 2382 6236 2388
rect 5920 1902 5948 2382
rect 6644 2304 6696 2310
rect 6644 2246 6696 2252
rect 5908 1896 5960 1902
rect 5908 1838 5960 1844
rect 5630 504 5686 513
rect 5630 439 5686 448
rect 6656 56 6684 2246
rect 6748 1358 6776 5034
rect 6840 4486 6868 5306
rect 6828 4480 6880 4486
rect 6828 4422 6880 4428
rect 6932 4282 6960 6598
rect 7024 6458 7052 7239
rect 7116 6458 7144 11194
rect 7288 10396 7340 10402
rect 7288 10338 7340 10344
rect 7196 9716 7248 9722
rect 7196 9658 7248 9664
rect 7208 8634 7236 9658
rect 7196 8628 7248 8634
rect 7196 8570 7248 8576
rect 7194 8392 7250 8401
rect 7194 8327 7250 8336
rect 7208 7206 7236 8327
rect 7196 7200 7248 7206
rect 7196 7142 7248 7148
rect 7012 6452 7064 6458
rect 7012 6394 7064 6400
rect 7104 6452 7156 6458
rect 7104 6394 7156 6400
rect 7300 6322 7328 10338
rect 7104 6316 7156 6322
rect 7104 6258 7156 6264
rect 7288 6316 7340 6322
rect 7288 6258 7340 6264
rect 7010 5400 7066 5409
rect 7010 5335 7012 5344
rect 7064 5335 7066 5344
rect 7012 5306 7064 5312
rect 7012 5228 7064 5234
rect 7012 5170 7064 5176
rect 7024 4282 7052 5170
rect 6920 4276 6972 4282
rect 6920 4218 6972 4224
rect 7012 4276 7064 4282
rect 7012 4218 7064 4224
rect 7012 4140 7064 4146
rect 7012 4082 7064 4088
rect 6826 3224 6882 3233
rect 6826 3159 6828 3168
rect 6880 3159 6882 3168
rect 6828 3130 6880 3136
rect 6920 2984 6972 2990
rect 6920 2926 6972 2932
rect 6932 2854 6960 2926
rect 6920 2848 6972 2854
rect 6920 2790 6972 2796
rect 7024 2446 7052 4082
rect 7012 2440 7064 2446
rect 7012 2382 7064 2388
rect 7116 2009 7144 6258
rect 7286 6080 7342 6089
rect 7286 6015 7342 6024
rect 7196 5840 7248 5846
rect 7196 5782 7248 5788
rect 7300 5794 7328 6015
rect 7392 5914 7420 11194
rect 7668 10010 7696 11194
rect 7484 9982 7696 10010
rect 7840 10056 7892 10062
rect 7840 9998 7892 10004
rect 7484 8294 7512 9982
rect 7562 9888 7618 9897
rect 7562 9823 7618 9832
rect 7472 8288 7524 8294
rect 7472 8230 7524 8236
rect 7472 7336 7524 7342
rect 7472 7278 7524 7284
rect 7484 6390 7512 7278
rect 7576 6458 7604 9823
rect 7654 9480 7710 9489
rect 7654 9415 7710 9424
rect 7668 8498 7696 9415
rect 7748 8968 7800 8974
rect 7748 8910 7800 8916
rect 7760 8634 7788 8910
rect 7748 8628 7800 8634
rect 7748 8570 7800 8576
rect 7656 8492 7708 8498
rect 7656 8434 7708 8440
rect 7746 8256 7802 8265
rect 7746 8191 7802 8200
rect 7654 8120 7710 8129
rect 7654 8055 7710 8064
rect 7668 8022 7696 8055
rect 7656 8016 7708 8022
rect 7656 7958 7708 7964
rect 7760 7886 7788 8191
rect 7748 7880 7800 7886
rect 7748 7822 7800 7828
rect 7748 7744 7800 7750
rect 7748 7686 7800 7692
rect 7656 7404 7708 7410
rect 7656 7346 7708 7352
rect 7668 6662 7696 7346
rect 7760 7002 7788 7686
rect 7748 6996 7800 7002
rect 7748 6938 7800 6944
rect 7748 6724 7800 6730
rect 7748 6666 7800 6672
rect 7656 6656 7708 6662
rect 7656 6598 7708 6604
rect 7760 6458 7788 6666
rect 7564 6452 7616 6458
rect 7564 6394 7616 6400
rect 7748 6452 7800 6458
rect 7748 6394 7800 6400
rect 7472 6384 7524 6390
rect 7472 6326 7524 6332
rect 7380 5908 7432 5914
rect 7380 5850 7432 5856
rect 7208 3738 7236 5782
rect 7300 5766 7420 5794
rect 7288 5704 7340 5710
rect 7288 5646 7340 5652
rect 7196 3732 7248 3738
rect 7196 3674 7248 3680
rect 7196 3460 7248 3466
rect 7196 3402 7248 3408
rect 7208 3194 7236 3402
rect 7196 3188 7248 3194
rect 7196 3130 7248 3136
rect 7102 2000 7158 2009
rect 7102 1935 7158 1944
rect 6736 1352 6788 1358
rect 6736 1294 6788 1300
rect 7300 610 7328 5646
rect 7392 3534 7420 5766
rect 7484 5642 7512 6326
rect 7564 6316 7616 6322
rect 7564 6258 7616 6264
rect 7472 5636 7524 5642
rect 7472 5578 7524 5584
rect 7472 5024 7524 5030
rect 7472 4966 7524 4972
rect 7484 4214 7512 4966
rect 7472 4208 7524 4214
rect 7472 4150 7524 4156
rect 7470 3768 7526 3777
rect 7470 3703 7526 3712
rect 7484 3602 7512 3703
rect 7472 3596 7524 3602
rect 7472 3538 7524 3544
rect 7380 3528 7432 3534
rect 7380 3470 7432 3476
rect 7392 882 7420 3470
rect 7472 3052 7524 3058
rect 7472 2994 7524 3000
rect 7484 2446 7512 2994
rect 7472 2440 7524 2446
rect 7472 2382 7524 2388
rect 7576 2258 7604 6258
rect 7656 6248 7708 6254
rect 7656 6190 7708 6196
rect 7668 4010 7696 6190
rect 7760 6186 7788 6394
rect 7748 6180 7800 6186
rect 7748 6122 7800 6128
rect 7852 5914 7880 9998
rect 7944 9858 7972 11194
rect 8220 10305 8248 11194
rect 8206 10296 8262 10305
rect 8206 10231 8262 10240
rect 8392 9988 8444 9994
rect 8392 9930 8444 9936
rect 7932 9852 7984 9858
rect 7932 9794 7984 9800
rect 7930 9752 7986 9761
rect 7930 9687 7986 9696
rect 7944 8362 7972 9687
rect 8024 9036 8076 9042
rect 8024 8978 8076 8984
rect 8036 8537 8064 8978
rect 8116 8900 8168 8906
rect 8116 8842 8168 8848
rect 8022 8528 8078 8537
rect 8128 8498 8156 8842
rect 8404 8634 8432 9930
rect 8496 9674 8524 11194
rect 8772 10198 8800 11194
rect 9048 10418 9076 11194
rect 9324 10441 9352 11194
rect 8864 10390 9076 10418
rect 9310 10432 9366 10441
rect 8760 10192 8812 10198
rect 8760 10134 8812 10140
rect 8576 9784 8628 9790
rect 8576 9726 8628 9732
rect 8588 9674 8616 9726
rect 8496 9646 8533 9674
rect 8505 9602 8533 9646
rect 8496 9574 8533 9602
rect 8568 9646 8616 9674
rect 8568 9602 8596 9646
rect 8568 9574 8616 9602
rect 8392 8628 8444 8634
rect 8392 8570 8444 8576
rect 8022 8463 8078 8472
rect 8116 8492 8168 8498
rect 8116 8434 8168 8440
rect 8392 8424 8444 8430
rect 8312 8384 8392 8412
rect 7932 8356 7984 8362
rect 7932 8298 7984 8304
rect 7950 8188 8258 8197
rect 7950 8186 7956 8188
rect 8012 8186 8036 8188
rect 8092 8186 8116 8188
rect 8172 8186 8196 8188
rect 8252 8186 8258 8188
rect 8012 8134 8014 8186
rect 8194 8134 8196 8186
rect 7950 8132 7956 8134
rect 8012 8132 8036 8134
rect 8092 8132 8116 8134
rect 8172 8132 8196 8134
rect 8252 8132 8258 8134
rect 7950 8123 8258 8132
rect 7932 7948 7984 7954
rect 7932 7890 7984 7896
rect 7944 7449 7972 7890
rect 8116 7880 8168 7886
rect 8116 7822 8168 7828
rect 7930 7440 7986 7449
rect 7930 7375 7986 7384
rect 7932 7268 7984 7274
rect 8128 7256 8156 7822
rect 8312 7410 8340 8384
rect 8392 8366 8444 8372
rect 8392 8288 8444 8294
rect 8390 8256 8392 8265
rect 8444 8256 8446 8265
rect 8390 8191 8446 8200
rect 8392 7880 8444 7886
rect 8392 7822 8444 7828
rect 8404 7478 8432 7822
rect 8392 7472 8444 7478
rect 8392 7414 8444 7420
rect 8300 7404 8352 7410
rect 8300 7346 8352 7352
rect 8496 7313 8524 9574
rect 8588 8634 8616 9574
rect 8864 9364 8892 10390
rect 9310 10367 9366 10376
rect 8944 10328 8996 10334
rect 8944 10270 8996 10276
rect 9402 10296 9458 10305
rect 8956 9654 8984 10270
rect 9402 10231 9458 10240
rect 9496 10260 9548 10266
rect 8944 9648 8996 9654
rect 8944 9590 8996 9596
rect 9036 9648 9088 9654
rect 9036 9590 9088 9596
rect 8680 9336 8892 9364
rect 8576 8628 8628 8634
rect 8576 8570 8628 8576
rect 8680 8378 8708 9336
rect 8852 8968 8904 8974
rect 8772 8928 8852 8956
rect 8772 8498 8800 8928
rect 8852 8910 8904 8916
rect 9048 8838 9076 9590
rect 9036 8832 9088 8838
rect 9416 8809 9444 10231
rect 9496 10202 9548 10208
rect 9036 8774 9088 8780
rect 9402 8800 9458 8809
rect 9010 8732 9318 8741
rect 9402 8735 9458 8744
rect 9010 8730 9016 8732
rect 9072 8730 9096 8732
rect 9152 8730 9176 8732
rect 9232 8730 9256 8732
rect 9312 8730 9318 8732
rect 9072 8678 9074 8730
rect 9254 8678 9256 8730
rect 9010 8676 9016 8678
rect 9072 8676 9096 8678
rect 9152 8676 9176 8678
rect 9232 8676 9256 8678
rect 9312 8676 9318 8678
rect 9010 8667 9318 8676
rect 9508 8650 9536 10202
rect 9600 10062 9628 11194
rect 9588 10056 9640 10062
rect 9588 9998 9640 10004
rect 9876 9897 9904 11194
rect 10046 10704 10102 10713
rect 10046 10639 10102 10648
rect 10060 9897 10088 10639
rect 9862 9888 9918 9897
rect 9588 9852 9640 9858
rect 9862 9823 9918 9832
rect 10046 9888 10102 9897
rect 10046 9823 10102 9832
rect 9588 9794 9640 9800
rect 9416 8622 9536 8650
rect 9600 8634 9628 9794
rect 9772 9512 9824 9518
rect 9772 9454 9824 9460
rect 9864 9512 9916 9518
rect 9864 9454 9916 9460
rect 9680 9172 9732 9178
rect 9680 9114 9732 9120
rect 9588 8628 9640 8634
rect 8760 8492 8812 8498
rect 8760 8434 8812 8440
rect 8944 8424 8996 8430
rect 8680 8350 8892 8378
rect 8944 8366 8996 8372
rect 9220 8424 9272 8430
rect 9272 8384 9352 8412
rect 9220 8366 9272 8372
rect 8760 8288 8812 8294
rect 8666 8256 8722 8265
rect 8760 8230 8812 8236
rect 8666 8191 8722 8200
rect 8574 7984 8630 7993
rect 8574 7919 8630 7928
rect 8588 7721 8616 7919
rect 8574 7712 8630 7721
rect 8574 7647 8630 7656
rect 8680 7585 8708 8191
rect 8666 7576 8722 7585
rect 8666 7511 8722 7520
rect 8772 7460 8800 8230
rect 8864 7546 8892 8350
rect 8956 7954 8984 8366
rect 9324 8106 9352 8384
rect 9416 8294 9444 8622
rect 9588 8570 9640 8576
rect 9496 8560 9548 8566
rect 9692 8514 9720 9114
rect 9496 8502 9548 8508
rect 9404 8288 9456 8294
rect 9404 8230 9456 8236
rect 9324 8078 9444 8106
rect 8944 7948 8996 7954
rect 8944 7890 8996 7896
rect 8956 7818 8984 7890
rect 8944 7812 8996 7818
rect 8944 7754 8996 7760
rect 9010 7644 9318 7653
rect 9010 7642 9016 7644
rect 9072 7642 9096 7644
rect 9152 7642 9176 7644
rect 9232 7642 9256 7644
rect 9312 7642 9318 7644
rect 9072 7590 9074 7642
rect 9254 7590 9256 7642
rect 9010 7588 9016 7590
rect 9072 7588 9096 7590
rect 9152 7588 9176 7590
rect 9232 7588 9256 7590
rect 9312 7588 9318 7590
rect 9010 7579 9318 7588
rect 8852 7540 8904 7546
rect 8852 7482 8904 7488
rect 8588 7432 8800 7460
rect 8482 7304 8538 7313
rect 7984 7228 8351 7256
rect 8482 7239 8538 7248
rect 7932 7210 7984 7216
rect 8323 7154 8351 7228
rect 8588 7188 8616 7432
rect 8852 7404 8904 7410
rect 8852 7346 8904 7352
rect 8312 7126 8351 7154
rect 8404 7160 8616 7188
rect 8668 7200 8720 7206
rect 7950 7100 8258 7109
rect 7950 7098 7956 7100
rect 8012 7098 8036 7100
rect 8092 7098 8116 7100
rect 8172 7098 8196 7100
rect 8252 7098 8258 7100
rect 8012 7046 8014 7098
rect 8194 7046 8196 7098
rect 7950 7044 7956 7046
rect 8012 7044 8036 7046
rect 8092 7044 8116 7046
rect 8172 7044 8196 7046
rect 8252 7044 8258 7046
rect 7950 7035 8258 7044
rect 8312 6848 8340 7126
rect 8036 6820 8340 6848
rect 8036 6186 8064 6820
rect 8116 6724 8168 6730
rect 8116 6666 8168 6672
rect 8128 6390 8156 6666
rect 8116 6384 8168 6390
rect 8116 6326 8168 6332
rect 8116 6248 8168 6254
rect 8168 6208 8340 6236
rect 8116 6190 8168 6196
rect 8024 6180 8076 6186
rect 8024 6122 8076 6128
rect 7950 6012 8258 6021
rect 7950 6010 7956 6012
rect 8012 6010 8036 6012
rect 8092 6010 8116 6012
rect 8172 6010 8196 6012
rect 8252 6010 8258 6012
rect 8012 5958 8014 6010
rect 8194 5958 8196 6010
rect 7950 5956 7956 5958
rect 8012 5956 8036 5958
rect 8092 5956 8116 5958
rect 8172 5956 8196 5958
rect 8252 5956 8258 5958
rect 7950 5947 8258 5956
rect 7840 5908 7892 5914
rect 7840 5850 7892 5856
rect 8312 5574 8340 6208
rect 8404 5914 8432 7160
rect 8668 7142 8720 7148
rect 8482 6896 8538 6905
rect 8680 6848 8708 7142
rect 8864 6934 8892 7346
rect 8852 6928 8904 6934
rect 8852 6870 8904 6876
rect 8482 6831 8538 6840
rect 8496 6633 8524 6831
rect 8588 6820 8708 6848
rect 8482 6624 8538 6633
rect 8482 6559 8538 6568
rect 8392 5908 8444 5914
rect 8392 5850 8444 5856
rect 8300 5568 8352 5574
rect 8300 5510 8352 5516
rect 7840 5228 7892 5234
rect 7840 5170 7892 5176
rect 7852 4826 7880 5170
rect 7950 4924 8258 4933
rect 7950 4922 7956 4924
rect 8012 4922 8036 4924
rect 8092 4922 8116 4924
rect 8172 4922 8196 4924
rect 8252 4922 8258 4924
rect 8012 4870 8014 4922
rect 8194 4870 8196 4922
rect 7950 4868 7956 4870
rect 8012 4868 8036 4870
rect 8092 4868 8116 4870
rect 8172 4868 8196 4870
rect 8252 4868 8258 4870
rect 7950 4859 8258 4868
rect 7840 4820 7892 4826
rect 7840 4762 7892 4768
rect 7748 4752 7800 4758
rect 7746 4720 7748 4729
rect 7800 4720 7802 4729
rect 8312 4672 8340 5510
rect 8390 5400 8446 5409
rect 8390 5335 8446 5344
rect 8404 4758 8432 5335
rect 8484 5160 8536 5166
rect 8484 5102 8536 5108
rect 8496 4865 8524 5102
rect 8482 4856 8538 4865
rect 8482 4791 8538 4800
rect 8392 4752 8444 4758
rect 8392 4694 8444 4700
rect 7746 4655 7802 4664
rect 8220 4644 8340 4672
rect 8116 4616 8168 4622
rect 8116 4558 8168 4564
rect 8128 4146 8156 4558
rect 8116 4140 8168 4146
rect 8116 4082 8168 4088
rect 7656 4004 7708 4010
rect 7656 3946 7708 3952
rect 8220 3924 8248 4644
rect 8588 4570 8616 6820
rect 8852 6792 8904 6798
rect 8852 6734 8904 6740
rect 8668 6724 8720 6730
rect 8668 6666 8720 6672
rect 8680 6322 8708 6666
rect 8758 6488 8814 6497
rect 8758 6423 8760 6432
rect 8812 6423 8814 6432
rect 8760 6394 8812 6400
rect 8668 6316 8720 6322
rect 8668 6258 8720 6264
rect 8760 6316 8812 6322
rect 8760 6258 8812 6264
rect 8668 5636 8720 5642
rect 8668 5578 8720 5584
rect 8312 4542 8616 4570
rect 8312 4214 8340 4542
rect 8576 4480 8628 4486
rect 8576 4422 8628 4428
rect 8588 4282 8616 4422
rect 8576 4276 8628 4282
rect 8576 4218 8628 4224
rect 8300 4208 8352 4214
rect 8300 4150 8352 4156
rect 8680 4126 8708 5578
rect 8496 4098 8708 4126
rect 8392 4072 8444 4078
rect 8392 4014 8444 4020
rect 8220 3896 8340 3924
rect 7950 3836 8258 3845
rect 7950 3834 7956 3836
rect 8012 3834 8036 3836
rect 8092 3834 8116 3836
rect 8172 3834 8196 3836
rect 8252 3834 8258 3836
rect 8012 3782 8014 3834
rect 8194 3782 8196 3834
rect 7950 3780 7956 3782
rect 8012 3780 8036 3782
rect 8092 3780 8116 3782
rect 8172 3780 8196 3782
rect 8252 3780 8258 3782
rect 7950 3771 8258 3780
rect 7656 3596 7708 3602
rect 7656 3538 7708 3544
rect 7668 3369 7696 3538
rect 8312 3534 8340 3896
rect 8404 3738 8432 4014
rect 8392 3732 8444 3738
rect 8392 3674 8444 3680
rect 8300 3528 8352 3534
rect 8300 3470 8352 3476
rect 8496 3448 8524 4098
rect 8576 4004 8628 4010
rect 8772 3992 8800 6258
rect 8864 5778 8892 6734
rect 9010 6556 9318 6565
rect 9010 6554 9016 6556
rect 9072 6554 9096 6556
rect 9152 6554 9176 6556
rect 9232 6554 9256 6556
rect 9312 6554 9318 6556
rect 9072 6502 9074 6554
rect 9254 6502 9256 6554
rect 9010 6500 9016 6502
rect 9072 6500 9096 6502
rect 9152 6500 9176 6502
rect 9232 6500 9256 6502
rect 9312 6500 9318 6502
rect 9010 6491 9318 6500
rect 9036 6384 9088 6390
rect 8956 6344 9036 6372
rect 8852 5772 8904 5778
rect 8852 5714 8904 5720
rect 8956 5658 8984 6344
rect 9036 6326 9088 6332
rect 9128 6316 9180 6322
rect 9128 6258 9180 6264
rect 9140 6089 9168 6258
rect 9416 6254 9444 8078
rect 9508 7546 9536 8502
rect 9600 8486 9720 8514
rect 9600 8430 9628 8486
rect 9588 8424 9640 8430
rect 9588 8366 9640 8372
rect 9784 8294 9812 9454
rect 9772 8288 9824 8294
rect 9772 8230 9824 8236
rect 9680 7812 9732 7818
rect 9680 7754 9732 7760
rect 9496 7540 9548 7546
rect 9496 7482 9548 7488
rect 9692 7478 9720 7754
rect 9680 7472 9732 7478
rect 9600 7432 9680 7460
rect 9496 7200 9548 7206
rect 9496 7142 9548 7148
rect 9508 6390 9536 7142
rect 9600 6798 9628 7432
rect 9680 7414 9732 7420
rect 9680 7336 9732 7342
rect 9680 7278 9732 7284
rect 9692 6798 9720 7278
rect 9588 6792 9640 6798
rect 9588 6734 9640 6740
rect 9680 6792 9732 6798
rect 9680 6734 9732 6740
rect 9496 6384 9548 6390
rect 9496 6326 9548 6332
rect 9586 6352 9642 6361
rect 9586 6287 9588 6296
rect 9640 6287 9642 6296
rect 9588 6258 9640 6264
rect 9404 6248 9456 6254
rect 9404 6190 9456 6196
rect 9126 6080 9182 6089
rect 9126 6015 9182 6024
rect 9494 6080 9550 6089
rect 9494 6015 9550 6024
rect 9312 5908 9364 5914
rect 9312 5850 9364 5856
rect 8628 3964 8800 3992
rect 8864 5630 8984 5658
rect 8576 3946 8628 3952
rect 8864 3913 8892 5630
rect 9324 5556 9352 5850
rect 9324 5528 9444 5556
rect 9010 5468 9318 5477
rect 9010 5466 9016 5468
rect 9072 5466 9096 5468
rect 9152 5466 9176 5468
rect 9232 5466 9256 5468
rect 9312 5466 9318 5468
rect 9072 5414 9074 5466
rect 9254 5414 9256 5466
rect 9010 5412 9016 5414
rect 9072 5412 9096 5414
rect 9152 5412 9176 5414
rect 9232 5412 9256 5414
rect 9312 5412 9318 5414
rect 9010 5403 9318 5412
rect 8944 5364 8996 5370
rect 9416 5352 9444 5528
rect 8996 5324 9168 5352
rect 8944 5306 8996 5312
rect 9140 5234 9168 5324
rect 9324 5324 9444 5352
rect 9036 5228 9088 5234
rect 9036 5170 9088 5176
rect 9128 5228 9180 5234
rect 9128 5170 9180 5176
rect 9048 4690 9076 5170
rect 9324 4690 9352 5324
rect 9508 4978 9536 6015
rect 9680 5704 9732 5710
rect 9416 4950 9536 4978
rect 9600 5664 9680 5692
rect 9416 4826 9444 4950
rect 9494 4856 9550 4865
rect 9404 4820 9456 4826
rect 9494 4791 9496 4800
rect 9404 4762 9456 4768
rect 9548 4791 9550 4800
rect 9496 4762 9548 4768
rect 9508 4690 9536 4762
rect 9036 4684 9088 4690
rect 9036 4626 9088 4632
rect 9312 4684 9364 4690
rect 9312 4626 9364 4632
rect 9496 4684 9548 4690
rect 9496 4626 9548 4632
rect 9010 4380 9318 4389
rect 9010 4378 9016 4380
rect 9072 4378 9096 4380
rect 9152 4378 9176 4380
rect 9232 4378 9256 4380
rect 9312 4378 9318 4380
rect 9072 4326 9074 4378
rect 9254 4326 9256 4378
rect 9010 4324 9016 4326
rect 9072 4324 9096 4326
rect 9152 4324 9176 4326
rect 9232 4324 9256 4326
rect 9312 4324 9318 4326
rect 9010 4315 9318 4324
rect 8944 4138 8996 4144
rect 8944 4080 8996 4086
rect 9220 4140 9272 4146
rect 9496 4140 9548 4146
rect 9272 4100 9352 4128
rect 9220 4082 9272 4088
rect 8956 3942 8984 4080
rect 9036 4004 9088 4010
rect 9220 4004 9272 4010
rect 9088 3964 9220 3992
rect 9036 3946 9088 3952
rect 9220 3946 9272 3952
rect 8944 3936 8996 3942
rect 8850 3904 8906 3913
rect 9324 3890 9352 4100
rect 9600 4128 9628 5664
rect 9680 5646 9732 5652
rect 9680 5364 9732 5370
rect 9680 5306 9732 5312
rect 9548 4100 9628 4128
rect 9496 4082 9548 4088
rect 9588 3936 9640 3942
rect 8944 3878 8996 3884
rect 8850 3839 8906 3848
rect 9232 3862 9352 3890
rect 9402 3904 9458 3913
rect 9036 3732 9088 3738
rect 8864 3692 9036 3720
rect 8496 3420 8708 3448
rect 7748 3392 7800 3398
rect 7654 3360 7710 3369
rect 7748 3334 7800 3340
rect 8482 3360 8538 3369
rect 7654 3295 7710 3304
rect 7760 3058 7788 3334
rect 8482 3295 8538 3304
rect 8496 3194 8524 3295
rect 7932 3188 7984 3194
rect 7932 3130 7984 3136
rect 8484 3188 8536 3194
rect 8484 3130 8536 3136
rect 7944 3058 7972 3130
rect 7748 3052 7800 3058
rect 7748 2994 7800 3000
rect 7932 3052 7984 3058
rect 7932 2994 7984 3000
rect 8496 2990 8524 3130
rect 8576 3052 8628 3058
rect 8576 2994 8628 3000
rect 8484 2984 8536 2990
rect 8484 2926 8536 2932
rect 7950 2748 8258 2757
rect 7950 2746 7956 2748
rect 8012 2746 8036 2748
rect 8092 2746 8116 2748
rect 8172 2746 8196 2748
rect 8252 2746 8258 2748
rect 8012 2694 8014 2746
rect 8194 2694 8196 2746
rect 7950 2692 7956 2694
rect 8012 2692 8036 2694
rect 8092 2692 8116 2694
rect 8172 2692 8196 2694
rect 8252 2692 8258 2694
rect 7950 2683 8258 2692
rect 8588 2446 8616 2994
rect 8680 2689 8708 3420
rect 8864 3233 8892 3692
rect 9036 3674 9088 3680
rect 9232 3534 9260 3862
rect 9586 3904 9588 3913
rect 9640 3904 9642 3913
rect 9458 3862 9536 3890
rect 9402 3839 9458 3848
rect 9310 3632 9366 3641
rect 9310 3567 9366 3576
rect 9324 3534 9352 3567
rect 9220 3528 9272 3534
rect 9220 3470 9272 3476
rect 9312 3528 9364 3534
rect 9312 3470 9364 3476
rect 9508 3398 9536 3862
rect 9586 3839 9642 3848
rect 9692 3602 9720 5306
rect 9784 4214 9812 8230
rect 9876 5234 9904 9454
rect 10152 9081 10180 11194
rect 10232 10124 10284 10130
rect 10232 10066 10284 10072
rect 10138 9072 10194 9081
rect 10138 9007 10194 9016
rect 9956 8424 10008 8430
rect 9956 8366 10008 8372
rect 9968 7206 9996 8366
rect 10244 7528 10272 10066
rect 10324 9376 10376 9382
rect 10324 9318 10376 9324
rect 10336 8498 10364 9318
rect 10324 8492 10376 8498
rect 10324 8434 10376 8440
rect 10324 7744 10376 7750
rect 10324 7686 10376 7692
rect 10336 7585 10364 7686
rect 10060 7500 10272 7528
rect 10322 7576 10378 7585
rect 10322 7511 10378 7520
rect 9956 7200 10008 7206
rect 9956 7142 10008 7148
rect 9864 5228 9916 5234
rect 9864 5170 9916 5176
rect 9864 5024 9916 5030
rect 9864 4966 9916 4972
rect 9956 5024 10008 5030
rect 9956 4966 10008 4972
rect 9772 4208 9824 4214
rect 9772 4150 9824 4156
rect 9876 4078 9904 4966
rect 9968 4554 9996 4966
rect 9956 4548 10008 4554
rect 9956 4490 10008 4496
rect 9954 4448 10010 4457
rect 10060 4434 10088 7500
rect 10428 7426 10456 11194
rect 10704 10577 10732 11194
rect 10690 10568 10746 10577
rect 10690 10503 10746 10512
rect 10874 10568 10930 10577
rect 10874 10503 10930 10512
rect 10784 9444 10836 9450
rect 10784 9386 10836 9392
rect 10508 9376 10560 9382
rect 10506 9344 10508 9353
rect 10560 9344 10562 9353
rect 10506 9279 10562 9288
rect 10598 8664 10654 8673
rect 10598 8599 10654 8608
rect 10508 8288 10560 8294
rect 10508 8230 10560 8236
rect 10520 7886 10548 8230
rect 10612 7886 10640 8599
rect 10796 8294 10824 9386
rect 10784 8288 10836 8294
rect 10888 8265 10916 10503
rect 10980 8945 11008 11194
rect 11256 10305 11284 11194
rect 11242 10296 11298 10305
rect 11242 10231 11298 10240
rect 11336 9172 11388 9178
rect 11336 9114 11388 9120
rect 10966 8936 11022 8945
rect 10966 8871 11022 8880
rect 11244 8628 11296 8634
rect 11244 8570 11296 8576
rect 10968 8492 11020 8498
rect 10968 8434 11020 8440
rect 10784 8230 10836 8236
rect 10874 8256 10930 8265
rect 10508 7880 10560 7886
rect 10508 7822 10560 7828
rect 10600 7880 10652 7886
rect 10600 7822 10652 7828
rect 10600 7540 10652 7546
rect 10600 7482 10652 7488
rect 10244 7398 10456 7426
rect 10508 7472 10560 7478
rect 10508 7414 10560 7420
rect 10140 6656 10192 6662
rect 10140 6598 10192 6604
rect 10152 6322 10180 6598
rect 10140 6316 10192 6322
rect 10140 6258 10192 6264
rect 10244 6118 10272 7398
rect 10324 7200 10376 7206
rect 10324 7142 10376 7148
rect 10336 6118 10364 7142
rect 10520 6458 10548 7414
rect 10612 6798 10640 7482
rect 10600 6792 10652 6798
rect 10600 6734 10652 6740
rect 10692 6792 10744 6798
rect 10692 6734 10744 6740
rect 10600 6656 10652 6662
rect 10600 6598 10652 6604
rect 10508 6452 10560 6458
rect 10508 6394 10560 6400
rect 10416 6384 10468 6390
rect 10416 6326 10468 6332
rect 10232 6112 10284 6118
rect 10232 6054 10284 6060
rect 10324 6112 10376 6118
rect 10324 6054 10376 6060
rect 10428 5914 10456 6326
rect 10416 5908 10468 5914
rect 10416 5850 10468 5856
rect 10324 5636 10376 5642
rect 10324 5578 10376 5584
rect 10336 5234 10364 5578
rect 10324 5228 10376 5234
rect 10324 5170 10376 5176
rect 10416 5228 10468 5234
rect 10416 5170 10468 5176
rect 10232 5092 10284 5098
rect 10232 5034 10284 5040
rect 10244 4865 10272 5034
rect 10230 4856 10286 4865
rect 10230 4791 10286 4800
rect 10060 4406 10180 4434
rect 9954 4383 10010 4392
rect 9968 4282 9996 4383
rect 9956 4276 10008 4282
rect 9956 4218 10008 4224
rect 10048 4276 10100 4282
rect 10048 4218 10100 4224
rect 10060 4146 10088 4218
rect 10048 4140 10100 4146
rect 10048 4082 10100 4088
rect 9864 4072 9916 4078
rect 9864 4014 9916 4020
rect 9772 4004 9824 4010
rect 9772 3946 9824 3952
rect 9784 3641 9812 3946
rect 10152 3738 10180 4406
rect 10428 4282 10456 5170
rect 10506 4992 10562 5001
rect 10506 4927 10562 4936
rect 10416 4276 10468 4282
rect 10416 4218 10468 4224
rect 10140 3732 10192 3738
rect 10140 3674 10192 3680
rect 9770 3632 9826 3641
rect 9680 3596 9732 3602
rect 9770 3567 9826 3576
rect 9680 3538 9732 3544
rect 9954 3496 10010 3505
rect 9954 3431 10010 3440
rect 9312 3392 9364 3398
rect 9496 3392 9548 3398
rect 9364 3352 9444 3380
rect 9312 3334 9364 3340
rect 9010 3292 9318 3301
rect 9010 3290 9016 3292
rect 9072 3290 9096 3292
rect 9152 3290 9176 3292
rect 9232 3290 9256 3292
rect 9312 3290 9318 3292
rect 9072 3238 9074 3290
rect 9254 3238 9256 3290
rect 9010 3236 9016 3238
rect 9072 3236 9096 3238
rect 9152 3236 9176 3238
rect 9232 3236 9256 3238
rect 9312 3236 9318 3238
rect 8850 3224 8906 3233
rect 9010 3227 9318 3236
rect 9416 3233 9444 3352
rect 9496 3334 9548 3340
rect 8850 3159 8906 3168
rect 9402 3224 9458 3233
rect 9402 3159 9458 3168
rect 9036 2848 9088 2854
rect 9036 2790 9088 2796
rect 8666 2680 8722 2689
rect 8666 2615 8722 2624
rect 9048 2514 9076 2790
rect 9508 2514 9536 3334
rect 9968 3194 9996 3431
rect 10232 3392 10284 3398
rect 10232 3334 10284 3340
rect 10324 3392 10376 3398
rect 10324 3334 10376 3340
rect 9956 3188 10008 3194
rect 9956 3130 10008 3136
rect 10140 3188 10192 3194
rect 10140 3130 10192 3136
rect 9772 3052 9824 3058
rect 9772 2994 9824 3000
rect 9036 2508 9088 2514
rect 9036 2450 9088 2456
rect 9496 2508 9548 2514
rect 9496 2450 9548 2456
rect 8576 2440 8628 2446
rect 8576 2382 8628 2388
rect 7656 2372 7708 2378
rect 7656 2314 7708 2320
rect 8760 2372 8812 2378
rect 8760 2314 8812 2320
rect 9496 2372 9548 2378
rect 9496 2314 9548 2320
rect 7484 2230 7604 2258
rect 7380 876 7432 882
rect 7380 818 7432 824
rect 7484 746 7512 2230
rect 7564 2100 7616 2106
rect 7564 2042 7616 2048
rect 7576 1154 7604 2042
rect 7668 1562 7696 2314
rect 7748 2304 7800 2310
rect 7748 2246 7800 2252
rect 8576 2304 8628 2310
rect 8576 2246 8628 2252
rect 7656 1556 7708 1562
rect 7656 1498 7708 1504
rect 7564 1148 7616 1154
rect 7564 1090 7616 1096
rect 7472 740 7524 746
rect 7472 682 7524 688
rect 7288 604 7340 610
rect 7288 546 7340 552
rect 7760 56 7788 2246
rect 1122 0 1178 56
rect 2226 0 2282 56
rect 3330 0 3386 56
rect 4434 0 4490 56
rect 5538 0 5594 56
rect 6642 0 6698 56
rect 7746 0 7802 56
rect 8588 42 8616 2246
rect 8772 950 8800 2314
rect 9010 2204 9318 2213
rect 9010 2202 9016 2204
rect 9072 2202 9096 2204
rect 9152 2202 9176 2204
rect 9232 2202 9256 2204
rect 9312 2202 9318 2204
rect 9072 2150 9074 2202
rect 9254 2150 9256 2202
rect 9010 2148 9016 2150
rect 9072 2148 9096 2150
rect 9152 2148 9176 2150
rect 9232 2148 9256 2150
rect 9312 2148 9318 2150
rect 9010 2139 9318 2148
rect 9508 2106 9536 2314
rect 9784 2310 9812 2994
rect 10152 2990 10180 3130
rect 10140 2984 10192 2990
rect 10140 2926 10192 2932
rect 10140 2440 10192 2446
rect 10140 2382 10192 2388
rect 9588 2304 9640 2310
rect 9588 2246 9640 2252
rect 9772 2304 9824 2310
rect 9772 2246 9824 2252
rect 9956 2304 10008 2310
rect 9956 2246 10008 2252
rect 9496 2100 9548 2106
rect 9496 2042 9548 2048
rect 9600 1601 9628 2246
rect 9586 1592 9642 1601
rect 9586 1527 9642 1536
rect 8760 944 8812 950
rect 8760 886 8812 892
rect 8772 56 8892 82
rect 9968 56 9996 2246
rect 10152 1698 10180 2382
rect 10140 1692 10192 1698
rect 10140 1634 10192 1640
rect 10244 1018 10272 3334
rect 10336 2582 10364 3334
rect 10520 3058 10548 4927
rect 10612 4146 10640 6598
rect 10704 6458 10732 6734
rect 10692 6452 10744 6458
rect 10692 6394 10744 6400
rect 10692 6180 10744 6186
rect 10692 6122 10744 6128
rect 10704 5914 10732 6122
rect 10692 5908 10744 5914
rect 10692 5850 10744 5856
rect 10692 5296 10744 5302
rect 10692 5238 10744 5244
rect 10704 4486 10732 5238
rect 10796 4690 10824 8230
rect 10874 8191 10930 8200
rect 10876 7540 10928 7546
rect 10876 7482 10928 7488
rect 10888 6934 10916 7482
rect 10876 6928 10928 6934
rect 10876 6870 10928 6876
rect 10876 6724 10928 6730
rect 10876 6666 10928 6672
rect 10888 6458 10916 6666
rect 10876 6452 10928 6458
rect 10876 6394 10928 6400
rect 10876 6112 10928 6118
rect 10876 6054 10928 6060
rect 10888 5846 10916 6054
rect 10876 5840 10928 5846
rect 10876 5782 10928 5788
rect 10784 4684 10836 4690
rect 10784 4626 10836 4632
rect 10692 4480 10744 4486
rect 10692 4422 10744 4428
rect 10600 4140 10652 4146
rect 10600 4082 10652 4088
rect 10600 3528 10652 3534
rect 10600 3470 10652 3476
rect 10612 3058 10640 3470
rect 10508 3052 10560 3058
rect 10508 2994 10560 3000
rect 10600 3052 10652 3058
rect 10600 2994 10652 3000
rect 10324 2576 10376 2582
rect 10324 2518 10376 2524
rect 10324 2440 10376 2446
rect 10324 2382 10376 2388
rect 10336 2281 10364 2382
rect 10322 2272 10378 2281
rect 10322 2207 10378 2216
rect 10520 2145 10548 2994
rect 10598 2816 10654 2825
rect 10598 2751 10654 2760
rect 10612 2446 10640 2751
rect 10600 2440 10652 2446
rect 10600 2382 10652 2388
rect 10506 2136 10562 2145
rect 10704 2106 10732 4422
rect 10782 4312 10838 4321
rect 10782 4247 10838 4256
rect 10796 4214 10824 4247
rect 10784 4208 10836 4214
rect 10784 4150 10836 4156
rect 10784 4072 10836 4078
rect 10784 4014 10836 4020
rect 10796 3738 10824 4014
rect 10980 3942 11008 8434
rect 11256 8430 11284 8570
rect 11244 8424 11296 8430
rect 11244 8366 11296 8372
rect 11060 8288 11112 8294
rect 11060 8230 11112 8236
rect 11072 8090 11100 8230
rect 11060 8084 11112 8090
rect 11060 8026 11112 8032
rect 11152 8084 11204 8090
rect 11152 8026 11204 8032
rect 11060 7812 11112 7818
rect 11060 7754 11112 7760
rect 11072 7002 11100 7754
rect 11060 6996 11112 7002
rect 11060 6938 11112 6944
rect 11164 6798 11192 8026
rect 11348 6984 11376 9114
rect 11428 8424 11480 8430
rect 11428 8366 11480 8372
rect 11440 7206 11468 8366
rect 11532 8362 11560 11194
rect 11808 9926 11836 11194
rect 11796 9920 11848 9926
rect 11796 9862 11848 9868
rect 11888 9920 11940 9926
rect 11888 9862 11940 9868
rect 11796 9580 11848 9586
rect 11796 9522 11848 9528
rect 11808 9246 11836 9522
rect 11704 9240 11756 9246
rect 11704 9182 11756 9188
rect 11796 9240 11848 9246
rect 11796 9182 11848 9188
rect 11612 8628 11664 8634
rect 11612 8570 11664 8576
rect 11520 8356 11572 8362
rect 11520 8298 11572 8304
rect 11520 7336 11572 7342
rect 11520 7278 11572 7284
rect 11428 7200 11480 7206
rect 11428 7142 11480 7148
rect 11256 6956 11376 6984
rect 11256 6905 11284 6956
rect 11242 6896 11298 6905
rect 11242 6831 11298 6840
rect 11336 6860 11388 6866
rect 11336 6802 11388 6808
rect 11152 6792 11204 6798
rect 11152 6734 11204 6740
rect 11060 5024 11112 5030
rect 11060 4966 11112 4972
rect 11072 4554 11100 4966
rect 11060 4548 11112 4554
rect 11060 4490 11112 4496
rect 10968 3936 11020 3942
rect 10968 3878 11020 3884
rect 10784 3732 10836 3738
rect 10784 3674 10836 3680
rect 11072 3534 11100 4490
rect 11164 4298 11192 6734
rect 11244 6656 11296 6662
rect 11244 6598 11296 6604
rect 11256 6322 11284 6598
rect 11244 6316 11296 6322
rect 11244 6258 11296 6264
rect 11348 6118 11376 6802
rect 11440 6254 11468 7142
rect 11428 6248 11480 6254
rect 11428 6190 11480 6196
rect 11336 6112 11388 6118
rect 11336 6054 11388 6060
rect 11426 6080 11482 6089
rect 11426 6015 11482 6024
rect 11440 5710 11468 6015
rect 11428 5704 11480 5710
rect 11428 5646 11480 5652
rect 11336 5636 11388 5642
rect 11336 5578 11388 5584
rect 11244 5296 11296 5302
rect 11244 5238 11296 5244
rect 11256 4457 11284 5238
rect 11348 4758 11376 5578
rect 11440 5574 11468 5646
rect 11428 5568 11480 5574
rect 11428 5510 11480 5516
rect 11440 5234 11468 5510
rect 11428 5228 11480 5234
rect 11428 5170 11480 5176
rect 11532 4758 11560 7278
rect 11624 5794 11652 8570
rect 11716 8498 11744 9182
rect 11796 8832 11848 8838
rect 11796 8774 11848 8780
rect 11808 8634 11836 8774
rect 11796 8628 11848 8634
rect 11796 8570 11848 8576
rect 11704 8492 11756 8498
rect 11704 8434 11756 8440
rect 11900 8294 11928 9862
rect 12084 9722 12112 11194
rect 12360 9790 12388 11194
rect 12636 9926 12664 11194
rect 12952 11194 12954 11212
rect 13174 11194 13230 11250
rect 13450 11194 13506 11250
rect 13726 11194 13782 11250
rect 14002 11194 14058 11250
rect 14278 11194 14334 11250
rect 14554 11194 14610 11250
rect 14830 11194 14886 11250
rect 15106 11194 15162 11250
rect 15382 11194 15438 11250
rect 15658 11194 15714 11250
rect 15934 11194 15990 11250
rect 16210 11194 16266 11250
rect 16486 11194 16542 11250
rect 16762 11194 16818 11250
rect 17038 11194 17094 11250
rect 17314 11194 17370 11250
rect 17590 11194 17646 11250
rect 17866 11194 17922 11250
rect 18142 11194 18198 11250
rect 18418 11194 18474 11250
rect 18694 11194 18750 11250
rect 18970 11194 19026 11250
rect 19246 11194 19302 11250
rect 19522 11194 19578 11250
rect 19798 11194 19854 11250
rect 20074 11194 20130 11250
rect 20350 11194 20406 11250
rect 20626 11194 20682 11250
rect 20902 11194 20958 11250
rect 21178 11194 21234 11250
rect 21454 11194 21510 11250
rect 21730 11194 21786 11250
rect 22006 11194 22062 11250
rect 22282 11194 22338 11250
rect 22558 11194 22614 11250
rect 22834 11194 22890 11250
rect 23110 11194 23166 11250
rect 23386 11194 23442 11250
rect 23662 11194 23718 11250
rect 23938 11194 23994 11250
rect 24214 11194 24270 11250
rect 24490 11194 24546 11250
rect 24766 11194 24822 11250
rect 25042 11194 25098 11250
rect 25318 11194 25374 11250
rect 25594 11194 25650 11250
rect 25870 11194 25926 11250
rect 26146 11194 26202 11250
rect 26422 11194 26478 11250
rect 26698 11194 26754 11250
rect 26974 11194 27030 11250
rect 27250 11194 27306 11250
rect 27526 11194 27582 11250
rect 27802 11194 27858 11250
rect 28078 11194 28134 11250
rect 28354 11194 28410 11250
rect 28630 11194 28686 11250
rect 28906 11194 28962 11250
rect 29182 11194 29238 11250
rect 29458 11194 29514 11250
rect 29734 11194 29790 11250
rect 30010 11194 30066 11250
rect 30286 11194 30342 11250
rect 30562 11194 30618 11250
rect 30838 11194 30894 11250
rect 31114 11194 31170 11250
rect 31390 11194 31446 11250
rect 31666 11194 31722 11250
rect 31942 11194 31998 11250
rect 32218 11194 32274 11250
rect 32494 11194 32550 11250
rect 32770 11194 32826 11250
rect 33046 11194 33102 11250
rect 33322 11194 33378 11250
rect 33598 11194 33654 11250
rect 33874 11194 33930 11250
rect 34150 11194 34206 11250
rect 34426 11194 34482 11250
rect 34702 11194 34758 11250
rect 34978 11194 35034 11250
rect 35254 11194 35310 11250
rect 35530 11194 35586 11250
rect 35806 11194 35862 11250
rect 36082 11194 36138 11250
rect 36358 11194 36414 11250
rect 36634 11194 36690 11250
rect 36910 11194 36966 11250
rect 37186 11194 37242 11250
rect 37462 11194 37518 11250
rect 37738 11194 37794 11250
rect 12900 11154 12952 11160
rect 12992 10736 13044 10742
rect 12992 10678 13044 10684
rect 12900 10532 12952 10538
rect 12900 10474 12952 10480
rect 12808 10192 12860 10198
rect 12808 10134 12860 10140
rect 12624 9920 12676 9926
rect 12624 9862 12676 9868
rect 12348 9784 12400 9790
rect 12348 9726 12400 9732
rect 12072 9716 12124 9722
rect 12072 9658 12124 9664
rect 12072 9036 12124 9042
rect 12072 8978 12124 8984
rect 12084 8566 12112 8978
rect 12072 8560 12124 8566
rect 12072 8502 12124 8508
rect 12820 8498 12848 10134
rect 11980 8492 12032 8498
rect 11980 8434 12032 8440
rect 12716 8492 12768 8498
rect 12716 8434 12768 8440
rect 12808 8492 12860 8498
rect 12808 8434 12860 8440
rect 11992 8362 12020 8434
rect 11980 8356 12032 8362
rect 11980 8298 12032 8304
rect 11888 8288 11940 8294
rect 11888 8230 11940 8236
rect 12624 8288 12676 8294
rect 12624 8230 12676 8236
rect 12530 8120 12586 8129
rect 12348 8084 12400 8090
rect 12530 8055 12586 8064
rect 12348 8026 12400 8032
rect 11704 7404 11756 7410
rect 11704 7346 11756 7352
rect 11716 7002 11744 7346
rect 11888 7200 11940 7206
rect 11888 7142 11940 7148
rect 11980 7200 12032 7206
rect 11980 7142 12032 7148
rect 11704 6996 11756 7002
rect 11704 6938 11756 6944
rect 11900 6322 11928 7142
rect 11992 6866 12020 7142
rect 12360 7041 12388 8026
rect 12440 7880 12492 7886
rect 12440 7822 12492 7828
rect 12346 7032 12402 7041
rect 12452 7002 12480 7822
rect 12346 6967 12402 6976
rect 12440 6996 12492 7002
rect 12440 6938 12492 6944
rect 11980 6860 12032 6866
rect 11980 6802 12032 6808
rect 12348 6792 12400 6798
rect 12348 6734 12400 6740
rect 12164 6724 12216 6730
rect 12164 6666 12216 6672
rect 12176 6458 12204 6666
rect 12164 6452 12216 6458
rect 12164 6394 12216 6400
rect 11888 6316 11940 6322
rect 11888 6258 11940 6264
rect 11900 6202 11928 6258
rect 11808 6174 11928 6202
rect 11624 5766 11744 5794
rect 11612 5704 11664 5710
rect 11612 5646 11664 5652
rect 11336 4752 11388 4758
rect 11520 4752 11572 4758
rect 11336 4694 11388 4700
rect 11440 4712 11520 4740
rect 11242 4448 11298 4457
rect 11242 4383 11298 4392
rect 11164 4270 11284 4298
rect 11060 3528 11112 3534
rect 11060 3470 11112 3476
rect 10784 3392 10836 3398
rect 10784 3334 10836 3340
rect 10796 3194 10824 3334
rect 10784 3188 10836 3194
rect 10784 3130 10836 3136
rect 10796 2446 10824 3130
rect 11060 2848 11112 2854
rect 10874 2816 10930 2825
rect 10874 2751 10930 2760
rect 11058 2816 11060 2825
rect 11112 2816 11114 2825
rect 11058 2751 11114 2760
rect 10888 2666 10916 2751
rect 11150 2680 11206 2689
rect 10888 2650 11100 2666
rect 10888 2644 11112 2650
rect 10888 2638 11060 2644
rect 11150 2615 11206 2624
rect 11060 2586 11112 2592
rect 10968 2576 11020 2582
rect 10968 2518 11020 2524
rect 10784 2440 10836 2446
rect 10784 2382 10836 2388
rect 10506 2071 10562 2080
rect 10692 2100 10744 2106
rect 10692 2042 10744 2048
rect 10980 1290 11008 2518
rect 11060 2304 11112 2310
rect 11060 2246 11112 2252
rect 10968 1284 11020 1290
rect 10968 1226 11020 1232
rect 10232 1012 10284 1018
rect 10232 954 10284 960
rect 11072 56 11100 2246
rect 11164 1766 11192 2615
rect 11152 1760 11204 1766
rect 11152 1702 11204 1708
rect 11256 1698 11284 4270
rect 11348 4214 11376 4694
rect 11440 4457 11468 4712
rect 11520 4694 11572 4700
rect 11520 4616 11572 4622
rect 11520 4558 11572 4564
rect 11426 4448 11482 4457
rect 11426 4383 11482 4392
rect 11336 4208 11388 4214
rect 11336 4150 11388 4156
rect 11532 4146 11560 4558
rect 11428 4140 11480 4146
rect 11428 4082 11480 4088
rect 11520 4140 11572 4146
rect 11520 4082 11572 4088
rect 11440 3602 11468 4082
rect 11624 3738 11652 5646
rect 11716 4026 11744 5766
rect 11808 5234 11836 6174
rect 11980 6112 12032 6118
rect 11980 6054 12032 6060
rect 11992 5794 12020 6054
rect 11992 5766 12204 5794
rect 11992 5250 12020 5766
rect 12176 5642 12204 5766
rect 12256 5704 12308 5710
rect 12256 5646 12308 5652
rect 12072 5636 12124 5642
rect 12072 5578 12124 5584
rect 12164 5636 12216 5642
rect 12164 5578 12216 5584
rect 11900 5234 12020 5250
rect 11796 5228 11848 5234
rect 11796 5170 11848 5176
rect 11900 5228 12032 5234
rect 11900 5222 11980 5228
rect 11900 4826 11928 5222
rect 11980 5170 12032 5176
rect 11888 4820 11940 4826
rect 11888 4762 11940 4768
rect 11716 3998 11836 4026
rect 11704 3936 11756 3942
rect 11704 3878 11756 3884
rect 11612 3732 11664 3738
rect 11612 3674 11664 3680
rect 11428 3596 11480 3602
rect 11428 3538 11480 3544
rect 11716 3058 11744 3878
rect 11808 3194 11836 3998
rect 11900 3602 11928 4762
rect 11888 3596 11940 3602
rect 11888 3538 11940 3544
rect 12084 3448 12112 5578
rect 12164 5092 12216 5098
rect 12164 5034 12216 5040
rect 12176 4554 12204 5034
rect 12164 4548 12216 4554
rect 12164 4490 12216 4496
rect 12164 3460 12216 3466
rect 12084 3420 12164 3448
rect 12164 3402 12216 3408
rect 12268 3398 12296 5646
rect 12360 5574 12388 6734
rect 12348 5568 12400 5574
rect 12348 5510 12400 5516
rect 12452 4622 12480 6938
rect 12440 4616 12492 4622
rect 12440 4558 12492 4564
rect 12544 4486 12572 8055
rect 12636 7886 12664 8230
rect 12624 7880 12676 7886
rect 12624 7822 12676 7828
rect 12728 7721 12756 8434
rect 12714 7712 12770 7721
rect 12770 7670 12848 7698
rect 12714 7647 12770 7656
rect 12716 7404 12768 7410
rect 12716 7346 12768 7352
rect 12728 6474 12756 7346
rect 12820 6934 12848 7670
rect 12808 6928 12860 6934
rect 12808 6870 12860 6876
rect 12808 6792 12860 6798
rect 12808 6734 12860 6740
rect 12636 6446 12756 6474
rect 12636 5216 12664 6446
rect 12716 6384 12768 6390
rect 12716 6326 12768 6332
rect 12728 6118 12756 6326
rect 12716 6112 12768 6118
rect 12716 6054 12768 6060
rect 12636 5188 12756 5216
rect 12624 5092 12676 5098
rect 12624 5034 12676 5040
rect 12636 4865 12664 5034
rect 12622 4856 12678 4865
rect 12622 4791 12678 4800
rect 12624 4752 12676 4758
rect 12624 4694 12676 4700
rect 12532 4480 12584 4486
rect 12532 4422 12584 4428
rect 12636 4282 12664 4694
rect 12624 4276 12676 4282
rect 12624 4218 12676 4224
rect 12530 4176 12586 4185
rect 12530 4111 12586 4120
rect 12348 3460 12400 3466
rect 12348 3402 12400 3408
rect 11980 3392 12032 3398
rect 11980 3334 12032 3340
rect 12256 3392 12308 3398
rect 12256 3334 12308 3340
rect 11796 3188 11848 3194
rect 11796 3130 11848 3136
rect 11888 3188 11940 3194
rect 11888 3130 11940 3136
rect 11900 3074 11928 3130
rect 11808 3058 11928 3074
rect 11992 3058 12020 3334
rect 12254 3088 12310 3097
rect 11612 3052 11664 3058
rect 11612 2994 11664 3000
rect 11704 3052 11756 3058
rect 11704 2994 11756 3000
rect 11796 3052 11928 3058
rect 11848 3046 11928 3052
rect 11980 3052 12032 3058
rect 11796 2994 11848 3000
rect 12360 3074 12388 3402
rect 12310 3046 12388 3074
rect 12254 3023 12310 3032
rect 11980 2994 12032 3000
rect 11336 2848 11388 2854
rect 11336 2790 11388 2796
rect 11348 2514 11376 2790
rect 11624 2582 11652 2994
rect 12162 2680 12218 2689
rect 12162 2615 12218 2624
rect 11612 2576 11664 2582
rect 11612 2518 11664 2524
rect 11886 2544 11942 2553
rect 11336 2508 11388 2514
rect 11886 2479 11942 2488
rect 11336 2450 11388 2456
rect 11900 2446 11928 2479
rect 11888 2440 11940 2446
rect 11888 2382 11940 2388
rect 11980 2372 12032 2378
rect 11980 2314 12032 2320
rect 12072 2372 12124 2378
rect 12072 2314 12124 2320
rect 11704 2304 11756 2310
rect 11704 2246 11756 2252
rect 11716 2038 11744 2246
rect 11704 2032 11756 2038
rect 11704 1974 11756 1980
rect 11992 1970 12020 2314
rect 12084 2106 12112 2314
rect 12176 2106 12204 2615
rect 12348 2508 12400 2514
rect 12348 2450 12400 2456
rect 12360 2310 12388 2450
rect 12348 2304 12400 2310
rect 12348 2246 12400 2252
rect 12440 2304 12492 2310
rect 12440 2246 12492 2252
rect 12072 2100 12124 2106
rect 12072 2042 12124 2048
rect 12164 2100 12216 2106
rect 12164 2042 12216 2048
rect 11980 1964 12032 1970
rect 11980 1906 12032 1912
rect 11992 1698 12020 1906
rect 11244 1692 11296 1698
rect 11244 1634 11296 1640
rect 11980 1692 12032 1698
rect 11980 1634 12032 1640
rect 11150 1592 11206 1601
rect 11150 1527 11206 1536
rect 11164 1494 11192 1527
rect 11152 1488 11204 1494
rect 11152 1430 11204 1436
rect 12176 56 12296 82
rect 8772 54 8906 56
rect 8772 42 8800 54
rect 8588 14 8800 42
rect 8850 0 8906 54
rect 9954 0 10010 56
rect 11058 0 11114 56
rect 12162 54 12296 56
rect 12162 0 12218 54
rect 12268 42 12296 54
rect 12452 42 12480 2246
rect 12544 1698 12572 4111
rect 12728 3505 12756 5188
rect 12714 3496 12770 3505
rect 12714 3431 12770 3440
rect 12532 1692 12584 1698
rect 12532 1634 12584 1640
rect 12820 1562 12848 6734
rect 12912 6225 12940 10474
rect 13004 8634 13032 10678
rect 13188 9761 13216 11194
rect 13464 10305 13492 11194
rect 13450 10296 13506 10305
rect 13450 10231 13506 10240
rect 13740 9994 13768 11194
rect 13728 9988 13780 9994
rect 13728 9930 13780 9936
rect 14016 9858 14044 11194
rect 14004 9852 14056 9858
rect 14004 9794 14056 9800
rect 13174 9752 13230 9761
rect 13174 9687 13230 9696
rect 13084 9036 13136 9042
rect 13084 8978 13136 8984
rect 13096 8906 13124 8978
rect 13084 8900 13136 8906
rect 13084 8842 13136 8848
rect 13268 8900 13320 8906
rect 13268 8842 13320 8848
rect 12992 8628 13044 8634
rect 12992 8570 13044 8576
rect 12992 8424 13044 8430
rect 12992 8366 13044 8372
rect 13004 7478 13032 8366
rect 13176 7880 13228 7886
rect 13176 7822 13228 7828
rect 12992 7472 13044 7478
rect 12992 7414 13044 7420
rect 12898 6216 12954 6225
rect 12898 6151 12954 6160
rect 12900 5160 12952 5166
rect 12900 5102 12952 5108
rect 12912 4282 12940 5102
rect 13004 4808 13032 7414
rect 13188 7177 13216 7822
rect 13174 7168 13230 7177
rect 13174 7103 13230 7112
rect 13174 6624 13230 6633
rect 13174 6559 13230 6568
rect 13084 6112 13136 6118
rect 13084 6054 13136 6060
rect 13096 5778 13124 6054
rect 13084 5772 13136 5778
rect 13084 5714 13136 5720
rect 13084 4820 13136 4826
rect 13004 4780 13084 4808
rect 13084 4762 13136 4768
rect 12900 4276 12952 4282
rect 12900 4218 12952 4224
rect 13084 4140 13136 4146
rect 13084 4082 13136 4088
rect 13096 3534 13124 4082
rect 13188 3738 13216 6559
rect 13280 5409 13308 8842
rect 13728 8560 13780 8566
rect 13728 8502 13780 8508
rect 13544 8492 13596 8498
rect 13544 8434 13596 8440
rect 13556 8401 13584 8434
rect 13542 8392 13598 8401
rect 13542 8327 13598 8336
rect 13634 7984 13690 7993
rect 13452 7948 13504 7954
rect 13634 7919 13690 7928
rect 13452 7890 13504 7896
rect 13464 7392 13492 7890
rect 13544 7404 13596 7410
rect 13464 7364 13544 7392
rect 13360 7336 13412 7342
rect 13360 7278 13412 7284
rect 13372 7002 13400 7278
rect 13360 6996 13412 7002
rect 13360 6938 13412 6944
rect 13358 6216 13414 6225
rect 13358 6151 13414 6160
rect 13372 5681 13400 6151
rect 13358 5672 13414 5681
rect 13358 5607 13414 5616
rect 13266 5400 13322 5409
rect 13266 5335 13322 5344
rect 13360 5296 13412 5302
rect 13360 5238 13412 5244
rect 13372 4758 13400 5238
rect 13360 4752 13412 4758
rect 13360 4694 13412 4700
rect 13268 4684 13320 4690
rect 13268 4626 13320 4632
rect 13280 4146 13308 4626
rect 13360 4548 13412 4554
rect 13360 4490 13412 4496
rect 13372 4282 13400 4490
rect 13464 4282 13492 7364
rect 13544 7346 13596 7352
rect 13648 6934 13676 7919
rect 13740 7886 13768 8502
rect 14096 8424 14148 8430
rect 13832 8372 14096 8378
rect 13832 8366 14148 8372
rect 13832 8350 14136 8366
rect 13728 7880 13780 7886
rect 13728 7822 13780 7828
rect 13728 7744 13780 7750
rect 13726 7712 13728 7721
rect 13780 7712 13782 7721
rect 13726 7647 13782 7656
rect 13832 7206 13860 8350
rect 13950 8188 14258 8197
rect 13950 8186 13956 8188
rect 14012 8186 14036 8188
rect 14092 8186 14116 8188
rect 14172 8186 14196 8188
rect 14252 8186 14258 8188
rect 14012 8134 14014 8186
rect 14194 8134 14196 8186
rect 13950 8132 13956 8134
rect 14012 8132 14036 8134
rect 14092 8132 14116 8134
rect 14172 8132 14196 8134
rect 14252 8132 14258 8134
rect 13950 8123 14258 8132
rect 13912 7812 13964 7818
rect 14188 7812 14240 7818
rect 13964 7772 14188 7800
rect 13912 7754 13964 7760
rect 14188 7754 14240 7760
rect 14292 7206 14320 11194
rect 14568 10742 14596 11194
rect 14556 10736 14608 10742
rect 14556 10678 14608 10684
rect 14844 10010 14872 11194
rect 14752 9982 14872 10010
rect 14752 8838 14780 9982
rect 14830 9752 14886 9761
rect 14830 9687 14886 9696
rect 14740 8832 14792 8838
rect 14740 8774 14792 8780
rect 14370 8664 14426 8673
rect 14370 8599 14426 8608
rect 14738 8664 14794 8673
rect 14738 8599 14794 8608
rect 13820 7200 13872 7206
rect 13820 7142 13872 7148
rect 14280 7200 14332 7206
rect 14280 7142 14332 7148
rect 13636 6928 13688 6934
rect 13634 6896 13636 6905
rect 13688 6896 13690 6905
rect 13634 6831 13690 6840
rect 13636 6724 13688 6730
rect 13636 6666 13688 6672
rect 13544 6656 13596 6662
rect 13544 6598 13596 6604
rect 13556 6390 13584 6598
rect 13544 6384 13596 6390
rect 13544 6326 13596 6332
rect 13544 6112 13596 6118
rect 13544 6054 13596 6060
rect 13360 4276 13412 4282
rect 13360 4218 13412 4224
rect 13452 4276 13504 4282
rect 13452 4218 13504 4224
rect 13556 4146 13584 6054
rect 13648 5710 13676 6666
rect 13832 6390 13860 7142
rect 13950 7100 14258 7109
rect 13950 7098 13956 7100
rect 14012 7098 14036 7100
rect 14092 7098 14116 7100
rect 14172 7098 14196 7100
rect 14252 7098 14258 7100
rect 14012 7046 14014 7098
rect 14194 7046 14196 7098
rect 13950 7044 13956 7046
rect 14012 7044 14036 7046
rect 14092 7044 14116 7046
rect 14172 7044 14196 7046
rect 14252 7044 14258 7046
rect 13950 7035 14258 7044
rect 13912 6792 13964 6798
rect 13912 6734 13964 6740
rect 13924 6390 13952 6734
rect 14188 6656 14240 6662
rect 14188 6598 14240 6604
rect 14280 6656 14332 6662
rect 14280 6598 14332 6604
rect 13820 6384 13872 6390
rect 13820 6326 13872 6332
rect 13912 6384 13964 6390
rect 13912 6326 13964 6332
rect 14200 6254 14228 6598
rect 14188 6248 14240 6254
rect 14188 6190 14240 6196
rect 13820 6180 13872 6186
rect 13820 6122 13872 6128
rect 13832 5914 13860 6122
rect 13950 6012 14258 6021
rect 13950 6010 13956 6012
rect 14012 6010 14036 6012
rect 14092 6010 14116 6012
rect 14172 6010 14196 6012
rect 14252 6010 14258 6012
rect 14012 5958 14014 6010
rect 14194 5958 14196 6010
rect 13950 5956 13956 5958
rect 14012 5956 14036 5958
rect 14092 5956 14116 5958
rect 14172 5956 14196 5958
rect 14252 5956 14258 5958
rect 13950 5947 14258 5956
rect 14292 5914 14320 6598
rect 13820 5908 13872 5914
rect 13820 5850 13872 5856
rect 14280 5908 14332 5914
rect 14280 5850 14332 5856
rect 13636 5704 13688 5710
rect 13636 5646 13688 5652
rect 14188 5160 14240 5166
rect 14188 5102 14240 5108
rect 14200 5030 14228 5102
rect 14188 5024 14240 5030
rect 14188 4966 14240 4972
rect 13950 4924 14258 4933
rect 13950 4922 13956 4924
rect 14012 4922 14036 4924
rect 14092 4922 14116 4924
rect 14172 4922 14196 4924
rect 14252 4922 14258 4924
rect 14012 4870 14014 4922
rect 14194 4870 14196 4922
rect 13950 4868 13956 4870
rect 14012 4868 14036 4870
rect 14092 4868 14116 4870
rect 14172 4868 14196 4870
rect 14252 4868 14258 4870
rect 13950 4859 14258 4868
rect 14292 4740 14320 5850
rect 14108 4712 14320 4740
rect 14108 4146 14136 4712
rect 14384 4622 14412 8599
rect 14752 8566 14780 8599
rect 14648 8560 14700 8566
rect 14648 8502 14700 8508
rect 14740 8560 14792 8566
rect 14740 8502 14792 8508
rect 14464 8288 14516 8294
rect 14464 8230 14516 8236
rect 14476 7886 14504 8230
rect 14660 8022 14688 8502
rect 14844 8498 14872 9687
rect 15120 8820 15148 11194
rect 15198 9072 15254 9081
rect 15198 9007 15254 9016
rect 15212 8906 15240 9007
rect 15200 8900 15252 8906
rect 15200 8842 15252 8848
rect 14936 8792 15148 8820
rect 14936 8634 14964 8792
rect 15010 8732 15318 8741
rect 15010 8730 15016 8732
rect 15072 8730 15096 8732
rect 15152 8730 15176 8732
rect 15232 8730 15256 8732
rect 15312 8730 15318 8732
rect 15072 8678 15074 8730
rect 15254 8678 15256 8730
rect 15010 8676 15016 8678
rect 15072 8676 15096 8678
rect 15152 8676 15176 8678
rect 15232 8676 15256 8678
rect 15312 8676 15318 8678
rect 15010 8667 15318 8676
rect 14924 8628 14976 8634
rect 14924 8570 14976 8576
rect 14832 8492 14884 8498
rect 14832 8434 14884 8440
rect 15292 8492 15344 8498
rect 15396 8480 15424 11194
rect 15566 9344 15622 9353
rect 15566 9279 15622 9288
rect 15580 8498 15608 9279
rect 15344 8452 15424 8480
rect 15568 8492 15620 8498
rect 15292 8434 15344 8440
rect 15568 8434 15620 8440
rect 15672 8362 15700 11194
rect 15750 9480 15806 9489
rect 15750 9415 15806 9424
rect 15764 8498 15792 9415
rect 15948 8566 15976 11194
rect 16118 10296 16174 10305
rect 16118 10231 16174 10240
rect 16028 8832 16080 8838
rect 16028 8774 16080 8780
rect 15936 8560 15988 8566
rect 15936 8502 15988 8508
rect 15752 8492 15804 8498
rect 15752 8434 15804 8440
rect 16040 8362 16068 8774
rect 15660 8356 15712 8362
rect 15660 8298 15712 8304
rect 16028 8356 16080 8362
rect 16028 8298 16080 8304
rect 14832 8288 14884 8294
rect 14738 8256 14794 8265
rect 14832 8230 14884 8236
rect 14924 8288 14976 8294
rect 14924 8230 14976 8236
rect 14738 8191 14794 8200
rect 14648 8016 14700 8022
rect 14554 7984 14610 7993
rect 14648 7958 14700 7964
rect 14554 7919 14610 7928
rect 14464 7880 14516 7886
rect 14464 7822 14516 7828
rect 14476 6322 14504 7822
rect 14568 7449 14596 7919
rect 14648 7880 14700 7886
rect 14648 7822 14700 7828
rect 14660 7478 14688 7822
rect 14648 7472 14700 7478
rect 14554 7440 14610 7449
rect 14648 7414 14700 7420
rect 14554 7375 14610 7384
rect 14556 7200 14608 7206
rect 14556 7142 14608 7148
rect 14568 6866 14596 7142
rect 14556 6860 14608 6866
rect 14556 6802 14608 6808
rect 14464 6316 14516 6322
rect 14464 6258 14516 6264
rect 14556 6112 14608 6118
rect 14462 6080 14518 6089
rect 14556 6054 14608 6060
rect 14462 6015 14518 6024
rect 14476 5846 14504 6015
rect 14464 5840 14516 5846
rect 14464 5782 14516 5788
rect 14568 5681 14596 6054
rect 14554 5672 14610 5681
rect 14554 5607 14610 5616
rect 14464 5024 14516 5030
rect 14464 4966 14516 4972
rect 14476 4758 14504 4966
rect 14464 4752 14516 4758
rect 14464 4694 14516 4700
rect 14188 4616 14240 4622
rect 14372 4616 14424 4622
rect 14240 4576 14320 4604
rect 14188 4558 14240 4564
rect 13268 4140 13320 4146
rect 13268 4082 13320 4088
rect 13544 4140 13596 4146
rect 13544 4082 13596 4088
rect 14096 4140 14148 4146
rect 14096 4082 14148 4088
rect 13820 4072 13872 4078
rect 13820 4014 13872 4020
rect 13176 3732 13228 3738
rect 13176 3674 13228 3680
rect 13728 3732 13780 3738
rect 13728 3674 13780 3680
rect 13268 3664 13320 3670
rect 13268 3606 13320 3612
rect 13084 3528 13136 3534
rect 13084 3470 13136 3476
rect 13174 3224 13230 3233
rect 13174 3159 13230 3168
rect 12898 3088 12954 3097
rect 13188 3058 13216 3159
rect 12898 3023 12900 3032
rect 12952 3023 12954 3032
rect 13176 3052 13228 3058
rect 12900 2994 12952 3000
rect 13176 2994 13228 3000
rect 13188 2514 13216 2994
rect 13176 2508 13228 2514
rect 13176 2450 13228 2456
rect 13084 2304 13136 2310
rect 13084 2246 13136 2252
rect 12808 1556 12860 1562
rect 12808 1498 12860 1504
rect 13096 1222 13124 2246
rect 13084 1216 13136 1222
rect 13084 1158 13136 1164
rect 13280 56 13308 3606
rect 13740 3602 13768 3674
rect 13728 3596 13780 3602
rect 13728 3538 13780 3544
rect 13452 3528 13504 3534
rect 13452 3470 13504 3476
rect 13634 3496 13690 3505
rect 13464 2650 13492 3470
rect 13634 3431 13690 3440
rect 13648 3398 13676 3431
rect 13636 3392 13688 3398
rect 13636 3334 13688 3340
rect 13832 3194 13860 4014
rect 13950 3836 14258 3845
rect 13950 3834 13956 3836
rect 14012 3834 14036 3836
rect 14092 3834 14116 3836
rect 14172 3834 14196 3836
rect 14252 3834 14258 3836
rect 14012 3782 14014 3834
rect 14194 3782 14196 3834
rect 13950 3780 13956 3782
rect 14012 3780 14036 3782
rect 14092 3780 14116 3782
rect 14172 3780 14196 3782
rect 14252 3780 14258 3782
rect 13950 3771 14258 3780
rect 14292 3534 14320 4576
rect 14372 4558 14424 4564
rect 14476 4214 14504 4694
rect 14372 4208 14424 4214
rect 14372 4150 14424 4156
rect 14464 4208 14516 4214
rect 14464 4150 14516 4156
rect 14280 3528 14332 3534
rect 14002 3496 14058 3505
rect 14280 3470 14332 3476
rect 14002 3431 14058 3440
rect 14096 3460 14148 3466
rect 14016 3398 14044 3431
rect 14096 3402 14148 3408
rect 14004 3392 14056 3398
rect 14004 3334 14056 3340
rect 13636 3188 13688 3194
rect 13636 3130 13688 3136
rect 13820 3188 13872 3194
rect 14004 3188 14056 3194
rect 13820 3130 13872 3136
rect 13924 3148 14004 3176
rect 13544 2984 13596 2990
rect 13544 2926 13596 2932
rect 13556 2825 13584 2926
rect 13648 2922 13676 3130
rect 13924 3074 13952 3148
rect 14004 3130 14056 3136
rect 13832 3046 13952 3074
rect 14002 3088 14058 3097
rect 13636 2916 13688 2922
rect 13636 2858 13688 2864
rect 13728 2848 13780 2854
rect 13542 2816 13598 2825
rect 13728 2790 13780 2796
rect 13542 2751 13598 2760
rect 13452 2644 13504 2650
rect 13452 2586 13504 2592
rect 13740 2514 13768 2790
rect 13728 2508 13780 2514
rect 13728 2450 13780 2456
rect 13832 1902 13860 3046
rect 14002 3023 14058 3032
rect 14016 2990 14044 3023
rect 13912 2984 13964 2990
rect 13912 2926 13964 2932
rect 14004 2984 14056 2990
rect 14004 2926 14056 2932
rect 13924 2836 13952 2926
rect 14108 2836 14136 3402
rect 13924 2808 14136 2836
rect 14384 2825 14412 4150
rect 14464 3732 14516 3738
rect 14464 3674 14516 3680
rect 14476 3602 14504 3674
rect 14464 3596 14516 3602
rect 14464 3538 14516 3544
rect 14568 3194 14596 5607
rect 14752 5352 14780 8191
rect 14844 8129 14872 8230
rect 14830 8120 14886 8129
rect 14830 8055 14886 8064
rect 14830 7712 14886 7721
rect 14830 7647 14886 7656
rect 14844 5953 14872 7647
rect 14936 6186 14964 8230
rect 15658 8120 15714 8129
rect 15658 8055 15714 8064
rect 15108 7880 15160 7886
rect 15160 7840 15424 7868
rect 15108 7822 15160 7828
rect 15010 7644 15318 7653
rect 15010 7642 15016 7644
rect 15072 7642 15096 7644
rect 15152 7642 15176 7644
rect 15232 7642 15256 7644
rect 15312 7642 15318 7644
rect 15072 7590 15074 7642
rect 15254 7590 15256 7642
rect 15010 7588 15016 7590
rect 15072 7588 15096 7590
rect 15152 7588 15176 7590
rect 15232 7588 15256 7590
rect 15312 7588 15318 7590
rect 15010 7579 15318 7588
rect 15396 7528 15424 7840
rect 15476 7744 15528 7750
rect 15476 7686 15528 7692
rect 15304 7500 15424 7528
rect 15304 7410 15332 7500
rect 15292 7404 15344 7410
rect 15292 7346 15344 7352
rect 15384 7404 15436 7410
rect 15384 7346 15436 7352
rect 15488 7392 15516 7686
rect 15568 7404 15620 7410
rect 15488 7364 15568 7392
rect 15010 6556 15318 6565
rect 15010 6554 15016 6556
rect 15072 6554 15096 6556
rect 15152 6554 15176 6556
rect 15232 6554 15256 6556
rect 15312 6554 15318 6556
rect 15072 6502 15074 6554
rect 15254 6502 15256 6554
rect 15010 6500 15016 6502
rect 15072 6500 15096 6502
rect 15152 6500 15176 6502
rect 15232 6500 15256 6502
rect 15312 6500 15318 6502
rect 15010 6491 15318 6500
rect 15108 6316 15160 6322
rect 15108 6258 15160 6264
rect 14924 6180 14976 6186
rect 14924 6122 14976 6128
rect 14830 5944 14886 5953
rect 14830 5879 14886 5888
rect 14660 5324 14780 5352
rect 14660 4282 14688 5324
rect 14740 5228 14792 5234
rect 14740 5170 14792 5176
rect 14752 4690 14780 5170
rect 14832 5160 14884 5166
rect 14832 5102 14884 5108
rect 14844 5001 14872 5102
rect 14830 4992 14886 5001
rect 14830 4927 14886 4936
rect 14936 4826 14964 6122
rect 15120 5914 15148 6258
rect 15108 5908 15160 5914
rect 15108 5850 15160 5856
rect 15120 5642 15148 5850
rect 15108 5636 15160 5642
rect 15108 5578 15160 5584
rect 15010 5468 15318 5477
rect 15010 5466 15016 5468
rect 15072 5466 15096 5468
rect 15152 5466 15176 5468
rect 15232 5466 15256 5468
rect 15312 5466 15318 5468
rect 15072 5414 15074 5466
rect 15254 5414 15256 5466
rect 15010 5412 15016 5414
rect 15072 5412 15096 5414
rect 15152 5412 15176 5414
rect 15232 5412 15256 5414
rect 15312 5412 15318 5414
rect 15010 5403 15318 5412
rect 14924 4820 14976 4826
rect 14924 4762 14976 4768
rect 14740 4684 14792 4690
rect 14740 4626 14792 4632
rect 15396 4486 15424 7346
rect 15488 6730 15516 7364
rect 15568 7346 15620 7352
rect 15672 7188 15700 8055
rect 15752 7880 15804 7886
rect 15752 7822 15804 7828
rect 15764 7256 15792 7822
rect 15844 7812 15896 7818
rect 15844 7754 15896 7760
rect 15856 7410 15884 7754
rect 16026 7712 16082 7721
rect 16026 7647 16082 7656
rect 15936 7540 15988 7546
rect 15936 7482 15988 7488
rect 15948 7449 15976 7482
rect 15934 7440 15990 7449
rect 15844 7404 15896 7410
rect 16040 7410 16068 7647
rect 15934 7375 15990 7384
rect 16028 7404 16080 7410
rect 15844 7346 15896 7352
rect 16028 7346 16080 7352
rect 15936 7268 15988 7274
rect 15764 7228 15884 7256
rect 15672 7160 15792 7188
rect 15660 6860 15712 6866
rect 15660 6802 15712 6808
rect 15476 6724 15528 6730
rect 15476 6666 15528 6672
rect 15488 6390 15516 6666
rect 15672 6662 15700 6802
rect 15660 6656 15712 6662
rect 15660 6598 15712 6604
rect 15476 6384 15528 6390
rect 15476 6326 15528 6332
rect 15568 6316 15620 6322
rect 15568 6258 15620 6264
rect 15580 5914 15608 6258
rect 15568 5908 15620 5914
rect 15568 5850 15620 5856
rect 15476 5704 15528 5710
rect 15660 5704 15712 5710
rect 15476 5646 15528 5652
rect 15658 5672 15660 5681
rect 15712 5672 15714 5681
rect 15488 5302 15516 5646
rect 15658 5607 15714 5616
rect 15764 5545 15792 7160
rect 15750 5536 15806 5545
rect 15750 5471 15806 5480
rect 15476 5296 15528 5302
rect 15476 5238 15528 5244
rect 15660 5296 15712 5302
rect 15660 5238 15712 5244
rect 15476 4820 15528 4826
rect 15476 4762 15528 4768
rect 14832 4480 14884 4486
rect 14738 4448 14794 4457
rect 14832 4422 14884 4428
rect 15384 4480 15436 4486
rect 15384 4422 15436 4428
rect 14738 4383 14794 4392
rect 14648 4276 14700 4282
rect 14648 4218 14700 4224
rect 14752 4060 14780 4383
rect 14844 4214 14872 4422
rect 15010 4380 15318 4389
rect 15010 4378 15016 4380
rect 15072 4378 15096 4380
rect 15152 4378 15176 4380
rect 15232 4378 15256 4380
rect 15312 4378 15318 4380
rect 15072 4326 15074 4378
rect 15254 4326 15256 4378
rect 15010 4324 15016 4326
rect 15072 4324 15096 4326
rect 15152 4324 15176 4326
rect 15232 4324 15256 4326
rect 15312 4324 15318 4326
rect 15010 4315 15318 4324
rect 15384 4276 15436 4282
rect 15384 4218 15436 4224
rect 14832 4208 14884 4214
rect 15396 4185 15424 4218
rect 14832 4150 14884 4156
rect 15382 4176 15438 4185
rect 15382 4111 15438 4120
rect 14832 4072 14884 4078
rect 14752 4032 14832 4060
rect 14832 4014 14884 4020
rect 14830 3904 14886 3913
rect 14830 3839 14886 3848
rect 14740 3732 14792 3738
rect 14740 3674 14792 3680
rect 14752 3534 14780 3674
rect 14844 3534 14872 3839
rect 15384 3596 15436 3602
rect 15384 3538 15436 3544
rect 14740 3528 14792 3534
rect 14740 3470 14792 3476
rect 14832 3528 14884 3534
rect 15108 3528 15160 3534
rect 14832 3470 14884 3476
rect 14936 3476 15108 3482
rect 14936 3470 15160 3476
rect 14936 3454 15148 3470
rect 14830 3224 14886 3233
rect 14556 3188 14608 3194
rect 14830 3159 14886 3168
rect 14556 3130 14608 3136
rect 14648 3120 14700 3126
rect 14568 3068 14648 3074
rect 14568 3062 14700 3068
rect 14568 3046 14688 3062
rect 14844 3058 14872 3159
rect 14832 3052 14884 3058
rect 14370 2816 14426 2825
rect 13950 2748 14258 2757
rect 14370 2751 14426 2760
rect 13950 2746 13956 2748
rect 14012 2746 14036 2748
rect 14092 2746 14116 2748
rect 14172 2746 14196 2748
rect 14252 2746 14258 2748
rect 14012 2694 14014 2746
rect 14194 2694 14196 2746
rect 13950 2692 13956 2694
rect 14012 2692 14036 2694
rect 14092 2692 14116 2694
rect 14172 2692 14196 2694
rect 14252 2692 14258 2694
rect 13950 2683 14258 2692
rect 14384 2394 14412 2751
rect 14568 2650 14596 3046
rect 14832 2994 14884 3000
rect 14936 2990 14964 3454
rect 15396 3398 15424 3538
rect 15488 3398 15516 4762
rect 15672 4672 15700 5238
rect 15764 5001 15792 5471
rect 15750 4992 15806 5001
rect 15750 4927 15806 4936
rect 15752 4684 15804 4690
rect 15672 4644 15752 4672
rect 15568 4480 15620 4486
rect 15568 4422 15620 4428
rect 15384 3392 15436 3398
rect 15384 3334 15436 3340
rect 15476 3392 15528 3398
rect 15476 3334 15528 3340
rect 15010 3292 15318 3301
rect 15010 3290 15016 3292
rect 15072 3290 15096 3292
rect 15152 3290 15176 3292
rect 15232 3290 15256 3292
rect 15312 3290 15318 3292
rect 15072 3238 15074 3290
rect 15254 3238 15256 3290
rect 15010 3236 15016 3238
rect 15072 3236 15096 3238
rect 15152 3236 15176 3238
rect 15232 3236 15256 3238
rect 15312 3236 15318 3238
rect 15010 3227 15318 3236
rect 14924 2984 14976 2990
rect 14924 2926 14976 2932
rect 14740 2848 14792 2854
rect 14740 2790 14792 2796
rect 15016 2848 15068 2854
rect 15016 2790 15068 2796
rect 14556 2644 14608 2650
rect 14556 2586 14608 2592
rect 14648 2644 14700 2650
rect 14648 2586 14700 2592
rect 14554 2544 14610 2553
rect 14554 2479 14610 2488
rect 14568 2446 14596 2479
rect 14292 2366 14412 2394
rect 14556 2440 14608 2446
rect 14556 2382 14608 2388
rect 14292 2281 14320 2366
rect 14372 2304 14424 2310
rect 14278 2272 14334 2281
rect 14372 2246 14424 2252
rect 14278 2207 14334 2216
rect 13820 1896 13872 1902
rect 13820 1838 13872 1844
rect 14384 56 14412 2246
rect 14660 2145 14688 2586
rect 14752 2446 14780 2790
rect 15028 2514 15056 2790
rect 15488 2650 15516 3334
rect 15476 2644 15528 2650
rect 15476 2586 15528 2592
rect 15580 2514 15608 4422
rect 15672 4185 15700 4644
rect 15752 4626 15804 4632
rect 15752 4276 15804 4282
rect 15752 4218 15804 4224
rect 15658 4176 15714 4185
rect 15658 4111 15714 4120
rect 15658 3768 15714 3777
rect 15658 3703 15714 3712
rect 15672 3398 15700 3703
rect 15660 3392 15712 3398
rect 15660 3334 15712 3340
rect 15016 2508 15068 2514
rect 15016 2450 15068 2456
rect 15568 2508 15620 2514
rect 15568 2450 15620 2456
rect 14740 2440 14792 2446
rect 14740 2382 14792 2388
rect 15476 2304 15528 2310
rect 15476 2246 15528 2252
rect 15010 2204 15318 2213
rect 15010 2202 15016 2204
rect 15072 2202 15096 2204
rect 15152 2202 15176 2204
rect 15232 2202 15256 2204
rect 15312 2202 15318 2204
rect 15072 2150 15074 2202
rect 15254 2150 15256 2202
rect 15010 2148 15016 2150
rect 15072 2148 15096 2150
rect 15152 2148 15176 2150
rect 15232 2148 15256 2150
rect 15312 2148 15318 2150
rect 14646 2136 14702 2145
rect 15010 2139 15318 2148
rect 14646 2071 14702 2080
rect 15488 56 15516 2246
rect 15764 2038 15792 4218
rect 15856 3618 15884 7228
rect 15936 7210 15988 7216
rect 15948 7041 15976 7210
rect 16028 7200 16080 7206
rect 16026 7168 16028 7177
rect 16080 7168 16082 7177
rect 16026 7103 16082 7112
rect 15934 7032 15990 7041
rect 15934 6967 15990 6976
rect 15948 5914 15976 6967
rect 16028 6656 16080 6662
rect 16028 6598 16080 6604
rect 16040 6497 16068 6598
rect 16026 6488 16082 6497
rect 16026 6423 16082 6432
rect 15936 5908 15988 5914
rect 15936 5850 15988 5856
rect 16028 5704 16080 5710
rect 15948 5664 16028 5692
rect 15948 5556 15976 5664
rect 16028 5646 16080 5652
rect 15948 5528 16068 5556
rect 16040 4264 16068 5528
rect 16132 5352 16160 10231
rect 16224 8634 16252 11194
rect 16304 9308 16356 9314
rect 16304 9250 16356 9256
rect 16212 8628 16264 8634
rect 16212 8570 16264 8576
rect 16316 8129 16344 9250
rect 16500 8838 16528 11194
rect 16488 8832 16540 8838
rect 16488 8774 16540 8780
rect 16776 8634 16804 11194
rect 16948 9852 17000 9858
rect 16948 9794 17000 9800
rect 16856 9308 16908 9314
rect 16856 9250 16908 9256
rect 16868 9110 16896 9250
rect 16856 9104 16908 9110
rect 16856 9046 16908 9052
rect 16764 8628 16816 8634
rect 16764 8570 16816 8576
rect 16856 8560 16908 8566
rect 16856 8502 16908 8508
rect 16396 8424 16448 8430
rect 16396 8366 16448 8372
rect 16672 8424 16724 8430
rect 16672 8366 16724 8372
rect 16302 8120 16358 8129
rect 16302 8055 16358 8064
rect 16212 7472 16264 7478
rect 16212 7414 16264 7420
rect 16224 6338 16252 7414
rect 16408 6390 16436 8366
rect 16684 8090 16712 8366
rect 16580 8084 16632 8090
rect 16580 8026 16632 8032
rect 16672 8084 16724 8090
rect 16672 8026 16724 8032
rect 16592 7750 16620 8026
rect 16580 7744 16632 7750
rect 16684 7721 16712 8026
rect 16580 7686 16632 7692
rect 16670 7712 16726 7721
rect 16670 7647 16726 7656
rect 16580 7540 16632 7546
rect 16580 7482 16632 7488
rect 16396 6384 16448 6390
rect 16224 6310 16344 6338
rect 16396 6326 16448 6332
rect 16486 6352 16542 6361
rect 16316 6118 16344 6310
rect 16592 6322 16620 7482
rect 16672 7472 16724 7478
rect 16672 7414 16724 7420
rect 16684 7206 16712 7414
rect 16868 7206 16896 8502
rect 16672 7200 16724 7206
rect 16672 7142 16724 7148
rect 16856 7200 16908 7206
rect 16856 7142 16908 7148
rect 16670 6896 16726 6905
rect 16670 6831 16726 6840
rect 16684 6798 16712 6831
rect 16672 6792 16724 6798
rect 16672 6734 16724 6740
rect 16764 6656 16816 6662
rect 16670 6624 16726 6633
rect 16764 6598 16816 6604
rect 16670 6559 16726 6568
rect 16486 6287 16542 6296
rect 16580 6316 16632 6322
rect 16396 6248 16448 6254
rect 16396 6190 16448 6196
rect 16304 6112 16356 6118
rect 16304 6054 16356 6060
rect 16212 5840 16264 5846
rect 16212 5782 16264 5788
rect 16304 5840 16356 5846
rect 16408 5828 16436 6190
rect 16356 5800 16436 5828
rect 16304 5782 16356 5788
rect 16224 5710 16252 5782
rect 16212 5704 16264 5710
rect 16500 5692 16528 6287
rect 16580 6258 16632 6264
rect 16580 5704 16632 5710
rect 16264 5664 16344 5692
rect 16212 5646 16264 5652
rect 16212 5364 16264 5370
rect 16132 5324 16212 5352
rect 16212 5306 16264 5312
rect 16212 5024 16264 5030
rect 16212 4966 16264 4972
rect 16040 4236 16160 4264
rect 16026 4176 16082 4185
rect 16026 4111 16028 4120
rect 16080 4111 16082 4120
rect 16028 4082 16080 4088
rect 16132 4078 16160 4236
rect 16120 4072 16172 4078
rect 16120 4014 16172 4020
rect 16028 4004 16080 4010
rect 16028 3946 16080 3952
rect 16040 3670 16068 3946
rect 16028 3664 16080 3670
rect 15856 3590 15976 3618
rect 16028 3606 16080 3612
rect 15844 3528 15896 3534
rect 15844 3470 15896 3476
rect 15856 2650 15884 3470
rect 15844 2644 15896 2650
rect 15844 2586 15896 2592
rect 15948 2446 15976 3590
rect 16224 3505 16252 4966
rect 16316 4604 16344 5664
rect 16500 5664 16580 5692
rect 16396 4616 16448 4622
rect 16316 4576 16396 4604
rect 16396 4558 16448 4564
rect 16304 4480 16356 4486
rect 16304 4422 16356 4428
rect 16396 4480 16448 4486
rect 16396 4422 16448 4428
rect 16210 3496 16266 3505
rect 16210 3431 16266 3440
rect 16118 3360 16174 3369
rect 16118 3295 16174 3304
rect 16028 3188 16080 3194
rect 16028 3130 16080 3136
rect 15844 2440 15896 2446
rect 15844 2382 15896 2388
rect 15936 2440 15988 2446
rect 15936 2382 15988 2388
rect 15856 2292 15884 2382
rect 16040 2292 16068 3130
rect 16132 3126 16160 3295
rect 16120 3120 16172 3126
rect 16120 3062 16172 3068
rect 15856 2264 16068 2292
rect 15752 2032 15804 2038
rect 15752 1974 15804 1980
rect 16316 1834 16344 4422
rect 16408 4282 16436 4422
rect 16396 4276 16448 4282
rect 16396 4218 16448 4224
rect 16500 4146 16528 5664
rect 16580 5646 16632 5652
rect 16684 5642 16712 6559
rect 16672 5636 16724 5642
rect 16672 5578 16724 5584
rect 16684 4826 16712 5578
rect 16672 4820 16724 4826
rect 16672 4762 16724 4768
rect 16672 4616 16724 4622
rect 16672 4558 16724 4564
rect 16684 4282 16712 4558
rect 16672 4276 16724 4282
rect 16672 4218 16724 4224
rect 16776 4214 16804 6598
rect 16960 6322 16988 9794
rect 17052 8634 17080 11194
rect 17224 10872 17276 10878
rect 17224 10814 17276 10820
rect 17132 10328 17184 10334
rect 17132 10270 17184 10276
rect 17144 9722 17172 10270
rect 17132 9716 17184 9722
rect 17132 9658 17184 9664
rect 17132 9512 17184 9518
rect 17132 9454 17184 9460
rect 17040 8628 17092 8634
rect 17040 8570 17092 8576
rect 17038 8528 17094 8537
rect 17038 8463 17094 8472
rect 17052 8022 17080 8463
rect 17040 8016 17092 8022
rect 17040 7958 17092 7964
rect 17040 7472 17092 7478
rect 17040 7414 17092 7420
rect 16856 6316 16908 6322
rect 16856 6258 16908 6264
rect 16948 6316 17000 6322
rect 16948 6258 17000 6264
rect 16868 5273 16896 6258
rect 17052 6254 17080 7414
rect 17144 6662 17172 9454
rect 17236 6798 17264 10814
rect 17328 8090 17356 11194
rect 17406 10296 17462 10305
rect 17406 10231 17462 10240
rect 17500 10260 17552 10266
rect 17420 9897 17448 10231
rect 17500 10202 17552 10208
rect 17512 10062 17540 10202
rect 17500 10056 17552 10062
rect 17500 9998 17552 10004
rect 17406 9888 17462 9897
rect 17406 9823 17462 9832
rect 17500 9512 17552 9518
rect 17500 9454 17552 9460
rect 17512 8498 17540 9454
rect 17500 8492 17552 8498
rect 17500 8434 17552 8440
rect 17408 8424 17460 8430
rect 17408 8366 17460 8372
rect 17316 8084 17368 8090
rect 17316 8026 17368 8032
rect 17420 7886 17448 8366
rect 17408 7880 17460 7886
rect 17408 7822 17460 7828
rect 17406 6896 17462 6905
rect 17316 6860 17368 6866
rect 17604 6866 17632 11194
rect 17682 10568 17738 10577
rect 17682 10503 17738 10512
rect 17696 9897 17724 10503
rect 17682 9888 17738 9897
rect 17682 9823 17738 9832
rect 17880 8514 17908 11194
rect 17960 9444 18012 9450
rect 17960 9386 18012 9392
rect 17972 8945 18000 9386
rect 18052 9172 18104 9178
rect 18052 9114 18104 9120
rect 17958 8936 18014 8945
rect 17958 8871 18014 8880
rect 17788 8486 17908 8514
rect 17406 6831 17462 6840
rect 17592 6860 17644 6866
rect 17316 6802 17368 6808
rect 17224 6792 17276 6798
rect 17224 6734 17276 6740
rect 17132 6656 17184 6662
rect 17132 6598 17184 6604
rect 17224 6656 17276 6662
rect 17224 6598 17276 6604
rect 17236 6474 17264 6598
rect 17144 6446 17264 6474
rect 17040 6248 17092 6254
rect 17040 6190 17092 6196
rect 16948 6180 17000 6186
rect 16948 6122 17000 6128
rect 16960 5574 16988 6122
rect 16948 5568 17000 5574
rect 16948 5510 17000 5516
rect 16854 5264 16910 5273
rect 16854 5199 16910 5208
rect 16948 5228 17000 5234
rect 16948 5170 17000 5176
rect 16960 4690 16988 5170
rect 16948 4684 17000 4690
rect 16948 4626 17000 4632
rect 16764 4208 16816 4214
rect 16764 4150 16816 4156
rect 16488 4140 16540 4146
rect 16488 4082 16540 4088
rect 16488 3936 16540 3942
rect 16488 3878 16540 3884
rect 16500 2553 16528 3878
rect 16960 3534 16988 4626
rect 17052 4622 17080 6190
rect 17144 5681 17172 6446
rect 17224 6384 17276 6390
rect 17224 6326 17276 6332
rect 17130 5672 17186 5681
rect 17130 5607 17186 5616
rect 17132 5568 17184 5574
rect 17132 5510 17184 5516
rect 17144 4826 17172 5510
rect 17132 4820 17184 4826
rect 17132 4762 17184 4768
rect 17040 4616 17092 4622
rect 17040 4558 17092 4564
rect 16948 3528 17000 3534
rect 17236 3482 17264 6326
rect 17328 5914 17356 6802
rect 17420 6390 17448 6831
rect 17592 6802 17644 6808
rect 17500 6792 17552 6798
rect 17500 6734 17552 6740
rect 17408 6384 17460 6390
rect 17512 6361 17540 6734
rect 17684 6656 17736 6662
rect 17684 6598 17736 6604
rect 17590 6488 17646 6497
rect 17590 6423 17646 6432
rect 17408 6326 17460 6332
rect 17498 6352 17554 6361
rect 17498 6287 17554 6296
rect 17408 6248 17460 6254
rect 17408 6190 17460 6196
rect 17316 5908 17368 5914
rect 17316 5850 17368 5856
rect 17420 5302 17448 6190
rect 17500 6112 17552 6118
rect 17500 6054 17552 6060
rect 17408 5296 17460 5302
rect 17314 5264 17370 5273
rect 17408 5238 17460 5244
rect 17314 5199 17370 5208
rect 16948 3470 17000 3476
rect 16486 2544 16542 2553
rect 16486 2479 16542 2488
rect 16580 2304 16632 2310
rect 16580 2246 16632 2252
rect 16304 1828 16356 1834
rect 16304 1770 16356 1776
rect 16592 56 16620 2246
rect 16960 474 16988 3470
rect 17052 3454 17264 3482
rect 17052 2582 17080 3454
rect 17132 3392 17184 3398
rect 17132 3334 17184 3340
rect 17224 3392 17276 3398
rect 17224 3334 17276 3340
rect 17040 2576 17092 2582
rect 17040 2518 17092 2524
rect 17144 1834 17172 3334
rect 17236 3126 17264 3334
rect 17224 3120 17276 3126
rect 17224 3062 17276 3068
rect 17132 1828 17184 1834
rect 17132 1770 17184 1776
rect 17328 1154 17356 5199
rect 17512 4185 17540 6054
rect 17604 5914 17632 6423
rect 17696 6118 17724 6598
rect 17684 6112 17736 6118
rect 17684 6054 17736 6060
rect 17592 5908 17644 5914
rect 17592 5850 17644 5856
rect 17788 5710 17816 8486
rect 18064 8401 18092 9114
rect 18050 8392 18106 8401
rect 18050 8327 18106 8336
rect 18156 8129 18184 11194
rect 18432 10878 18460 11194
rect 18420 10872 18472 10878
rect 18420 10814 18472 10820
rect 18604 9308 18656 9314
rect 18604 9250 18656 9256
rect 18236 8968 18288 8974
rect 18236 8910 18288 8916
rect 18248 8498 18276 8910
rect 18326 8800 18382 8809
rect 18326 8735 18382 8744
rect 18340 8634 18368 8735
rect 18328 8628 18380 8634
rect 18328 8570 18380 8576
rect 18420 8628 18472 8634
rect 18420 8570 18472 8576
rect 18236 8492 18288 8498
rect 18236 8434 18288 8440
rect 17958 8120 18014 8129
rect 17958 8055 18014 8064
rect 18142 8120 18198 8129
rect 18142 8055 18198 8064
rect 18328 8084 18380 8090
rect 17972 7970 18000 8055
rect 18328 8026 18380 8032
rect 17972 7942 18184 7970
rect 18052 7880 18104 7886
rect 18052 7822 18104 7828
rect 17960 7744 18012 7750
rect 17958 7712 17960 7721
rect 18012 7712 18014 7721
rect 17958 7647 18014 7656
rect 17868 7540 17920 7546
rect 17868 7482 17920 7488
rect 17880 7018 17908 7482
rect 18064 7478 18092 7822
rect 18052 7472 18104 7478
rect 18052 7414 18104 7420
rect 18156 7154 18184 7942
rect 18156 7126 18276 7154
rect 17880 6990 18000 7018
rect 18248 7002 18276 7126
rect 17972 6916 18000 6990
rect 18236 6996 18288 7002
rect 18236 6938 18288 6944
rect 18144 6928 18196 6934
rect 17972 6888 18144 6916
rect 18144 6870 18196 6876
rect 18236 6860 18288 6866
rect 18236 6802 18288 6808
rect 17960 6792 18012 6798
rect 17960 6734 18012 6740
rect 17868 6724 17920 6730
rect 17868 6666 17920 6672
rect 17880 6633 17908 6666
rect 17866 6624 17922 6633
rect 17866 6559 17922 6568
rect 17868 6384 17920 6390
rect 17868 6326 17920 6332
rect 17776 5704 17828 5710
rect 17776 5646 17828 5652
rect 17776 5568 17828 5574
rect 17776 5510 17828 5516
rect 17592 5296 17644 5302
rect 17592 5238 17644 5244
rect 17498 4176 17554 4185
rect 17498 4111 17554 4120
rect 17604 3602 17632 5238
rect 17684 4208 17736 4214
rect 17684 4150 17736 4156
rect 17592 3596 17644 3602
rect 17592 3538 17644 3544
rect 17498 3224 17554 3233
rect 17498 3159 17554 3168
rect 17512 2990 17540 3159
rect 17604 2990 17632 3538
rect 17500 2984 17552 2990
rect 17500 2926 17552 2932
rect 17592 2984 17644 2990
rect 17592 2926 17644 2932
rect 17500 2848 17552 2854
rect 17500 2790 17552 2796
rect 17512 2446 17540 2790
rect 17500 2440 17552 2446
rect 17500 2382 17552 2388
rect 17500 2304 17552 2310
rect 17500 2246 17552 2252
rect 17512 1465 17540 2246
rect 17498 1456 17554 1465
rect 17498 1391 17554 1400
rect 17316 1148 17368 1154
rect 17316 1090 17368 1096
rect 16948 468 17000 474
rect 16948 410 17000 416
rect 17696 56 17724 4150
rect 17788 3058 17816 5510
rect 17880 4010 17908 6326
rect 17972 4078 18000 6734
rect 18248 6458 18276 6802
rect 18340 6633 18368 8026
rect 18326 6624 18382 6633
rect 18326 6559 18382 6568
rect 18236 6452 18288 6458
rect 18236 6394 18288 6400
rect 18328 6452 18380 6458
rect 18328 6394 18380 6400
rect 18142 6352 18198 6361
rect 18198 6310 18276 6338
rect 18142 6287 18198 6296
rect 18144 6248 18196 6254
rect 18144 6190 18196 6196
rect 18156 6089 18184 6190
rect 18142 6080 18198 6089
rect 18142 6015 18198 6024
rect 18156 5273 18184 6015
rect 18142 5264 18198 5273
rect 18142 5199 18198 5208
rect 18052 4752 18104 4758
rect 18052 4694 18104 4700
rect 17960 4072 18012 4078
rect 17960 4014 18012 4020
rect 17868 4004 17920 4010
rect 17868 3946 17920 3952
rect 17960 3528 18012 3534
rect 17960 3470 18012 3476
rect 17776 3052 17828 3058
rect 17776 2994 17828 3000
rect 17868 2100 17920 2106
rect 17868 2042 17920 2048
rect 17880 1737 17908 2042
rect 17866 1728 17922 1737
rect 17866 1663 17922 1672
rect 17972 1630 18000 3470
rect 17960 1624 18012 1630
rect 17960 1566 18012 1572
rect 18064 678 18092 4694
rect 18248 4622 18276 6310
rect 18340 5710 18368 6394
rect 18432 6254 18460 8570
rect 18616 8362 18644 9250
rect 18708 8673 18736 11194
rect 18984 9858 19012 11194
rect 19064 10192 19116 10198
rect 19064 10134 19116 10140
rect 19076 9858 19104 10134
rect 19156 10124 19208 10130
rect 19156 10066 19208 10072
rect 18972 9852 19024 9858
rect 18972 9794 19024 9800
rect 19064 9852 19116 9858
rect 19064 9794 19116 9800
rect 18972 8900 19024 8906
rect 18972 8842 19024 8848
rect 18694 8664 18750 8673
rect 18694 8599 18750 8608
rect 18984 8498 19012 8842
rect 18972 8492 19024 8498
rect 18972 8434 19024 8440
rect 19064 8492 19116 8498
rect 19064 8434 19116 8440
rect 18696 8424 18748 8430
rect 18696 8366 18748 8372
rect 18604 8356 18656 8362
rect 18604 8298 18656 8304
rect 18604 8084 18656 8090
rect 18604 8026 18656 8032
rect 18512 7948 18564 7954
rect 18512 7890 18564 7896
rect 18524 7546 18552 7890
rect 18616 7886 18644 8026
rect 18604 7880 18656 7886
rect 18604 7822 18656 7828
rect 18512 7540 18564 7546
rect 18512 7482 18564 7488
rect 18604 7540 18656 7546
rect 18604 7482 18656 7488
rect 18616 7206 18644 7482
rect 18604 7200 18656 7206
rect 18510 7168 18566 7177
rect 18604 7142 18656 7148
rect 18510 7103 18566 7112
rect 18524 7018 18552 7103
rect 18524 6990 18644 7018
rect 18512 6928 18564 6934
rect 18510 6896 18512 6905
rect 18564 6896 18566 6905
rect 18616 6866 18644 6990
rect 18510 6831 18566 6840
rect 18604 6860 18656 6866
rect 18604 6802 18656 6808
rect 18510 6760 18566 6769
rect 18510 6695 18566 6704
rect 18420 6248 18472 6254
rect 18420 6190 18472 6196
rect 18524 6202 18552 6695
rect 18602 6624 18658 6633
rect 18602 6559 18658 6568
rect 18616 6322 18644 6559
rect 18604 6316 18656 6322
rect 18604 6258 18656 6264
rect 18524 6174 18644 6202
rect 18420 6112 18472 6118
rect 18420 6054 18472 6060
rect 18512 6112 18564 6118
rect 18616 6089 18644 6174
rect 18512 6054 18564 6060
rect 18602 6080 18658 6089
rect 18432 5778 18460 6054
rect 18524 5846 18552 6054
rect 18602 6015 18658 6024
rect 18512 5840 18564 5846
rect 18512 5782 18564 5788
rect 18420 5772 18472 5778
rect 18420 5714 18472 5720
rect 18328 5704 18380 5710
rect 18328 5646 18380 5652
rect 18328 5568 18380 5574
rect 18328 5510 18380 5516
rect 18512 5568 18564 5574
rect 18512 5510 18564 5516
rect 18340 5370 18368 5510
rect 18328 5364 18380 5370
rect 18328 5306 18380 5312
rect 18236 4616 18288 4622
rect 18236 4558 18288 4564
rect 18328 4480 18380 4486
rect 18328 4422 18380 4428
rect 18236 4276 18288 4282
rect 18236 4218 18288 4224
rect 18248 4078 18276 4218
rect 18340 4146 18368 4422
rect 18328 4140 18380 4146
rect 18328 4082 18380 4088
rect 18236 4072 18288 4078
rect 18236 4014 18288 4020
rect 18328 3936 18380 3942
rect 18328 3878 18380 3884
rect 18234 3768 18290 3777
rect 18234 3703 18290 3712
rect 18248 3670 18276 3703
rect 18236 3664 18288 3670
rect 18236 3606 18288 3612
rect 18236 3528 18288 3534
rect 18236 3470 18288 3476
rect 18248 3398 18276 3470
rect 18236 3392 18288 3398
rect 18236 3334 18288 3340
rect 18340 2990 18368 3878
rect 18524 3534 18552 5510
rect 18708 5370 18736 8366
rect 18972 8356 19024 8362
rect 18972 8298 19024 8304
rect 18878 8120 18934 8129
rect 18878 8055 18934 8064
rect 18892 7886 18920 8055
rect 18984 7936 19012 8298
rect 19076 8129 19104 8434
rect 19062 8120 19118 8129
rect 19062 8055 19118 8064
rect 18984 7908 19104 7936
rect 18880 7880 18932 7886
rect 18880 7822 18932 7828
rect 18972 7744 19024 7750
rect 18892 7704 18972 7732
rect 18892 7698 18920 7704
rect 18857 7670 18920 7698
rect 18972 7686 19024 7692
rect 18857 7562 18885 7670
rect 18800 7534 18885 7562
rect 18800 7426 18828 7534
rect 18800 7398 19012 7426
rect 19076 7410 19104 7908
rect 18788 7268 18840 7274
rect 18840 7228 18920 7256
rect 18788 7210 18840 7216
rect 18786 7032 18842 7041
rect 18786 6967 18842 6976
rect 18800 5710 18828 6967
rect 18892 5778 18920 7228
rect 18880 5772 18932 5778
rect 18880 5714 18932 5720
rect 18788 5704 18840 5710
rect 18788 5646 18840 5652
rect 18788 5568 18840 5574
rect 18788 5510 18840 5516
rect 18696 5364 18748 5370
rect 18696 5306 18748 5312
rect 18694 5264 18750 5273
rect 18694 5199 18750 5208
rect 18708 4622 18736 5199
rect 18696 4616 18748 4622
rect 18696 4558 18748 4564
rect 18800 4162 18828 5510
rect 18984 5234 19012 7398
rect 19064 7404 19116 7410
rect 19064 7346 19116 7352
rect 19064 6928 19116 6934
rect 19062 6896 19064 6905
rect 19116 6896 19118 6905
rect 19062 6831 19118 6840
rect 19168 6798 19196 10066
rect 19156 6792 19208 6798
rect 19156 6734 19208 6740
rect 19062 6488 19118 6497
rect 19062 6423 19118 6432
rect 19076 6186 19104 6423
rect 19260 6322 19288 11194
rect 19536 9761 19564 11194
rect 19522 9752 19578 9761
rect 19522 9687 19578 9696
rect 19812 9330 19840 11194
rect 19628 9302 19840 9330
rect 19524 8356 19576 8362
rect 19524 8298 19576 8304
rect 19430 8256 19486 8265
rect 19430 8191 19486 8200
rect 19444 7818 19472 8191
rect 19340 7812 19392 7818
rect 19340 7754 19392 7760
rect 19432 7812 19484 7818
rect 19432 7754 19484 7760
rect 19248 6316 19300 6322
rect 19248 6258 19300 6264
rect 19064 6180 19116 6186
rect 19064 6122 19116 6128
rect 19248 6112 19300 6118
rect 19246 6080 19248 6089
rect 19300 6080 19302 6089
rect 19246 6015 19302 6024
rect 19352 5710 19380 7754
rect 19432 6724 19484 6730
rect 19432 6666 19484 6672
rect 19444 6118 19472 6666
rect 19432 6112 19484 6118
rect 19432 6054 19484 6060
rect 19430 5944 19486 5953
rect 19430 5879 19486 5888
rect 19340 5704 19392 5710
rect 19340 5646 19392 5652
rect 19064 5568 19116 5574
rect 19064 5510 19116 5516
rect 18972 5228 19024 5234
rect 18972 5170 19024 5176
rect 19076 5114 19104 5510
rect 19444 5370 19472 5879
rect 19432 5364 19484 5370
rect 19432 5306 19484 5312
rect 19338 5264 19394 5273
rect 19156 5228 19208 5234
rect 19338 5199 19394 5208
rect 19156 5170 19208 5176
rect 18616 4134 18828 4162
rect 18984 5086 19104 5114
rect 19168 5098 19196 5170
rect 19352 5098 19380 5199
rect 19432 5160 19484 5166
rect 19432 5102 19484 5108
rect 19156 5092 19208 5098
rect 18512 3528 18564 3534
rect 18512 3470 18564 3476
rect 18512 3392 18564 3398
rect 18432 3352 18512 3380
rect 18328 2984 18380 2990
rect 18328 2926 18380 2932
rect 18236 2916 18288 2922
rect 18236 2858 18288 2864
rect 18248 2650 18276 2858
rect 18236 2644 18288 2650
rect 18236 2586 18288 2592
rect 18340 2514 18368 2926
rect 18328 2508 18380 2514
rect 18328 2450 18380 2456
rect 18340 2106 18368 2450
rect 18328 2100 18380 2106
rect 18328 2042 18380 2048
rect 18432 814 18460 3352
rect 18512 3334 18564 3340
rect 18616 2774 18644 4134
rect 18984 4078 19012 5086
rect 19156 5034 19208 5040
rect 19340 5092 19392 5098
rect 19340 5034 19392 5040
rect 19064 5024 19116 5030
rect 19064 4966 19116 4972
rect 18880 4072 18932 4078
rect 18880 4014 18932 4020
rect 18972 4072 19024 4078
rect 18972 4014 19024 4020
rect 18892 3942 18920 4014
rect 18788 3936 18840 3942
rect 18788 3878 18840 3884
rect 18880 3936 18932 3942
rect 18880 3878 18932 3884
rect 18800 3534 18828 3878
rect 18972 3596 19024 3602
rect 18972 3538 19024 3544
rect 18788 3528 18840 3534
rect 18694 3496 18750 3505
rect 18788 3470 18840 3476
rect 18878 3496 18934 3505
rect 18694 3431 18750 3440
rect 18878 3431 18934 3440
rect 18708 3398 18736 3431
rect 18696 3392 18748 3398
rect 18696 3334 18748 3340
rect 18786 3224 18842 3233
rect 18786 3159 18842 3168
rect 18800 3058 18828 3159
rect 18788 3052 18840 3058
rect 18788 2994 18840 3000
rect 18694 2952 18750 2961
rect 18694 2887 18750 2896
rect 18524 2746 18644 2774
rect 18524 2689 18552 2746
rect 18510 2680 18566 2689
rect 18510 2615 18566 2624
rect 18708 2446 18736 2887
rect 18696 2440 18748 2446
rect 18696 2382 18748 2388
rect 18892 1714 18920 3431
rect 18984 2514 19012 3538
rect 19076 3534 19104 4966
rect 19248 4752 19300 4758
rect 19248 4694 19300 4700
rect 19156 3664 19208 3670
rect 19156 3606 19208 3612
rect 19064 3528 19116 3534
rect 19064 3470 19116 3476
rect 19168 3369 19196 3606
rect 19154 3360 19210 3369
rect 19154 3295 19210 3304
rect 19260 2922 19288 4694
rect 19444 4690 19472 5102
rect 19432 4684 19484 4690
rect 19432 4626 19484 4632
rect 19536 4146 19564 8298
rect 19628 7546 19656 9302
rect 20088 8480 20116 11194
rect 20364 9058 20392 11194
rect 20364 9030 20484 9058
rect 19720 8452 20116 8480
rect 19616 7540 19668 7546
rect 19616 7482 19668 7488
rect 19616 6792 19668 6798
rect 19616 6734 19668 6740
rect 19628 5234 19656 6734
rect 19720 5642 19748 8452
rect 20352 8424 20404 8430
rect 20352 8366 20404 8372
rect 19950 8188 20258 8197
rect 19950 8186 19956 8188
rect 20012 8186 20036 8188
rect 20092 8186 20116 8188
rect 20172 8186 20196 8188
rect 20252 8186 20258 8188
rect 20012 8134 20014 8186
rect 20194 8134 20196 8186
rect 19950 8132 19956 8134
rect 20012 8132 20036 8134
rect 20092 8132 20116 8134
rect 20172 8132 20196 8134
rect 20252 8132 20258 8134
rect 19950 8123 20258 8132
rect 20168 8084 20220 8090
rect 20168 8026 20220 8032
rect 20180 7818 20208 8026
rect 20260 7880 20312 7886
rect 20260 7822 20312 7828
rect 20168 7812 20220 7818
rect 20168 7754 20220 7760
rect 19800 7744 19852 7750
rect 19800 7686 19852 7692
rect 19708 5636 19760 5642
rect 19708 5578 19760 5584
rect 19616 5228 19668 5234
rect 19616 5170 19668 5176
rect 19524 4140 19576 4146
rect 19524 4082 19576 4088
rect 19708 3596 19760 3602
rect 19708 3538 19760 3544
rect 19340 3392 19392 3398
rect 19340 3334 19392 3340
rect 19248 2916 19300 2922
rect 19248 2858 19300 2864
rect 18972 2508 19024 2514
rect 18972 2450 19024 2456
rect 19246 2408 19302 2417
rect 19246 2343 19302 2352
rect 19260 2310 19288 2343
rect 19248 2304 19300 2310
rect 19248 2246 19300 2252
rect 19352 2009 19380 3334
rect 19432 3120 19484 3126
rect 19432 3062 19484 3068
rect 19444 2961 19472 3062
rect 19720 3058 19748 3538
rect 19708 3052 19760 3058
rect 19708 2994 19760 3000
rect 19430 2952 19486 2961
rect 19430 2887 19486 2896
rect 19432 2848 19484 2854
rect 19432 2790 19484 2796
rect 19444 2446 19472 2790
rect 19432 2440 19484 2446
rect 19432 2382 19484 2388
rect 19338 2000 19394 2009
rect 19338 1935 19394 1944
rect 19812 1873 19840 7686
rect 20180 7206 20208 7754
rect 20272 7392 20300 7822
rect 20364 7818 20392 8366
rect 20352 7812 20404 7818
rect 20352 7754 20404 7760
rect 20352 7404 20404 7410
rect 20272 7364 20352 7392
rect 20352 7346 20404 7352
rect 20168 7200 20220 7206
rect 20168 7142 20220 7148
rect 19950 7100 20258 7109
rect 19950 7098 19956 7100
rect 20012 7098 20036 7100
rect 20092 7098 20116 7100
rect 20172 7098 20196 7100
rect 20252 7098 20258 7100
rect 20012 7046 20014 7098
rect 20194 7046 20196 7098
rect 19950 7044 19956 7046
rect 20012 7044 20036 7046
rect 20092 7044 20116 7046
rect 20172 7044 20196 7046
rect 20252 7044 20258 7046
rect 19950 7035 20258 7044
rect 20364 6866 20392 7346
rect 20456 6905 20484 9030
rect 20536 9036 20588 9042
rect 20536 8978 20588 8984
rect 20442 6896 20498 6905
rect 20352 6860 20404 6866
rect 20442 6831 20498 6840
rect 20352 6802 20404 6808
rect 20260 6724 20312 6730
rect 20312 6684 20392 6712
rect 20260 6666 20312 6672
rect 20364 6089 20392 6684
rect 20350 6080 20406 6089
rect 19950 6012 20258 6021
rect 20350 6015 20406 6024
rect 19950 6010 19956 6012
rect 20012 6010 20036 6012
rect 20092 6010 20116 6012
rect 20172 6010 20196 6012
rect 20252 6010 20258 6012
rect 20012 5958 20014 6010
rect 20194 5958 20196 6010
rect 19950 5956 19956 5958
rect 20012 5956 20036 5958
rect 20092 5956 20116 5958
rect 20172 5956 20196 5958
rect 20252 5956 20258 5958
rect 19950 5947 20258 5956
rect 20364 5166 20392 6015
rect 20444 5228 20496 5234
rect 20444 5170 20496 5176
rect 20352 5160 20404 5166
rect 20352 5102 20404 5108
rect 19950 4924 20258 4933
rect 19950 4922 19956 4924
rect 20012 4922 20036 4924
rect 20092 4922 20116 4924
rect 20172 4922 20196 4924
rect 20252 4922 20258 4924
rect 20012 4870 20014 4922
rect 20194 4870 20196 4922
rect 19950 4868 19956 4870
rect 20012 4868 20036 4870
rect 20092 4868 20116 4870
rect 20172 4868 20196 4870
rect 20252 4868 20258 4870
rect 19950 4859 20258 4868
rect 20456 4622 20484 5170
rect 20444 4616 20496 4622
rect 20444 4558 20496 4564
rect 20548 4486 20576 8978
rect 20640 6322 20668 11194
rect 20916 10130 20944 11194
rect 20996 10532 21048 10538
rect 20996 10474 21048 10480
rect 21008 10130 21036 10474
rect 20904 10124 20956 10130
rect 20904 10066 20956 10072
rect 20996 10124 21048 10130
rect 20996 10066 21048 10072
rect 21192 9874 21220 11194
rect 20916 9846 21220 9874
rect 20916 8498 20944 9846
rect 21010 8732 21318 8741
rect 21010 8730 21016 8732
rect 21072 8730 21096 8732
rect 21152 8730 21176 8732
rect 21232 8730 21256 8732
rect 21312 8730 21318 8732
rect 21072 8678 21074 8730
rect 21254 8678 21256 8730
rect 21010 8676 21016 8678
rect 21072 8676 21096 8678
rect 21152 8676 21176 8678
rect 21232 8676 21256 8678
rect 21312 8676 21318 8678
rect 21010 8667 21318 8676
rect 21468 8498 21496 11194
rect 21548 8832 21600 8838
rect 21548 8774 21600 8780
rect 20904 8492 20956 8498
rect 20904 8434 20956 8440
rect 21456 8492 21508 8498
rect 21456 8434 21508 8440
rect 21088 8424 21140 8430
rect 21088 8366 21140 8372
rect 21364 8424 21416 8430
rect 21364 8366 21416 8372
rect 20904 8288 20956 8294
rect 20904 8230 20956 8236
rect 20810 7712 20866 7721
rect 20810 7647 20866 7656
rect 20718 7576 20774 7585
rect 20718 7511 20774 7520
rect 20732 7313 20760 7511
rect 20718 7304 20774 7313
rect 20718 7239 20774 7248
rect 20824 7177 20852 7647
rect 20810 7168 20866 7177
rect 20810 7103 20866 7112
rect 20628 6316 20680 6322
rect 20628 6258 20680 6264
rect 20626 5944 20682 5953
rect 20626 5879 20682 5888
rect 20720 5908 20772 5914
rect 20640 5681 20668 5879
rect 20720 5850 20772 5856
rect 20626 5672 20682 5681
rect 20626 5607 20682 5616
rect 20640 4690 20668 5607
rect 20628 4684 20680 4690
rect 20628 4626 20680 4632
rect 20444 4480 20496 4486
rect 20444 4422 20496 4428
rect 20536 4480 20588 4486
rect 20536 4422 20588 4428
rect 19950 3836 20258 3845
rect 19950 3834 19956 3836
rect 20012 3834 20036 3836
rect 20092 3834 20116 3836
rect 20172 3834 20196 3836
rect 20252 3834 20258 3836
rect 20012 3782 20014 3834
rect 20194 3782 20196 3834
rect 19950 3780 19956 3782
rect 20012 3780 20036 3782
rect 20092 3780 20116 3782
rect 20172 3780 20196 3782
rect 20252 3780 20258 3782
rect 19950 3771 20258 3780
rect 20352 3664 20404 3670
rect 20352 3606 20404 3612
rect 20364 3058 20392 3606
rect 20352 3052 20404 3058
rect 20352 2994 20404 3000
rect 20352 2916 20404 2922
rect 20352 2858 20404 2864
rect 20364 2825 20392 2858
rect 20350 2816 20406 2825
rect 19950 2748 20258 2757
rect 20350 2751 20406 2760
rect 19950 2746 19956 2748
rect 20012 2746 20036 2748
rect 20092 2746 20116 2748
rect 20172 2746 20196 2748
rect 20252 2746 20258 2748
rect 20012 2694 20014 2746
rect 20194 2694 20196 2746
rect 19950 2692 19956 2694
rect 20012 2692 20036 2694
rect 20092 2692 20116 2694
rect 20172 2692 20196 2694
rect 20252 2692 20258 2694
rect 19950 2683 20258 2692
rect 19892 2440 19944 2446
rect 19892 2382 19944 2388
rect 19798 1864 19854 1873
rect 19798 1799 19854 1808
rect 18800 1686 18920 1714
rect 18420 808 18472 814
rect 18420 750 18472 756
rect 18052 672 18104 678
rect 18052 614 18104 620
rect 18800 56 18828 1686
rect 19904 56 19932 2382
rect 20456 1970 20484 4422
rect 20732 4214 20760 5850
rect 20916 4842 20944 8230
rect 20994 7984 21050 7993
rect 20994 7919 21050 7928
rect 21008 7750 21036 7919
rect 21100 7750 21128 8366
rect 20996 7744 21048 7750
rect 20996 7686 21048 7692
rect 21088 7744 21140 7750
rect 21088 7686 21140 7692
rect 21010 7644 21318 7653
rect 21010 7642 21016 7644
rect 21072 7642 21096 7644
rect 21152 7642 21176 7644
rect 21232 7642 21256 7644
rect 21312 7642 21318 7644
rect 21072 7590 21074 7642
rect 21254 7590 21256 7642
rect 21010 7588 21016 7590
rect 21072 7588 21096 7590
rect 21152 7588 21176 7590
rect 21232 7588 21256 7590
rect 21312 7588 21318 7590
rect 21010 7579 21318 7588
rect 21376 7410 21404 8366
rect 21456 7948 21508 7954
rect 21456 7890 21508 7896
rect 21468 7585 21496 7890
rect 21454 7576 21510 7585
rect 21454 7511 21510 7520
rect 21364 7404 21416 7410
rect 21364 7346 21416 7352
rect 21364 6792 21416 6798
rect 21364 6734 21416 6740
rect 21010 6556 21318 6565
rect 21010 6554 21016 6556
rect 21072 6554 21096 6556
rect 21152 6554 21176 6556
rect 21232 6554 21256 6556
rect 21312 6554 21318 6556
rect 21072 6502 21074 6554
rect 21254 6502 21256 6554
rect 21010 6500 21016 6502
rect 21072 6500 21096 6502
rect 21152 6500 21176 6502
rect 21232 6500 21256 6502
rect 21312 6500 21318 6502
rect 21010 6491 21318 6500
rect 21376 6390 21404 6734
rect 21560 6440 21588 8774
rect 21640 8424 21692 8430
rect 21640 8366 21692 8372
rect 21652 7546 21680 8366
rect 21744 8362 21772 11194
rect 21822 9208 21878 9217
rect 21822 9143 21878 9152
rect 21732 8356 21784 8362
rect 21732 8298 21784 8304
rect 21640 7540 21692 7546
rect 21640 7482 21692 7488
rect 21732 6656 21784 6662
rect 21732 6598 21784 6604
rect 21468 6412 21588 6440
rect 21364 6384 21416 6390
rect 21364 6326 21416 6332
rect 21468 6118 21496 6412
rect 21548 6316 21600 6322
rect 21548 6258 21600 6264
rect 21456 6112 21508 6118
rect 21456 6054 21508 6060
rect 21364 5636 21416 5642
rect 21364 5578 21416 5584
rect 21010 5468 21318 5477
rect 21010 5466 21016 5468
rect 21072 5466 21096 5468
rect 21152 5466 21176 5468
rect 21232 5466 21256 5468
rect 21312 5466 21318 5468
rect 21072 5414 21074 5466
rect 21254 5414 21256 5466
rect 21010 5412 21016 5414
rect 21072 5412 21096 5414
rect 21152 5412 21176 5414
rect 21232 5412 21256 5414
rect 21312 5412 21318 5414
rect 21010 5403 21318 5412
rect 21180 5296 21232 5302
rect 21180 5238 21232 5244
rect 21192 4865 21220 5238
rect 21272 5024 21324 5030
rect 21270 4992 21272 5001
rect 21324 4992 21326 5001
rect 21270 4927 21326 4936
rect 21178 4856 21234 4865
rect 20916 4814 21036 4842
rect 20904 4752 20956 4758
rect 20904 4694 20956 4700
rect 20812 4616 20864 4622
rect 20812 4558 20864 4564
rect 20720 4208 20772 4214
rect 20720 4150 20772 4156
rect 20720 4072 20772 4078
rect 20720 4014 20772 4020
rect 20732 3738 20760 4014
rect 20824 4010 20852 4558
rect 20916 4060 20944 4694
rect 21008 4486 21036 4814
rect 21178 4791 21234 4800
rect 20996 4480 21048 4486
rect 20996 4422 21048 4428
rect 21010 4380 21318 4389
rect 21010 4378 21016 4380
rect 21072 4378 21096 4380
rect 21152 4378 21176 4380
rect 21232 4378 21256 4380
rect 21312 4378 21318 4380
rect 21072 4326 21074 4378
rect 21254 4326 21256 4378
rect 21010 4324 21016 4326
rect 21072 4324 21096 4326
rect 21152 4324 21176 4326
rect 21232 4324 21256 4326
rect 21312 4324 21318 4326
rect 21010 4315 21318 4324
rect 20996 4072 21048 4078
rect 20916 4032 20996 4060
rect 20996 4014 21048 4020
rect 21376 4010 21404 5578
rect 21456 5568 21508 5574
rect 21456 5510 21508 5516
rect 21468 5302 21496 5510
rect 21560 5370 21588 6258
rect 21640 5704 21692 5710
rect 21640 5646 21692 5652
rect 21548 5364 21600 5370
rect 21548 5306 21600 5312
rect 21456 5296 21508 5302
rect 21456 5238 21508 5244
rect 21652 5148 21680 5646
rect 21468 5120 21680 5148
rect 21468 4826 21496 5120
rect 21744 5030 21772 6598
rect 21548 5024 21600 5030
rect 21548 4966 21600 4972
rect 21640 5024 21692 5030
rect 21640 4966 21692 4972
rect 21732 5024 21784 5030
rect 21732 4966 21784 4972
rect 21456 4820 21508 4826
rect 21456 4762 21508 4768
rect 21560 4690 21588 4966
rect 21652 4690 21680 4966
rect 21548 4684 21600 4690
rect 21548 4626 21600 4632
rect 21640 4684 21692 4690
rect 21640 4626 21692 4632
rect 21548 4480 21600 4486
rect 21548 4422 21600 4428
rect 20812 4004 20864 4010
rect 20812 3946 20864 3952
rect 21364 4004 21416 4010
rect 21364 3946 21416 3952
rect 20994 3768 21050 3777
rect 20720 3732 20772 3738
rect 20994 3703 20996 3712
rect 20720 3674 20772 3680
rect 21048 3703 21050 3712
rect 20996 3674 21048 3680
rect 21364 3528 21416 3534
rect 21364 3470 21416 3476
rect 21456 3528 21508 3534
rect 21456 3470 21508 3476
rect 21010 3292 21318 3301
rect 21010 3290 21016 3292
rect 21072 3290 21096 3292
rect 21152 3290 21176 3292
rect 21232 3290 21256 3292
rect 21312 3290 21318 3292
rect 21072 3238 21074 3290
rect 21254 3238 21256 3290
rect 21010 3236 21016 3238
rect 21072 3236 21096 3238
rect 21152 3236 21176 3238
rect 21232 3236 21256 3238
rect 21312 3236 21318 3238
rect 21010 3227 21318 3236
rect 20904 3120 20956 3126
rect 20732 3068 20904 3074
rect 20732 3062 20956 3068
rect 20732 3058 20944 3062
rect 20720 3052 20944 3058
rect 20772 3046 20944 3052
rect 20720 2994 20772 3000
rect 21376 2650 21404 3470
rect 21468 3058 21496 3470
rect 21456 3052 21508 3058
rect 21456 2994 21508 3000
rect 21456 2848 21508 2854
rect 21456 2790 21508 2796
rect 21364 2644 21416 2650
rect 21364 2586 21416 2592
rect 21468 2514 21496 2790
rect 21456 2508 21508 2514
rect 21456 2450 21508 2456
rect 20904 2440 20956 2446
rect 20904 2382 20956 2388
rect 21086 2408 21142 2417
rect 20812 2304 20864 2310
rect 20812 2246 20864 2252
rect 20444 1964 20496 1970
rect 20444 1906 20496 1912
rect 20824 1902 20852 2246
rect 20812 1896 20864 1902
rect 20812 1838 20864 1844
rect 20916 1170 20944 2382
rect 21086 2343 21142 2352
rect 21100 2310 21128 2343
rect 21560 2310 21588 4422
rect 21640 3392 21692 3398
rect 21640 3334 21692 3340
rect 21652 2514 21680 3334
rect 21836 3126 21864 9143
rect 21916 7880 21968 7886
rect 21916 7822 21968 7828
rect 21928 4690 21956 7822
rect 22020 6934 22048 11194
rect 22100 7540 22152 7546
rect 22100 7482 22152 7488
rect 22008 6928 22060 6934
rect 22008 6870 22060 6876
rect 22008 6656 22060 6662
rect 22008 6598 22060 6604
rect 22020 6202 22048 6598
rect 22112 6322 22140 7482
rect 22192 7200 22244 7206
rect 22192 7142 22244 7148
rect 22204 6390 22232 7142
rect 22296 7002 22324 11194
rect 22466 10432 22522 10441
rect 22376 10396 22428 10402
rect 22466 10367 22522 10376
rect 22376 10338 22428 10344
rect 22388 8022 22416 10338
rect 22480 10033 22508 10367
rect 22466 10024 22522 10033
rect 22466 9959 22522 9968
rect 22572 9761 22600 11194
rect 22848 9897 22876 11194
rect 23020 10464 23072 10470
rect 23020 10406 23072 10412
rect 22834 9888 22890 9897
rect 22834 9823 22890 9832
rect 22558 9752 22614 9761
rect 22558 9687 22614 9696
rect 22744 9376 22796 9382
rect 22744 9318 22796 9324
rect 22756 8378 22784 9318
rect 22836 9308 22888 9314
rect 22836 9250 22888 9256
rect 22848 8838 22876 9250
rect 22836 8832 22888 8838
rect 22836 8774 22888 8780
rect 22848 8498 22876 8774
rect 22836 8492 22888 8498
rect 22836 8434 22888 8440
rect 22928 8424 22980 8430
rect 22756 8350 22876 8378
rect 22928 8366 22980 8372
rect 22376 8016 22428 8022
rect 22376 7958 22428 7964
rect 22560 7812 22612 7818
rect 22560 7754 22612 7760
rect 22466 7712 22522 7721
rect 22466 7647 22522 7656
rect 22376 7268 22428 7274
rect 22376 7210 22428 7216
rect 22284 6996 22336 7002
rect 22284 6938 22336 6944
rect 22284 6860 22336 6866
rect 22284 6802 22336 6808
rect 22296 6730 22324 6802
rect 22284 6724 22336 6730
rect 22284 6666 22336 6672
rect 22192 6384 22244 6390
rect 22192 6326 22244 6332
rect 22100 6316 22152 6322
rect 22100 6258 22152 6264
rect 22020 6174 22140 6202
rect 22008 5772 22060 5778
rect 22008 5714 22060 5720
rect 22020 5574 22048 5714
rect 22008 5568 22060 5574
rect 22008 5510 22060 5516
rect 22112 5166 22140 6174
rect 22284 6180 22336 6186
rect 22284 6122 22336 6128
rect 22296 5778 22324 6122
rect 22284 5772 22336 5778
rect 22284 5714 22336 5720
rect 22388 5250 22416 7210
rect 22480 6322 22508 7647
rect 22468 6316 22520 6322
rect 22468 6258 22520 6264
rect 22572 6186 22600 7754
rect 22744 7744 22796 7750
rect 22744 7686 22796 7692
rect 22652 7404 22704 7410
rect 22652 7346 22704 7352
rect 22664 7206 22692 7346
rect 22652 7200 22704 7206
rect 22652 7142 22704 7148
rect 22756 6798 22784 7686
rect 22744 6792 22796 6798
rect 22744 6734 22796 6740
rect 22652 6656 22704 6662
rect 22652 6598 22704 6604
rect 22664 6390 22692 6598
rect 22652 6384 22704 6390
rect 22652 6326 22704 6332
rect 22560 6180 22612 6186
rect 22560 6122 22612 6128
rect 22664 5778 22692 6326
rect 22652 5772 22704 5778
rect 22652 5714 22704 5720
rect 22468 5704 22520 5710
rect 22468 5646 22520 5652
rect 22204 5222 22416 5250
rect 22100 5160 22152 5166
rect 22100 5102 22152 5108
rect 21916 4684 21968 4690
rect 21916 4626 21968 4632
rect 21824 3120 21876 3126
rect 21824 3062 21876 3068
rect 21928 2961 21956 4626
rect 22204 4282 22232 5222
rect 22376 5160 22428 5166
rect 22376 5102 22428 5108
rect 22284 5024 22336 5030
rect 22388 5001 22416 5102
rect 22284 4966 22336 4972
rect 22374 4992 22430 5001
rect 22296 4690 22324 4966
rect 22374 4927 22430 4936
rect 22284 4684 22336 4690
rect 22284 4626 22336 4632
rect 22480 4457 22508 5646
rect 22466 4448 22522 4457
rect 22466 4383 22522 4392
rect 22374 4312 22430 4321
rect 22192 4276 22244 4282
rect 22374 4247 22430 4256
rect 22192 4218 22244 4224
rect 22388 4078 22416 4247
rect 22480 4078 22508 4383
rect 22376 4072 22428 4078
rect 22376 4014 22428 4020
rect 22468 4072 22520 4078
rect 22468 4014 22520 4020
rect 22100 3528 22152 3534
rect 22100 3470 22152 3476
rect 22112 3398 22140 3470
rect 22100 3392 22152 3398
rect 22100 3334 22152 3340
rect 22008 2984 22060 2990
rect 21914 2952 21970 2961
rect 22112 2972 22140 3334
rect 22060 2944 22140 2972
rect 22008 2926 22060 2932
rect 21914 2887 21970 2896
rect 22848 2774 22876 8350
rect 22940 7478 22968 8366
rect 23032 8106 23060 10406
rect 23124 9330 23152 11194
rect 23400 10169 23428 11194
rect 23572 10192 23624 10198
rect 23386 10160 23442 10169
rect 23572 10134 23624 10140
rect 23386 10095 23442 10104
rect 23584 9858 23612 10134
rect 23572 9852 23624 9858
rect 23572 9794 23624 9800
rect 23676 9450 23704 11194
rect 23664 9444 23716 9450
rect 23664 9386 23716 9392
rect 23124 9302 23520 9330
rect 23204 8560 23256 8566
rect 23204 8502 23256 8508
rect 23294 8528 23350 8537
rect 23216 8430 23244 8502
rect 23294 8463 23350 8472
rect 23204 8424 23256 8430
rect 23204 8366 23256 8372
rect 23112 8288 23164 8294
rect 23110 8256 23112 8265
rect 23204 8288 23256 8294
rect 23164 8256 23166 8265
rect 23204 8230 23256 8236
rect 23110 8191 23166 8200
rect 23032 8078 23152 8106
rect 23020 8016 23072 8022
rect 23020 7958 23072 7964
rect 22928 7472 22980 7478
rect 22928 7414 22980 7420
rect 22928 6792 22980 6798
rect 22928 6734 22980 6740
rect 22940 6662 22968 6734
rect 22928 6656 22980 6662
rect 23032 6644 23060 7958
rect 23124 6746 23152 8078
rect 23216 7478 23244 8230
rect 23308 7546 23336 8463
rect 23388 8356 23440 8362
rect 23388 8298 23440 8304
rect 23296 7540 23348 7546
rect 23296 7482 23348 7488
rect 23204 7472 23256 7478
rect 23204 7414 23256 7420
rect 23400 7410 23428 8298
rect 23492 7546 23520 9302
rect 23664 9308 23716 9314
rect 23664 9250 23716 9256
rect 23572 8424 23624 8430
rect 23572 8366 23624 8372
rect 23584 7721 23612 8366
rect 23570 7712 23626 7721
rect 23570 7647 23626 7656
rect 23480 7540 23532 7546
rect 23480 7482 23532 7488
rect 23388 7404 23440 7410
rect 23388 7346 23440 7352
rect 23572 6996 23624 7002
rect 23572 6938 23624 6944
rect 23478 6896 23534 6905
rect 23478 6831 23534 6840
rect 23492 6798 23520 6831
rect 23584 6798 23612 6938
rect 23480 6792 23532 6798
rect 23124 6718 23336 6746
rect 23480 6734 23532 6740
rect 23572 6792 23624 6798
rect 23572 6734 23624 6740
rect 23112 6656 23164 6662
rect 23032 6616 23112 6644
rect 22928 6598 22980 6604
rect 23112 6598 23164 6604
rect 23112 6316 23164 6322
rect 23112 6258 23164 6264
rect 22928 6112 22980 6118
rect 22928 6054 22980 6060
rect 23020 6112 23072 6118
rect 23020 6054 23072 6060
rect 22940 5658 22968 6054
rect 23032 5953 23060 6054
rect 23018 5944 23074 5953
rect 23018 5879 23074 5888
rect 23124 5846 23152 6258
rect 23112 5840 23164 5846
rect 23112 5782 23164 5788
rect 23112 5704 23164 5710
rect 22940 5630 23060 5658
rect 23112 5646 23164 5652
rect 23202 5672 23258 5681
rect 23032 5234 23060 5630
rect 23020 5228 23072 5234
rect 23020 5170 23072 5176
rect 23124 4826 23152 5646
rect 23202 5607 23258 5616
rect 23216 5574 23244 5607
rect 23204 5568 23256 5574
rect 23204 5510 23256 5516
rect 23204 5296 23256 5302
rect 23204 5238 23256 5244
rect 23112 4820 23164 4826
rect 23112 4762 23164 4768
rect 22928 4752 22980 4758
rect 22928 4694 22980 4700
rect 22940 3942 22968 4694
rect 23216 4298 23244 5238
rect 23308 5030 23336 6718
rect 23492 6322 23520 6734
rect 23480 6316 23532 6322
rect 23480 6258 23532 6264
rect 23388 6248 23440 6254
rect 23388 6190 23440 6196
rect 23572 6248 23624 6254
rect 23572 6190 23624 6196
rect 23400 5681 23428 6190
rect 23480 6180 23532 6186
rect 23480 6122 23532 6128
rect 23386 5672 23442 5681
rect 23386 5607 23442 5616
rect 23400 5234 23428 5607
rect 23492 5370 23520 6122
rect 23584 5574 23612 6190
rect 23572 5568 23624 5574
rect 23572 5510 23624 5516
rect 23480 5364 23532 5370
rect 23480 5306 23532 5312
rect 23388 5228 23440 5234
rect 23388 5170 23440 5176
rect 23572 5228 23624 5234
rect 23572 5170 23624 5176
rect 23296 5024 23348 5030
rect 23296 4966 23348 4972
rect 23584 4826 23612 5170
rect 23572 4820 23624 4826
rect 23572 4762 23624 4768
rect 23676 4706 23704 9250
rect 23848 9104 23900 9110
rect 23848 9046 23900 9052
rect 23860 8922 23888 9046
rect 23768 8894 23888 8922
rect 23768 8566 23796 8894
rect 23848 8832 23900 8838
rect 23848 8774 23900 8780
rect 23756 8560 23808 8566
rect 23756 8502 23808 8508
rect 23860 8294 23888 8774
rect 23848 8288 23900 8294
rect 23768 8248 23848 8276
rect 23768 6186 23796 8248
rect 23848 8230 23900 8236
rect 23952 7721 23980 11194
rect 24124 9852 24176 9858
rect 24124 9794 24176 9800
rect 24136 9722 24164 9794
rect 24124 9716 24176 9722
rect 24124 9658 24176 9664
rect 24032 8968 24084 8974
rect 24032 8910 24084 8916
rect 23938 7712 23994 7721
rect 23938 7647 23994 7656
rect 23848 6928 23900 6934
rect 23848 6870 23900 6876
rect 23756 6180 23808 6186
rect 23756 6122 23808 6128
rect 23756 5636 23808 5642
rect 23756 5578 23808 5584
rect 23768 5234 23796 5578
rect 23756 5228 23808 5234
rect 23756 5170 23808 5176
rect 23768 4758 23796 5170
rect 23400 4678 23704 4706
rect 23756 4752 23808 4758
rect 23756 4694 23808 4700
rect 23296 4548 23348 4554
rect 23296 4490 23348 4496
rect 23124 4282 23244 4298
rect 23112 4276 23244 4282
rect 23164 4270 23244 4276
rect 23112 4218 23164 4224
rect 23020 4208 23072 4214
rect 23020 4150 23072 4156
rect 22928 3936 22980 3942
rect 22928 3878 22980 3884
rect 23032 3738 23060 4150
rect 23308 4146 23336 4490
rect 23296 4140 23348 4146
rect 23296 4082 23348 4088
rect 23112 4072 23164 4078
rect 23112 4014 23164 4020
rect 23124 3738 23152 4014
rect 23020 3732 23072 3738
rect 23020 3674 23072 3680
rect 23112 3732 23164 3738
rect 23112 3674 23164 3680
rect 23400 3058 23428 4678
rect 23572 4616 23624 4622
rect 23572 4558 23624 4564
rect 23584 4457 23612 4558
rect 23570 4448 23626 4457
rect 23570 4383 23626 4392
rect 23756 4140 23808 4146
rect 23756 4082 23808 4088
rect 23664 3936 23716 3942
rect 23768 3924 23796 4082
rect 23716 3896 23796 3924
rect 23664 3878 23716 3884
rect 23480 3528 23532 3534
rect 23480 3470 23532 3476
rect 23388 3052 23440 3058
rect 23388 2994 23440 3000
rect 23204 2848 23256 2854
rect 23204 2790 23256 2796
rect 22848 2746 22968 2774
rect 22940 2650 22968 2746
rect 22928 2644 22980 2650
rect 22928 2586 22980 2592
rect 21640 2508 21692 2514
rect 21640 2450 21692 2456
rect 23216 2446 23244 2790
rect 23204 2440 23256 2446
rect 23204 2382 23256 2388
rect 21088 2304 21140 2310
rect 21088 2246 21140 2252
rect 21548 2304 21600 2310
rect 21548 2246 21600 2252
rect 21010 2204 21318 2213
rect 21010 2202 21016 2204
rect 21072 2202 21096 2204
rect 21152 2202 21176 2204
rect 21232 2202 21256 2204
rect 21312 2202 21318 2204
rect 21072 2150 21074 2202
rect 21254 2150 21256 2202
rect 21010 2148 21016 2150
rect 21072 2148 21096 2150
rect 21152 2148 21176 2150
rect 21232 2148 21256 2150
rect 21312 2148 21318 2150
rect 21010 2139 21318 2148
rect 20916 1142 21036 1170
rect 21008 56 21036 1142
rect 23492 882 23520 3470
rect 23860 3194 23888 6870
rect 23940 6656 23992 6662
rect 23940 6598 23992 6604
rect 23952 5642 23980 6598
rect 24044 5846 24072 8910
rect 24124 8628 24176 8634
rect 24124 8570 24176 8576
rect 24136 8265 24164 8570
rect 24122 8256 24178 8265
rect 24122 8191 24178 8200
rect 24228 8004 24256 11194
rect 24504 10033 24532 11194
rect 24490 10024 24546 10033
rect 24490 9959 24546 9968
rect 24400 9512 24452 9518
rect 24400 9454 24452 9460
rect 24308 9036 24360 9042
rect 24308 8978 24360 8984
rect 24320 8430 24348 8978
rect 24308 8424 24360 8430
rect 24308 8366 24360 8372
rect 24228 7976 24348 8004
rect 24124 7880 24176 7886
rect 24124 7822 24176 7828
rect 24136 7410 24164 7822
rect 24214 7576 24270 7585
rect 24214 7511 24270 7520
rect 24124 7404 24176 7410
rect 24124 7346 24176 7352
rect 24124 7268 24176 7274
rect 24124 7210 24176 7216
rect 24136 7177 24164 7210
rect 24122 7168 24178 7177
rect 24122 7103 24178 7112
rect 24124 6724 24176 6730
rect 24124 6666 24176 6672
rect 24136 6089 24164 6666
rect 24122 6080 24178 6089
rect 24122 6015 24178 6024
rect 24228 5846 24256 7511
rect 24320 6769 24348 7976
rect 24306 6760 24362 6769
rect 24306 6695 24362 6704
rect 24032 5840 24084 5846
rect 24032 5782 24084 5788
rect 24216 5840 24268 5846
rect 24216 5782 24268 5788
rect 24412 5794 24440 9454
rect 24492 8560 24544 8566
rect 24490 8528 24492 8537
rect 24584 8560 24636 8566
rect 24544 8528 24546 8537
rect 24584 8502 24636 8508
rect 24490 8463 24546 8472
rect 24596 7954 24624 8502
rect 24676 8424 24728 8430
rect 24676 8366 24728 8372
rect 24688 8294 24716 8366
rect 24780 8294 24808 11194
rect 24860 8356 24912 8362
rect 24860 8298 24912 8304
rect 24676 8288 24728 8294
rect 24676 8230 24728 8236
rect 24768 8288 24820 8294
rect 24768 8230 24820 8236
rect 24584 7948 24636 7954
rect 24584 7890 24636 7896
rect 24492 7812 24544 7818
rect 24492 7754 24544 7760
rect 24504 5914 24532 7754
rect 24676 6792 24728 6798
rect 24676 6734 24728 6740
rect 24768 6792 24820 6798
rect 24768 6734 24820 6740
rect 24688 6322 24716 6734
rect 24780 6662 24808 6734
rect 24872 6662 24900 8298
rect 25056 8090 25084 11194
rect 25134 9752 25190 9761
rect 25134 9687 25190 9696
rect 25044 8084 25096 8090
rect 25044 8026 25096 8032
rect 25044 7948 25096 7954
rect 25044 7890 25096 7896
rect 24952 7812 25004 7818
rect 24952 7754 25004 7760
rect 24964 7546 24992 7754
rect 24952 7540 25004 7546
rect 24952 7482 25004 7488
rect 24768 6656 24820 6662
rect 24768 6598 24820 6604
rect 24860 6656 24912 6662
rect 24860 6598 24912 6604
rect 25056 6610 25084 7890
rect 25148 6798 25176 9687
rect 25332 8838 25360 11194
rect 25412 9308 25464 9314
rect 25412 9250 25464 9256
rect 25320 8832 25372 8838
rect 25320 8774 25372 8780
rect 25228 8628 25280 8634
rect 25228 8570 25280 8576
rect 25240 8537 25268 8570
rect 25226 8528 25282 8537
rect 25226 8463 25282 8472
rect 25228 8356 25280 8362
rect 25228 8298 25280 8304
rect 25320 8356 25372 8362
rect 25320 8298 25372 8304
rect 25136 6792 25188 6798
rect 25136 6734 25188 6740
rect 25056 6582 25176 6610
rect 25042 6488 25098 6497
rect 25042 6423 25098 6432
rect 24676 6316 24728 6322
rect 24676 6258 24728 6264
rect 25056 6118 25084 6423
rect 24952 6112 25004 6118
rect 24952 6054 25004 6060
rect 25044 6112 25096 6118
rect 25044 6054 25096 6060
rect 24492 5908 24544 5914
rect 24492 5850 24544 5856
rect 24412 5766 24532 5794
rect 24964 5778 24992 6054
rect 24400 5704 24452 5710
rect 24400 5646 24452 5652
rect 23940 5636 23992 5642
rect 23940 5578 23992 5584
rect 24412 5574 24440 5646
rect 24216 5568 24268 5574
rect 24216 5510 24268 5516
rect 24400 5568 24452 5574
rect 24400 5510 24452 5516
rect 23938 4720 23994 4729
rect 23938 4655 23940 4664
rect 23992 4655 23994 4664
rect 23940 4626 23992 4632
rect 23940 3936 23992 3942
rect 23940 3878 23992 3884
rect 23848 3188 23900 3194
rect 23848 3130 23900 3136
rect 23572 2984 23624 2990
rect 23572 2926 23624 2932
rect 23584 2417 23612 2926
rect 23570 2408 23626 2417
rect 23570 2343 23626 2352
rect 23480 876 23532 882
rect 23480 818 23532 824
rect 23952 610 23980 3878
rect 24228 3466 24256 5510
rect 24400 4480 24452 4486
rect 24400 4422 24452 4428
rect 24412 4146 24440 4422
rect 24400 4140 24452 4146
rect 24400 4082 24452 4088
rect 24504 3670 24532 5766
rect 24584 5772 24636 5778
rect 24584 5714 24636 5720
rect 24952 5772 25004 5778
rect 24952 5714 25004 5720
rect 24596 4282 24624 5714
rect 24768 5704 24820 5710
rect 24768 5646 24820 5652
rect 24780 4622 24808 5646
rect 24860 5568 24912 5574
rect 24860 5510 24912 5516
rect 24872 4622 24900 5510
rect 24768 4616 24820 4622
rect 24768 4558 24820 4564
rect 24860 4616 24912 4622
rect 24860 4558 24912 4564
rect 24584 4276 24636 4282
rect 24584 4218 24636 4224
rect 24676 4140 24728 4146
rect 24676 4082 24728 4088
rect 24688 3777 24716 4082
rect 24674 3768 24730 3777
rect 24674 3703 24730 3712
rect 24492 3664 24544 3670
rect 24492 3606 24544 3612
rect 24216 3460 24268 3466
rect 24216 3402 24268 3408
rect 24122 3224 24178 3233
rect 24122 3159 24124 3168
rect 24176 3159 24178 3168
rect 24124 3130 24176 3136
rect 24228 2990 24256 3402
rect 25148 3126 25176 6582
rect 25240 6322 25268 8298
rect 25228 6316 25280 6322
rect 25228 6258 25280 6264
rect 25332 5370 25360 8298
rect 25424 7002 25452 9250
rect 25608 8906 25636 11194
rect 25884 9761 25912 11194
rect 25870 9752 25926 9761
rect 25870 9687 25926 9696
rect 26160 9246 26188 11194
rect 26436 10146 26464 11194
rect 26436 10118 26556 10146
rect 26424 9444 26476 9450
rect 26424 9386 26476 9392
rect 26148 9240 26200 9246
rect 26148 9182 26200 9188
rect 26332 9172 26384 9178
rect 26332 9114 26384 9120
rect 25596 8900 25648 8906
rect 25596 8842 25648 8848
rect 25872 8560 25924 8566
rect 25872 8502 25924 8508
rect 25688 8492 25740 8498
rect 25608 8452 25688 8480
rect 25504 7948 25556 7954
rect 25504 7890 25556 7896
rect 25412 6996 25464 7002
rect 25412 6938 25464 6944
rect 25516 6746 25544 7890
rect 25608 6916 25636 8452
rect 25688 8434 25740 8440
rect 25780 8424 25832 8430
rect 25780 8366 25832 8372
rect 25688 8288 25740 8294
rect 25792 8265 25820 8366
rect 25688 8230 25740 8236
rect 25778 8256 25834 8265
rect 25700 7410 25728 8230
rect 25778 8191 25834 8200
rect 25884 7818 25912 8502
rect 25950 8188 26258 8197
rect 25950 8186 25956 8188
rect 26012 8186 26036 8188
rect 26092 8186 26116 8188
rect 26172 8186 26196 8188
rect 26252 8186 26258 8188
rect 26012 8134 26014 8186
rect 26194 8134 26196 8186
rect 25950 8132 25956 8134
rect 26012 8132 26036 8134
rect 26092 8132 26116 8134
rect 26172 8132 26196 8134
rect 26252 8132 26258 8134
rect 25950 8123 26258 8132
rect 25872 7812 25924 7818
rect 25872 7754 25924 7760
rect 26240 7812 26292 7818
rect 26240 7754 26292 7760
rect 25870 7712 25926 7721
rect 25870 7647 25926 7656
rect 25688 7404 25740 7410
rect 25688 7346 25740 7352
rect 25780 7200 25832 7206
rect 25780 7142 25832 7148
rect 25792 7041 25820 7142
rect 25778 7032 25834 7041
rect 25778 6967 25834 6976
rect 25608 6888 25820 6916
rect 25424 6718 25544 6746
rect 25686 6760 25742 6769
rect 25320 5364 25372 5370
rect 25320 5306 25372 5312
rect 25228 5024 25280 5030
rect 25228 4966 25280 4972
rect 25240 4690 25268 4966
rect 25228 4684 25280 4690
rect 25228 4626 25280 4632
rect 25332 4486 25360 5306
rect 25320 4480 25372 4486
rect 25320 4422 25372 4428
rect 25424 4282 25452 6718
rect 25686 6695 25742 6704
rect 25504 6656 25556 6662
rect 25504 6598 25556 6604
rect 25516 6390 25544 6598
rect 25504 6384 25556 6390
rect 25504 6326 25556 6332
rect 25700 6322 25728 6695
rect 25792 6390 25820 6888
rect 25780 6384 25832 6390
rect 25780 6326 25832 6332
rect 25688 6316 25740 6322
rect 25688 6258 25740 6264
rect 25504 6112 25556 6118
rect 25504 6054 25556 6060
rect 25688 6112 25740 6118
rect 25688 6054 25740 6060
rect 25516 5302 25544 6054
rect 25504 5296 25556 5302
rect 25504 5238 25556 5244
rect 25596 5228 25648 5234
rect 25596 5170 25648 5176
rect 25504 4548 25556 4554
rect 25504 4490 25556 4496
rect 25516 4282 25544 4490
rect 25412 4276 25464 4282
rect 25412 4218 25464 4224
rect 25504 4276 25556 4282
rect 25504 4218 25556 4224
rect 25228 4072 25280 4078
rect 25228 4014 25280 4020
rect 25320 4072 25372 4078
rect 25320 4014 25372 4020
rect 25240 3194 25268 4014
rect 25332 3466 25360 4014
rect 25424 3670 25452 4218
rect 25504 3936 25556 3942
rect 25504 3878 25556 3884
rect 25412 3664 25464 3670
rect 25412 3606 25464 3612
rect 25320 3460 25372 3466
rect 25320 3402 25372 3408
rect 25412 3460 25464 3466
rect 25412 3402 25464 3408
rect 25332 3369 25360 3402
rect 25318 3360 25374 3369
rect 25318 3295 25374 3304
rect 25228 3188 25280 3194
rect 25228 3130 25280 3136
rect 25136 3120 25188 3126
rect 25136 3062 25188 3068
rect 24216 2984 24268 2990
rect 24216 2926 24268 2932
rect 23940 604 23992 610
rect 23940 546 23992 552
rect 23204 196 23256 202
rect 23204 138 23256 144
rect 24308 196 24360 202
rect 24308 138 24360 144
rect 22112 66 22232 82
rect 22112 60 22244 66
rect 22112 56 22192 60
rect 12268 14 12480 42
rect 13266 0 13322 56
rect 14370 0 14426 56
rect 15474 0 15530 56
rect 16578 0 16634 56
rect 17682 0 17738 56
rect 18786 0 18842 56
rect 19890 0 19946 56
rect 20994 0 21050 56
rect 22098 54 22192 56
rect 22098 0 22154 54
rect 23216 56 23244 138
rect 24320 56 24348 138
rect 25424 56 25452 3402
rect 25516 3058 25544 3878
rect 25608 3584 25636 5170
rect 25700 5166 25728 6054
rect 25792 5216 25820 6326
rect 25884 6322 25912 7647
rect 26252 7478 26280 7754
rect 26240 7472 26292 7478
rect 26240 7414 26292 7420
rect 25950 7100 26258 7109
rect 25950 7098 25956 7100
rect 26012 7098 26036 7100
rect 26092 7098 26116 7100
rect 26172 7098 26196 7100
rect 26252 7098 26258 7100
rect 26012 7046 26014 7098
rect 26194 7046 26196 7098
rect 25950 7044 25956 7046
rect 26012 7044 26036 7046
rect 26092 7044 26116 7046
rect 26172 7044 26196 7046
rect 26252 7044 26258 7046
rect 25950 7035 26258 7044
rect 26240 6792 26292 6798
rect 26238 6760 26240 6769
rect 26292 6760 26294 6769
rect 25964 6724 26016 6730
rect 26238 6695 26294 6704
rect 25964 6666 26016 6672
rect 25976 6458 26004 6666
rect 25964 6452 26016 6458
rect 25964 6394 26016 6400
rect 26252 6322 26280 6695
rect 25872 6316 25924 6322
rect 25872 6258 25924 6264
rect 26240 6316 26292 6322
rect 26240 6258 26292 6264
rect 25872 6112 25924 6118
rect 26344 6089 26372 9114
rect 26436 7342 26464 9386
rect 26528 8974 26556 10118
rect 26608 10056 26660 10062
rect 26608 9998 26660 10004
rect 26516 8968 26568 8974
rect 26516 8910 26568 8916
rect 26514 8664 26570 8673
rect 26514 8599 26570 8608
rect 26528 7546 26556 8599
rect 26516 7540 26568 7546
rect 26516 7482 26568 7488
rect 26424 7336 26476 7342
rect 26424 7278 26476 7284
rect 26422 7168 26478 7177
rect 26422 7103 26478 7112
rect 26436 6458 26464 7103
rect 26424 6452 26476 6458
rect 26424 6394 26476 6400
rect 25872 6054 25924 6060
rect 26330 6080 26386 6089
rect 25884 5710 25912 6054
rect 26528 6066 26556 7482
rect 26620 6440 26648 9998
rect 26712 7002 26740 11194
rect 26988 10305 27016 11194
rect 26974 10296 27030 10305
rect 26974 10231 27030 10240
rect 26792 9920 26844 9926
rect 26792 9862 26844 9868
rect 27264 9874 27292 11194
rect 27434 10568 27490 10577
rect 27434 10503 27490 10512
rect 26804 8537 26832 9862
rect 27264 9846 27384 9874
rect 27356 9450 27384 9846
rect 27344 9444 27396 9450
rect 27344 9386 27396 9392
rect 26884 8900 26936 8906
rect 26884 8842 26936 8848
rect 26790 8528 26846 8537
rect 26790 8463 26846 8472
rect 26896 8430 26924 8842
rect 27010 8732 27318 8741
rect 27010 8730 27016 8732
rect 27072 8730 27096 8732
rect 27152 8730 27176 8732
rect 27232 8730 27256 8732
rect 27312 8730 27318 8732
rect 27072 8678 27074 8730
rect 27254 8678 27256 8730
rect 27010 8676 27016 8678
rect 27072 8676 27096 8678
rect 27152 8676 27176 8678
rect 27232 8676 27256 8678
rect 27312 8676 27318 8678
rect 27010 8667 27318 8676
rect 27068 8492 27120 8498
rect 27068 8434 27120 8440
rect 26884 8424 26936 8430
rect 26884 8366 26936 8372
rect 26792 8288 26844 8294
rect 26792 8230 26844 8236
rect 26804 7410 26832 8230
rect 27080 7886 27108 8434
rect 27252 8424 27304 8430
rect 27252 8366 27304 8372
rect 27264 8276 27292 8366
rect 27264 8248 27384 8276
rect 27068 7880 27120 7886
rect 27068 7822 27120 7828
rect 27010 7644 27318 7653
rect 27010 7642 27016 7644
rect 27072 7642 27096 7644
rect 27152 7642 27176 7644
rect 27232 7642 27256 7644
rect 27312 7642 27318 7644
rect 27072 7590 27074 7642
rect 27254 7590 27256 7642
rect 27010 7588 27016 7590
rect 27072 7588 27096 7590
rect 27152 7588 27176 7590
rect 27232 7588 27256 7590
rect 27312 7588 27318 7590
rect 27010 7579 27318 7588
rect 26792 7404 26844 7410
rect 26792 7346 26844 7352
rect 27068 7200 27120 7206
rect 27068 7142 27120 7148
rect 26882 7032 26938 7041
rect 26700 6996 26752 7002
rect 26882 6967 26938 6976
rect 26700 6938 26752 6944
rect 26896 6934 26924 6967
rect 26884 6928 26936 6934
rect 26884 6870 26936 6876
rect 27080 6798 27108 7142
rect 27158 7032 27214 7041
rect 27158 6967 27214 6976
rect 27068 6792 27120 6798
rect 27172 6769 27200 6967
rect 27356 6798 27384 8248
rect 27448 7041 27476 10503
rect 27540 8906 27568 11194
rect 27618 9752 27674 9761
rect 27816 9722 27844 11194
rect 27988 9988 28040 9994
rect 27988 9930 28040 9936
rect 27618 9687 27674 9696
rect 27804 9716 27856 9722
rect 27528 8900 27580 8906
rect 27528 8842 27580 8848
rect 27528 7880 27580 7886
rect 27528 7822 27580 7828
rect 27540 7478 27568 7822
rect 27528 7472 27580 7478
rect 27528 7414 27580 7420
rect 27434 7032 27490 7041
rect 27434 6967 27490 6976
rect 27540 6866 27568 7414
rect 27528 6860 27580 6866
rect 27528 6802 27580 6808
rect 27632 6798 27660 9687
rect 27804 9658 27856 9664
rect 27710 9208 27766 9217
rect 27710 9143 27766 9152
rect 27804 9172 27856 9178
rect 27724 8401 27752 9143
rect 27804 9114 27856 9120
rect 27710 8392 27766 8401
rect 27710 8327 27766 8336
rect 27712 8288 27764 8294
rect 27710 8256 27712 8265
rect 27764 8256 27766 8265
rect 27710 8191 27766 8200
rect 27816 8129 27844 9114
rect 27896 9104 27948 9110
rect 27896 9046 27948 9052
rect 27802 8120 27858 8129
rect 27802 8055 27858 8064
rect 27804 8016 27856 8022
rect 27804 7958 27856 7964
rect 27344 6792 27396 6798
rect 27068 6734 27120 6740
rect 27158 6760 27214 6769
rect 26700 6724 26752 6730
rect 26752 6684 26832 6712
rect 27344 6734 27396 6740
rect 27620 6792 27672 6798
rect 27620 6734 27672 6740
rect 27158 6695 27214 6704
rect 27712 6724 27764 6730
rect 26700 6666 26752 6672
rect 26804 6644 26832 6684
rect 27712 6666 27764 6672
rect 26884 6656 26936 6662
rect 26804 6616 26884 6644
rect 26884 6598 26936 6604
rect 27344 6656 27396 6662
rect 27344 6598 27396 6604
rect 27010 6556 27318 6565
rect 27010 6554 27016 6556
rect 27072 6554 27096 6556
rect 27152 6554 27176 6556
rect 27232 6554 27256 6556
rect 27312 6554 27318 6556
rect 27072 6502 27074 6554
rect 27254 6502 27256 6554
rect 27010 6500 27016 6502
rect 27072 6500 27096 6502
rect 27152 6500 27176 6502
rect 27232 6500 27256 6502
rect 27312 6500 27318 6502
rect 27010 6491 27318 6500
rect 26792 6452 26844 6458
rect 26620 6412 26740 6440
rect 26606 6352 26662 6361
rect 26606 6287 26608 6296
rect 26660 6287 26662 6296
rect 26608 6258 26660 6264
rect 25950 6012 26258 6021
rect 26330 6015 26386 6024
rect 26436 6038 26556 6066
rect 25950 6010 25956 6012
rect 26012 6010 26036 6012
rect 26092 6010 26116 6012
rect 26172 6010 26196 6012
rect 26252 6010 26258 6012
rect 26012 5958 26014 6010
rect 26194 5958 26196 6010
rect 25950 5956 25956 5958
rect 26012 5956 26036 5958
rect 26092 5956 26116 5958
rect 26172 5956 26196 5958
rect 26252 5956 26258 5958
rect 25950 5947 26258 5956
rect 26344 5710 26372 6015
rect 25872 5704 25924 5710
rect 25872 5646 25924 5652
rect 26332 5704 26384 5710
rect 26332 5646 26384 5652
rect 26436 5574 26464 6038
rect 26516 5908 26568 5914
rect 26516 5850 26568 5856
rect 26424 5568 26476 5574
rect 26424 5510 26476 5516
rect 26332 5296 26384 5302
rect 26332 5238 26384 5244
rect 26424 5296 26476 5302
rect 26424 5238 26476 5244
rect 25964 5228 26016 5234
rect 25792 5188 25964 5216
rect 25688 5160 25740 5166
rect 25688 5102 25740 5108
rect 25792 4049 25820 5188
rect 25964 5170 26016 5176
rect 25950 4924 26258 4933
rect 25950 4922 25956 4924
rect 26012 4922 26036 4924
rect 26092 4922 26116 4924
rect 26172 4922 26196 4924
rect 26252 4922 26258 4924
rect 26012 4870 26014 4922
rect 26194 4870 26196 4922
rect 25950 4868 25956 4870
rect 26012 4868 26036 4870
rect 26092 4868 26116 4870
rect 26172 4868 26196 4870
rect 26252 4868 26258 4870
rect 25950 4859 26258 4868
rect 26240 4616 26292 4622
rect 26344 4604 26372 5238
rect 26292 4576 26372 4604
rect 26240 4558 26292 4564
rect 26252 4214 26280 4558
rect 26436 4321 26464 5238
rect 26422 4312 26478 4321
rect 26422 4247 26478 4256
rect 26240 4208 26292 4214
rect 26240 4150 26292 4156
rect 26332 4072 26384 4078
rect 25778 4040 25834 4049
rect 26528 4049 26556 5850
rect 26606 5536 26662 5545
rect 26606 5471 26662 5480
rect 26620 4622 26648 5471
rect 26712 5370 26740 6412
rect 26976 6452 27028 6458
rect 26844 6412 26924 6440
rect 26792 6394 26844 6400
rect 26790 6352 26846 6361
rect 26790 6287 26846 6296
rect 26700 5364 26752 5370
rect 26700 5306 26752 5312
rect 26804 5166 26832 6287
rect 26792 5160 26844 5166
rect 26792 5102 26844 5108
rect 26700 5024 26752 5030
rect 26792 5024 26844 5030
rect 26700 4966 26752 4972
rect 26790 4992 26792 5001
rect 26844 4992 26846 5001
rect 26608 4616 26660 4622
rect 26608 4558 26660 4564
rect 26606 4448 26662 4457
rect 26606 4383 26662 4392
rect 26332 4014 26384 4020
rect 26514 4040 26570 4049
rect 25778 3975 25834 3984
rect 25950 3836 26258 3845
rect 25950 3834 25956 3836
rect 26012 3834 26036 3836
rect 26092 3834 26116 3836
rect 26172 3834 26196 3836
rect 26252 3834 26258 3836
rect 26012 3782 26014 3834
rect 26194 3782 26196 3834
rect 25950 3780 25956 3782
rect 26012 3780 26036 3782
rect 26092 3780 26116 3782
rect 26172 3780 26196 3782
rect 26252 3780 26258 3782
rect 25950 3771 26258 3780
rect 25964 3664 26016 3670
rect 25964 3606 26016 3612
rect 26146 3632 26202 3641
rect 25780 3596 25832 3602
rect 25608 3556 25780 3584
rect 25780 3538 25832 3544
rect 25792 3194 25820 3538
rect 25976 3534 26004 3606
rect 26146 3567 26202 3576
rect 25964 3528 26016 3534
rect 25964 3470 26016 3476
rect 26160 3466 26188 3567
rect 26148 3460 26200 3466
rect 26148 3402 26200 3408
rect 25780 3188 25832 3194
rect 25780 3130 25832 3136
rect 26160 3126 26188 3402
rect 26148 3120 26200 3126
rect 26148 3062 26200 3068
rect 26344 3058 26372 4014
rect 26514 3975 26570 3984
rect 26620 3913 26648 4383
rect 26712 4010 26740 4966
rect 26790 4927 26846 4936
rect 26792 4208 26844 4214
rect 26792 4150 26844 4156
rect 26700 4004 26752 4010
rect 26700 3946 26752 3952
rect 26606 3904 26662 3913
rect 26606 3839 26662 3848
rect 26514 3768 26570 3777
rect 26514 3703 26570 3712
rect 26422 3632 26478 3641
rect 26528 3602 26556 3703
rect 26804 3602 26832 4150
rect 26422 3567 26478 3576
rect 26516 3596 26568 3602
rect 26436 3369 26464 3567
rect 26516 3538 26568 3544
rect 26792 3596 26844 3602
rect 26792 3538 26844 3544
rect 26422 3360 26478 3369
rect 26422 3295 26478 3304
rect 25504 3052 25556 3058
rect 25504 2994 25556 3000
rect 25780 3052 25832 3058
rect 25780 2994 25832 3000
rect 26332 3052 26384 3058
rect 26332 2994 26384 3000
rect 26792 3052 26844 3058
rect 26792 2994 26844 3000
rect 25792 2825 25820 2994
rect 25962 2952 26018 2961
rect 25962 2887 26018 2896
rect 26606 2952 26662 2961
rect 26606 2887 26662 2896
rect 25976 2854 26004 2887
rect 26620 2854 26648 2887
rect 25964 2848 26016 2854
rect 25778 2816 25834 2825
rect 25964 2790 26016 2796
rect 26608 2848 26660 2854
rect 26608 2790 26660 2796
rect 25778 2751 25834 2760
rect 25950 2748 26258 2757
rect 25950 2746 25956 2748
rect 26012 2746 26036 2748
rect 26092 2746 26116 2748
rect 26172 2746 26196 2748
rect 26252 2746 26258 2748
rect 26012 2694 26014 2746
rect 26194 2694 26196 2746
rect 25950 2692 25956 2694
rect 26012 2692 26036 2694
rect 26092 2692 26116 2694
rect 26172 2692 26196 2694
rect 26252 2692 26258 2694
rect 25950 2683 26258 2692
rect 26804 2650 26832 2994
rect 26896 2774 26924 6412
rect 26976 6394 27028 6400
rect 26988 6118 27016 6394
rect 26976 6112 27028 6118
rect 26976 6054 27028 6060
rect 27160 6112 27212 6118
rect 27160 6054 27212 6060
rect 27172 5914 27200 6054
rect 27160 5908 27212 5914
rect 27160 5850 27212 5856
rect 27356 5817 27384 6598
rect 27528 6452 27580 6458
rect 27528 6394 27580 6400
rect 27540 6254 27568 6394
rect 27618 6352 27674 6361
rect 27618 6287 27620 6296
rect 27672 6287 27674 6296
rect 27620 6258 27672 6264
rect 27528 6248 27580 6254
rect 27528 6190 27580 6196
rect 27342 5808 27398 5817
rect 27342 5743 27398 5752
rect 27436 5772 27488 5778
rect 27436 5714 27488 5720
rect 27344 5568 27396 5574
rect 27344 5510 27396 5516
rect 27010 5468 27318 5477
rect 27010 5466 27016 5468
rect 27072 5466 27096 5468
rect 27152 5466 27176 5468
rect 27232 5466 27256 5468
rect 27312 5466 27318 5468
rect 27072 5414 27074 5466
rect 27254 5414 27256 5466
rect 27010 5412 27016 5414
rect 27072 5412 27096 5414
rect 27152 5412 27176 5414
rect 27232 5412 27256 5414
rect 27312 5412 27318 5414
rect 27010 5403 27318 5412
rect 27160 5364 27212 5370
rect 27160 5306 27212 5312
rect 27068 5160 27120 5166
rect 27068 5102 27120 5108
rect 27080 4758 27108 5102
rect 27172 4826 27200 5306
rect 27356 5234 27384 5510
rect 27448 5370 27476 5714
rect 27436 5364 27488 5370
rect 27436 5306 27488 5312
rect 27344 5228 27396 5234
rect 27344 5170 27396 5176
rect 27540 5114 27568 6190
rect 27620 5568 27672 5574
rect 27620 5510 27672 5516
rect 27632 5234 27660 5510
rect 27620 5228 27672 5234
rect 27620 5170 27672 5176
rect 27356 5086 27568 5114
rect 27160 4820 27212 4826
rect 27160 4762 27212 4768
rect 27068 4752 27120 4758
rect 27068 4694 27120 4700
rect 26976 4684 27028 4690
rect 26976 4626 27028 4632
rect 26988 4554 27016 4626
rect 26976 4548 27028 4554
rect 26976 4490 27028 4496
rect 27010 4380 27318 4389
rect 27010 4378 27016 4380
rect 27072 4378 27096 4380
rect 27152 4378 27176 4380
rect 27232 4378 27256 4380
rect 27312 4378 27318 4380
rect 27072 4326 27074 4378
rect 27254 4326 27256 4378
rect 27010 4324 27016 4326
rect 27072 4324 27096 4326
rect 27152 4324 27176 4326
rect 27232 4324 27256 4326
rect 27312 4324 27318 4326
rect 27010 4315 27318 4324
rect 27356 4078 27384 5086
rect 27436 5024 27488 5030
rect 27436 4966 27488 4972
rect 27528 5024 27580 5030
rect 27528 4966 27580 4972
rect 27448 4622 27476 4966
rect 27436 4616 27488 4622
rect 27436 4558 27488 4564
rect 27344 4072 27396 4078
rect 27344 4014 27396 4020
rect 27344 3936 27396 3942
rect 27344 3878 27396 3884
rect 27010 3292 27318 3301
rect 27010 3290 27016 3292
rect 27072 3290 27096 3292
rect 27152 3290 27176 3292
rect 27232 3290 27256 3292
rect 27312 3290 27318 3292
rect 27072 3238 27074 3290
rect 27254 3238 27256 3290
rect 27010 3236 27016 3238
rect 27072 3236 27096 3238
rect 27152 3236 27176 3238
rect 27232 3236 27256 3238
rect 27312 3236 27318 3238
rect 27010 3227 27318 3236
rect 27252 2848 27304 2854
rect 27250 2816 27252 2825
rect 27304 2816 27306 2825
rect 26896 2746 27108 2774
rect 27250 2751 27306 2760
rect 26792 2644 26844 2650
rect 26792 2586 26844 2592
rect 26884 2508 26936 2514
rect 26804 2468 26884 2496
rect 25872 2304 25924 2310
rect 25872 2246 25924 2252
rect 25884 1630 25912 2246
rect 26804 2106 26832 2468
rect 26884 2450 26936 2456
rect 27080 2394 27108 2746
rect 26896 2366 27108 2394
rect 26792 2100 26844 2106
rect 26792 2042 26844 2048
rect 26896 2038 26924 2366
rect 27010 2204 27318 2213
rect 27010 2202 27016 2204
rect 27072 2202 27096 2204
rect 27152 2202 27176 2204
rect 27232 2202 27256 2204
rect 27312 2202 27318 2204
rect 27072 2150 27074 2202
rect 27254 2150 27256 2202
rect 27010 2148 27016 2150
rect 27072 2148 27096 2150
rect 27152 2148 27176 2150
rect 27232 2148 27256 2150
rect 27312 2148 27318 2150
rect 27010 2139 27318 2148
rect 26884 2032 26936 2038
rect 26514 2000 26570 2009
rect 26884 1974 26936 1980
rect 26514 1935 26570 1944
rect 25872 1624 25924 1630
rect 25872 1566 25924 1572
rect 26528 56 26556 1935
rect 27356 1601 27384 3878
rect 27540 3738 27568 4966
rect 27620 4752 27672 4758
rect 27620 4694 27672 4700
rect 27632 4146 27660 4694
rect 27620 4140 27672 4146
rect 27620 4082 27672 4088
rect 27528 3732 27580 3738
rect 27528 3674 27580 3680
rect 27724 3602 27752 6666
rect 27712 3596 27764 3602
rect 27712 3538 27764 3544
rect 27434 3224 27490 3233
rect 27434 3159 27490 3168
rect 27448 2394 27476 3159
rect 27618 2952 27674 2961
rect 27618 2887 27674 2896
rect 27526 2816 27582 2825
rect 27526 2751 27582 2760
rect 27540 2514 27568 2751
rect 27528 2508 27580 2514
rect 27528 2450 27580 2456
rect 27448 2366 27568 2394
rect 27342 1592 27398 1601
rect 27342 1527 27398 1536
rect 27540 746 27568 2366
rect 27528 740 27580 746
rect 27528 682 27580 688
rect 27632 56 27660 2887
rect 27816 2446 27844 7958
rect 27908 5914 27936 9046
rect 28000 7750 28028 9930
rect 28092 8673 28120 11194
rect 28368 10282 28396 11194
rect 28368 10254 28580 10282
rect 28446 10160 28502 10169
rect 28446 10095 28502 10104
rect 28354 10024 28410 10033
rect 28354 9959 28410 9968
rect 28170 9888 28226 9897
rect 28170 9823 28226 9832
rect 28078 8664 28134 8673
rect 28078 8599 28134 8608
rect 28080 8560 28132 8566
rect 28184 8548 28212 9823
rect 28262 8664 28318 8673
rect 28262 8599 28264 8608
rect 28316 8599 28318 8608
rect 28264 8570 28316 8576
rect 28132 8520 28212 8548
rect 28080 8502 28132 8508
rect 28264 8492 28316 8498
rect 28184 8452 28264 8480
rect 28184 8265 28212 8452
rect 28264 8434 28316 8440
rect 28264 8356 28316 8362
rect 28264 8298 28316 8304
rect 28170 8256 28226 8265
rect 28170 8191 28226 8200
rect 27988 7744 28040 7750
rect 27988 7686 28040 7692
rect 28276 6798 28304 8298
rect 28368 7886 28396 9959
rect 28460 7886 28488 10095
rect 28356 7880 28408 7886
rect 28356 7822 28408 7828
rect 28448 7880 28500 7886
rect 28448 7822 28500 7828
rect 28552 7721 28580 10254
rect 28538 7712 28594 7721
rect 28538 7647 28594 7656
rect 28540 7404 28592 7410
rect 28540 7346 28592 7352
rect 28552 7177 28580 7346
rect 28538 7168 28594 7177
rect 28538 7103 28594 7112
rect 28264 6792 28316 6798
rect 28264 6734 28316 6740
rect 28644 6730 28672 11194
rect 28920 10334 28948 11194
rect 28908 10328 28960 10334
rect 28908 10270 28960 10276
rect 29000 9444 29052 9450
rect 29000 9386 29052 9392
rect 28816 9240 28868 9246
rect 28816 9182 28868 9188
rect 28724 8288 28776 8294
rect 28724 8230 28776 8236
rect 28736 8129 28764 8230
rect 28722 8120 28778 8129
rect 28722 8055 28778 8064
rect 28724 8016 28776 8022
rect 28722 7984 28724 7993
rect 28776 7984 28778 7993
rect 28722 7919 28778 7928
rect 28828 7818 28856 9182
rect 28906 8664 28962 8673
rect 29012 8634 29040 9386
rect 29090 8664 29146 8673
rect 28906 8599 28908 8608
rect 28960 8599 28962 8608
rect 29000 8628 29052 8634
rect 28908 8570 28960 8576
rect 29090 8599 29146 8608
rect 29000 8570 29052 8576
rect 29104 8498 29132 8599
rect 29000 8492 29052 8498
rect 29000 8434 29052 8440
rect 29092 8492 29144 8498
rect 29196 8480 29224 11194
rect 29472 10418 29500 11194
rect 29472 10390 29684 10418
rect 29458 10296 29514 10305
rect 29458 10231 29514 10240
rect 29368 9104 29420 9110
rect 29368 9046 29420 9052
rect 29196 8452 29316 8480
rect 29092 8434 29144 8440
rect 28908 8356 28960 8362
rect 28908 8298 28960 8304
rect 28920 8265 28948 8298
rect 28906 8256 28962 8265
rect 28906 8191 28962 8200
rect 28908 8084 28960 8090
rect 28908 8026 28960 8032
rect 28920 7886 28948 8026
rect 28908 7880 28960 7886
rect 28908 7822 28960 7828
rect 28816 7812 28868 7818
rect 28816 7754 28868 7760
rect 29012 7546 29040 8434
rect 29092 8356 29144 8362
rect 29092 8298 29144 8304
rect 29000 7540 29052 7546
rect 29000 7482 29052 7488
rect 29104 6866 29132 8298
rect 29184 8016 29236 8022
rect 29184 7958 29236 7964
rect 29196 7041 29224 7958
rect 29182 7032 29238 7041
rect 29182 6967 29238 6976
rect 29092 6860 29144 6866
rect 29092 6802 29144 6808
rect 28632 6724 28684 6730
rect 28632 6666 28684 6672
rect 29000 6656 29052 6662
rect 29000 6598 29052 6604
rect 27986 6488 28042 6497
rect 27986 6423 28042 6432
rect 27896 5908 27948 5914
rect 27896 5850 27948 5856
rect 27896 5092 27948 5098
rect 27896 5034 27948 5040
rect 27908 5001 27936 5034
rect 27894 4992 27950 5001
rect 27894 4927 27950 4936
rect 28000 4298 28028 6423
rect 28814 6352 28870 6361
rect 28724 6316 28776 6322
rect 28814 6287 28870 6296
rect 28724 6258 28776 6264
rect 28632 6112 28684 6118
rect 28736 6089 28764 6258
rect 28632 6054 28684 6060
rect 28722 6080 28778 6089
rect 28264 5908 28316 5914
rect 28184 5868 28264 5896
rect 28080 5840 28132 5846
rect 28080 5782 28132 5788
rect 27908 4270 28028 4298
rect 27908 4214 27936 4270
rect 27896 4208 27948 4214
rect 27988 4208 28040 4214
rect 27896 4150 27948 4156
rect 27986 4176 27988 4185
rect 28040 4176 28042 4185
rect 27986 4111 28042 4120
rect 27804 2440 27856 2446
rect 27804 2382 27856 2388
rect 27712 2100 27764 2106
rect 27712 2042 27764 2048
rect 27724 785 27752 2042
rect 28092 1902 28120 5782
rect 28184 3777 28212 5868
rect 28264 5850 28316 5856
rect 28644 5710 28672 6054
rect 28722 6015 28778 6024
rect 28632 5704 28684 5710
rect 28632 5646 28684 5652
rect 28724 5704 28776 5710
rect 28724 5646 28776 5652
rect 28264 5636 28316 5642
rect 28264 5578 28316 5584
rect 28276 4622 28304 5578
rect 28368 5234 28672 5250
rect 28356 5228 28672 5234
rect 28408 5222 28672 5228
rect 28356 5170 28408 5176
rect 28448 5160 28500 5166
rect 28448 5102 28500 5108
rect 28264 4616 28316 4622
rect 28264 4558 28316 4564
rect 28356 4616 28408 4622
rect 28356 4558 28408 4564
rect 28368 4214 28396 4558
rect 28356 4208 28408 4214
rect 28356 4150 28408 4156
rect 28264 4072 28316 4078
rect 28264 4014 28316 4020
rect 28170 3768 28226 3777
rect 28276 3738 28304 4014
rect 28170 3703 28226 3712
rect 28264 3732 28316 3738
rect 28264 3674 28316 3680
rect 28172 3528 28224 3534
rect 28172 3470 28224 3476
rect 28080 1896 28132 1902
rect 28080 1838 28132 1844
rect 28184 1086 28212 3470
rect 28460 3398 28488 5102
rect 28540 4616 28592 4622
rect 28540 4558 28592 4564
rect 28448 3392 28500 3398
rect 28448 3334 28500 3340
rect 28552 3194 28580 4558
rect 28540 3188 28592 3194
rect 28540 3130 28592 3136
rect 28552 3058 28580 3130
rect 28644 3126 28672 5222
rect 28736 4078 28764 5646
rect 28724 4072 28776 4078
rect 28724 4014 28776 4020
rect 28632 3120 28684 3126
rect 28632 3062 28684 3068
rect 28540 3052 28592 3058
rect 28540 2994 28592 3000
rect 28644 2417 28672 3062
rect 28828 2774 28856 6287
rect 29012 5710 29040 6598
rect 29184 5840 29236 5846
rect 29184 5782 29236 5788
rect 29000 5704 29052 5710
rect 29000 5646 29052 5652
rect 29092 5704 29144 5710
rect 29092 5646 29144 5652
rect 29000 5568 29052 5574
rect 29000 5510 29052 5516
rect 28908 5092 28960 5098
rect 28908 5034 28960 5040
rect 28920 4690 28948 5034
rect 29012 4826 29040 5510
rect 29104 5370 29132 5646
rect 29196 5370 29224 5782
rect 29288 5778 29316 8452
rect 29380 8362 29408 9046
rect 29368 8356 29420 8362
rect 29368 8298 29420 8304
rect 29368 8016 29420 8022
rect 29368 7958 29420 7964
rect 29380 7750 29408 7958
rect 29368 7744 29420 7750
rect 29368 7686 29420 7692
rect 29368 7404 29420 7410
rect 29368 7346 29420 7352
rect 29380 7177 29408 7346
rect 29366 7168 29422 7177
rect 29366 7103 29422 7112
rect 29472 6798 29500 10231
rect 29552 9512 29604 9518
rect 29552 9454 29604 9460
rect 29564 8498 29592 9454
rect 29552 8492 29604 8498
rect 29552 8434 29604 8440
rect 29552 8288 29604 8294
rect 29552 8230 29604 8236
rect 29564 7478 29592 8230
rect 29656 7970 29684 10390
rect 29748 9246 29776 11194
rect 30024 9382 30052 11194
rect 29828 9376 29880 9382
rect 29828 9318 29880 9324
rect 30012 9376 30064 9382
rect 30012 9318 30064 9324
rect 29736 9240 29788 9246
rect 29736 9182 29788 9188
rect 29840 8820 29868 9318
rect 30104 9036 30156 9042
rect 30104 8978 30156 8984
rect 29840 8792 29960 8820
rect 29826 8664 29882 8673
rect 29826 8599 29882 8608
rect 29840 8566 29868 8599
rect 29828 8560 29880 8566
rect 29828 8502 29880 8508
rect 29736 8288 29788 8294
rect 29736 8230 29788 8236
rect 29748 8090 29776 8230
rect 29840 8090 29868 8502
rect 29932 8294 29960 8792
rect 30116 8566 30144 8978
rect 30196 8832 30248 8838
rect 30196 8774 30248 8780
rect 30104 8560 30156 8566
rect 30104 8502 30156 8508
rect 30208 8498 30236 8774
rect 30196 8492 30248 8498
rect 30196 8434 30248 8440
rect 30012 8424 30064 8430
rect 30012 8366 30064 8372
rect 29920 8288 29972 8294
rect 29920 8230 29972 8236
rect 29736 8084 29788 8090
rect 29736 8026 29788 8032
rect 29828 8084 29880 8090
rect 29828 8026 29880 8032
rect 29656 7942 29776 7970
rect 29644 7880 29696 7886
rect 29644 7822 29696 7828
rect 29552 7472 29604 7478
rect 29552 7414 29604 7420
rect 29656 7410 29684 7822
rect 29748 7585 29776 7942
rect 29734 7576 29790 7585
rect 30024 7546 30052 8366
rect 30196 8084 30248 8090
rect 30196 8026 30248 8032
rect 29734 7511 29790 7520
rect 30012 7540 30064 7546
rect 30012 7482 30064 7488
rect 29828 7472 29880 7478
rect 29828 7414 29880 7420
rect 29644 7404 29696 7410
rect 29644 7346 29696 7352
rect 29736 7336 29788 7342
rect 29736 7278 29788 7284
rect 29460 6792 29512 6798
rect 29460 6734 29512 6740
rect 29642 6760 29698 6769
rect 29642 6695 29698 6704
rect 29656 6662 29684 6695
rect 29644 6656 29696 6662
rect 29644 6598 29696 6604
rect 29748 6458 29776 7278
rect 29840 6798 29868 7414
rect 30104 7404 30156 7410
rect 30104 7346 30156 7352
rect 30116 7002 30144 7346
rect 30104 6996 30156 7002
rect 30104 6938 30156 6944
rect 30208 6798 30236 8026
rect 30300 7993 30328 11194
rect 30472 10192 30524 10198
rect 30472 10134 30524 10140
rect 30380 8492 30432 8498
rect 30380 8434 30432 8440
rect 30286 7984 30342 7993
rect 30286 7919 30342 7928
rect 30286 7712 30342 7721
rect 30286 7647 30342 7656
rect 29828 6792 29880 6798
rect 29828 6734 29880 6740
rect 30196 6792 30248 6798
rect 30196 6734 30248 6740
rect 29920 6656 29972 6662
rect 29920 6598 29972 6604
rect 29736 6452 29788 6458
rect 29736 6394 29788 6400
rect 29552 6112 29604 6118
rect 29552 6054 29604 6060
rect 29564 5914 29592 6054
rect 29552 5908 29604 5914
rect 29552 5850 29604 5856
rect 29276 5772 29328 5778
rect 29276 5714 29328 5720
rect 29644 5636 29696 5642
rect 29644 5578 29696 5584
rect 29552 5568 29604 5574
rect 29552 5510 29604 5516
rect 29092 5364 29144 5370
rect 29092 5306 29144 5312
rect 29184 5364 29236 5370
rect 29184 5306 29236 5312
rect 29460 5296 29512 5302
rect 29460 5238 29512 5244
rect 29000 4820 29052 4826
rect 29000 4762 29052 4768
rect 28908 4684 28960 4690
rect 28908 4626 28960 4632
rect 28920 4214 28948 4626
rect 28908 4208 28960 4214
rect 28908 4150 28960 4156
rect 28908 4004 28960 4010
rect 28908 3946 28960 3952
rect 28920 3913 28948 3946
rect 28906 3904 28962 3913
rect 28906 3839 28962 3848
rect 28736 2746 28856 2774
rect 28630 2408 28686 2417
rect 28630 2343 28686 2352
rect 28172 1080 28224 1086
rect 28172 1022 28224 1028
rect 27710 776 27766 785
rect 27710 711 27766 720
rect 28736 56 28764 2746
rect 29472 2650 29500 5238
rect 29460 2644 29512 2650
rect 29460 2586 29512 2592
rect 29564 542 29592 5510
rect 29656 5370 29684 5578
rect 29644 5364 29696 5370
rect 29644 5306 29696 5312
rect 29828 5024 29880 5030
rect 29828 4966 29880 4972
rect 29736 4548 29788 4554
rect 29736 4490 29788 4496
rect 29748 3942 29776 4490
rect 29736 3936 29788 3942
rect 29736 3878 29788 3884
rect 29644 3392 29696 3398
rect 29644 3334 29696 3340
rect 29656 2990 29684 3334
rect 29748 3097 29776 3878
rect 29734 3088 29790 3097
rect 29734 3023 29790 3032
rect 29644 2984 29696 2990
rect 29644 2926 29696 2932
rect 29840 950 29868 4966
rect 29932 4282 29960 6598
rect 30300 6322 30328 7647
rect 30104 6316 30156 6322
rect 30104 6258 30156 6264
rect 30288 6316 30340 6322
rect 30288 6258 30340 6264
rect 30012 6248 30064 6254
rect 30012 6190 30064 6196
rect 30024 6089 30052 6190
rect 30010 6080 30066 6089
rect 30010 6015 30066 6024
rect 30024 5710 30052 6015
rect 30012 5704 30064 5710
rect 30116 5692 30144 6258
rect 30196 5840 30248 5846
rect 30392 5828 30420 8434
rect 30484 8129 30512 10134
rect 30576 10033 30604 11194
rect 30748 10124 30800 10130
rect 30748 10066 30800 10072
rect 30562 10024 30618 10033
rect 30562 9959 30618 9968
rect 30656 8560 30708 8566
rect 30656 8502 30708 8508
rect 30470 8120 30526 8129
rect 30470 8055 30526 8064
rect 30472 7948 30524 7954
rect 30472 7890 30524 7896
rect 30484 7410 30512 7890
rect 30564 7880 30616 7886
rect 30564 7822 30616 7828
rect 30576 7750 30604 7822
rect 30564 7744 30616 7750
rect 30564 7686 30616 7692
rect 30472 7404 30524 7410
rect 30472 7346 30524 7352
rect 30472 6860 30524 6866
rect 30472 6802 30524 6808
rect 30248 5800 30420 5828
rect 30196 5782 30248 5788
rect 30380 5704 30432 5710
rect 30116 5664 30236 5692
rect 30012 5646 30064 5652
rect 29920 4276 29972 4282
rect 29920 4218 29972 4224
rect 29920 4140 29972 4146
rect 29920 4082 29972 4088
rect 29932 3505 29960 4082
rect 29918 3496 29974 3505
rect 29918 3431 29974 3440
rect 30024 1630 30052 5646
rect 30208 5352 30236 5664
rect 30380 5646 30432 5652
rect 30288 5364 30340 5370
rect 30208 5324 30288 5352
rect 30288 5306 30340 5312
rect 30392 4622 30420 5646
rect 30380 4616 30432 4622
rect 30380 4558 30432 4564
rect 30104 4072 30156 4078
rect 30104 4014 30156 4020
rect 30116 3194 30144 4014
rect 30380 3936 30432 3942
rect 30380 3878 30432 3884
rect 30194 3632 30250 3641
rect 30194 3567 30250 3576
rect 30208 3398 30236 3567
rect 30196 3392 30248 3398
rect 30196 3334 30248 3340
rect 30104 3188 30156 3194
rect 30104 3130 30156 3136
rect 30392 2854 30420 3878
rect 30484 2854 30512 6802
rect 30576 6798 30604 7686
rect 30564 6792 30616 6798
rect 30564 6734 30616 6740
rect 30668 6662 30696 8502
rect 30656 6656 30708 6662
rect 30656 6598 30708 6604
rect 30656 6316 30708 6322
rect 30656 6258 30708 6264
rect 30668 6225 30696 6258
rect 30654 6216 30710 6225
rect 30654 6151 30710 6160
rect 30668 5642 30696 6151
rect 30760 5710 30788 10066
rect 30852 6730 30880 11194
rect 31128 9897 31156 11194
rect 31114 9888 31170 9897
rect 31114 9823 31170 9832
rect 31404 9382 31432 11194
rect 31680 9761 31708 11194
rect 31666 9752 31722 9761
rect 31666 9687 31722 9696
rect 31300 9376 31352 9382
rect 31300 9318 31352 9324
rect 31392 9376 31444 9382
rect 31392 9318 31444 9324
rect 30932 9172 30984 9178
rect 30932 9114 30984 9120
rect 30944 8673 30972 9114
rect 30930 8664 30986 8673
rect 30930 8599 30986 8608
rect 30932 8560 30984 8566
rect 30932 8502 30984 8508
rect 30840 6724 30892 6730
rect 30840 6666 30892 6672
rect 30838 5808 30894 5817
rect 30838 5743 30894 5752
rect 30748 5704 30800 5710
rect 30748 5646 30800 5652
rect 30656 5636 30708 5642
rect 30656 5578 30708 5584
rect 30668 5234 30696 5578
rect 30656 5228 30708 5234
rect 30656 5170 30708 5176
rect 30562 4856 30618 4865
rect 30562 4791 30618 4800
rect 30656 4820 30708 4826
rect 30576 3194 30604 4791
rect 30656 4762 30708 4768
rect 30668 4554 30696 4762
rect 30656 4548 30708 4554
rect 30656 4490 30708 4496
rect 30668 4146 30696 4490
rect 30656 4140 30708 4146
rect 30656 4082 30708 4088
rect 30656 4004 30708 4010
rect 30656 3946 30708 3952
rect 30668 3670 30696 3946
rect 30656 3664 30708 3670
rect 30656 3606 30708 3612
rect 30564 3188 30616 3194
rect 30564 3130 30616 3136
rect 30748 3188 30800 3194
rect 30748 3130 30800 3136
rect 30760 2922 30788 3130
rect 30748 2916 30800 2922
rect 30748 2858 30800 2864
rect 30380 2848 30432 2854
rect 30380 2790 30432 2796
rect 30472 2848 30524 2854
rect 30472 2790 30524 2796
rect 30392 2582 30420 2790
rect 30380 2576 30432 2582
rect 30380 2518 30432 2524
rect 30012 1624 30064 1630
rect 30012 1566 30064 1572
rect 30852 1442 30880 5743
rect 30944 2650 30972 8502
rect 31116 8424 31168 8430
rect 31116 8366 31168 8372
rect 31024 8356 31076 8362
rect 31024 8298 31076 8304
rect 31036 6934 31064 8298
rect 31128 7002 31156 8366
rect 31208 8356 31260 8362
rect 31208 8298 31260 8304
rect 31220 8090 31248 8298
rect 31208 8084 31260 8090
rect 31208 8026 31260 8032
rect 31116 6996 31168 7002
rect 31116 6938 31168 6944
rect 31024 6928 31076 6934
rect 31024 6870 31076 6876
rect 31208 6860 31260 6866
rect 31208 6802 31260 6808
rect 31114 6760 31170 6769
rect 31114 6695 31170 6704
rect 31128 6390 31156 6695
rect 31116 6384 31168 6390
rect 31116 6326 31168 6332
rect 31024 6316 31076 6322
rect 31024 6258 31076 6264
rect 31036 6089 31064 6258
rect 31022 6080 31078 6089
rect 31022 6015 31078 6024
rect 31220 5914 31248 6802
rect 31312 6338 31340 9318
rect 31956 9246 31984 11194
rect 31576 9240 31628 9246
rect 31576 9182 31628 9188
rect 31944 9240 31996 9246
rect 31944 9182 31996 9188
rect 32034 9208 32090 9217
rect 31588 9024 31616 9182
rect 32034 9143 32090 9152
rect 31588 8996 31708 9024
rect 31392 8492 31444 8498
rect 31576 8492 31628 8498
rect 31392 8434 31444 8440
rect 31496 8452 31576 8480
rect 31404 7750 31432 8434
rect 31496 7886 31524 8452
rect 31576 8434 31628 8440
rect 31576 8084 31628 8090
rect 31576 8026 31628 8032
rect 31484 7880 31536 7886
rect 31484 7822 31536 7828
rect 31392 7744 31444 7750
rect 31392 7686 31444 7692
rect 31496 7546 31524 7822
rect 31484 7540 31536 7546
rect 31484 7482 31536 7488
rect 31392 6860 31444 6866
rect 31392 6802 31444 6808
rect 31404 6458 31432 6802
rect 31496 6798 31524 7482
rect 31484 6792 31536 6798
rect 31484 6734 31536 6740
rect 31588 6458 31616 8026
rect 31680 6866 31708 8996
rect 31760 8968 31812 8974
rect 31760 8910 31812 8916
rect 31772 8498 31800 8910
rect 32048 8537 32076 9143
rect 32232 9042 32260 11194
rect 32404 10328 32456 10334
rect 32404 10270 32456 10276
rect 32312 9716 32364 9722
rect 32312 9658 32364 9664
rect 32220 9036 32272 9042
rect 32220 8978 32272 8984
rect 32128 8900 32180 8906
rect 32128 8842 32180 8848
rect 32034 8528 32090 8537
rect 31760 8492 31812 8498
rect 32140 8498 32168 8842
rect 32034 8463 32090 8472
rect 32128 8492 32180 8498
rect 31760 8434 31812 8440
rect 32128 8434 32180 8440
rect 31944 8356 31996 8362
rect 31864 8316 31944 8344
rect 31760 8288 31812 8294
rect 31760 8230 31812 8236
rect 31772 8022 31800 8230
rect 31864 8072 31892 8316
rect 31944 8298 31996 8304
rect 31950 8188 32258 8197
rect 31950 8186 31956 8188
rect 32012 8186 32036 8188
rect 32092 8186 32116 8188
rect 32172 8186 32196 8188
rect 32252 8186 32258 8188
rect 32012 8134 32014 8186
rect 32194 8134 32196 8186
rect 31950 8132 31956 8134
rect 32012 8132 32036 8134
rect 32092 8132 32116 8134
rect 32172 8132 32196 8134
rect 32252 8132 32258 8134
rect 31950 8123 32258 8132
rect 32324 8072 32352 9658
rect 32416 8537 32444 10270
rect 32402 8528 32458 8537
rect 32402 8463 32458 8472
rect 32508 8430 32536 11194
rect 32588 9376 32640 9382
rect 32588 9318 32640 9324
rect 32404 8424 32456 8430
rect 32404 8366 32456 8372
rect 32496 8424 32548 8430
rect 32496 8366 32548 8372
rect 32416 8265 32444 8366
rect 32402 8256 32458 8265
rect 32402 8191 32458 8200
rect 32600 8106 32628 9318
rect 32784 8362 32812 11194
rect 33060 8974 33088 11194
rect 33048 8968 33100 8974
rect 33048 8910 33100 8916
rect 33336 8838 33364 11194
rect 33506 9888 33562 9897
rect 33506 9823 33562 9832
rect 33414 9616 33470 9625
rect 33414 9551 33470 9560
rect 33324 8832 33376 8838
rect 33324 8774 33376 8780
rect 33010 8732 33318 8741
rect 33010 8730 33016 8732
rect 33072 8730 33096 8732
rect 33152 8730 33176 8732
rect 33232 8730 33256 8732
rect 33312 8730 33318 8732
rect 33072 8678 33074 8730
rect 33254 8678 33256 8730
rect 33010 8676 33016 8678
rect 33072 8676 33096 8678
rect 33152 8676 33176 8678
rect 33232 8676 33256 8678
rect 33312 8676 33318 8678
rect 32862 8664 32918 8673
rect 33010 8667 33318 8676
rect 32862 8599 32864 8608
rect 32916 8599 32918 8608
rect 32864 8570 32916 8576
rect 32954 8528 33010 8537
rect 32954 8463 33010 8472
rect 33048 8492 33100 8498
rect 32772 8356 32824 8362
rect 32772 8298 32824 8304
rect 32864 8288 32916 8294
rect 31864 8044 31984 8072
rect 31760 8016 31812 8022
rect 31760 7958 31812 7964
rect 31760 7880 31812 7886
rect 31760 7822 31812 7828
rect 31772 7324 31800 7822
rect 31956 7750 31984 8044
rect 32232 8044 32352 8072
rect 32416 8078 32628 8106
rect 32692 8236 32864 8242
rect 32692 8230 32916 8236
rect 32692 8214 32904 8230
rect 32232 7886 32260 8044
rect 32220 7880 32272 7886
rect 32220 7822 32272 7828
rect 31944 7744 31996 7750
rect 31944 7686 31996 7692
rect 32128 7744 32180 7750
rect 32128 7686 32180 7692
rect 32218 7712 32274 7721
rect 32140 7478 32168 7686
rect 32218 7647 32274 7656
rect 32232 7478 32260 7647
rect 32128 7472 32180 7478
rect 32128 7414 32180 7420
rect 32220 7472 32272 7478
rect 32220 7414 32272 7420
rect 31944 7336 31996 7342
rect 31772 7296 31944 7324
rect 31944 7278 31996 7284
rect 32220 7268 32272 7274
rect 32272 7228 32352 7256
rect 32220 7210 32272 7216
rect 31944 7200 31996 7206
rect 31758 7168 31814 7177
rect 31864 7160 31944 7188
rect 31864 7154 31892 7160
rect 31814 7126 31892 7154
rect 31944 7142 31996 7148
rect 31758 7103 31814 7112
rect 31950 7100 32258 7109
rect 31950 7098 31956 7100
rect 32012 7098 32036 7100
rect 32092 7098 32116 7100
rect 32172 7098 32196 7100
rect 32252 7098 32258 7100
rect 32012 7046 32014 7098
rect 32194 7046 32196 7098
rect 31950 7044 31956 7046
rect 32012 7044 32036 7046
rect 32092 7044 32116 7046
rect 32172 7044 32196 7046
rect 32252 7044 32258 7046
rect 31758 7032 31814 7041
rect 31950 7035 32258 7044
rect 32324 7002 32352 7228
rect 31758 6967 31814 6976
rect 32312 6996 32364 7002
rect 31668 6860 31720 6866
rect 31668 6802 31720 6808
rect 31666 6760 31722 6769
rect 31772 6746 31800 6967
rect 32312 6938 32364 6944
rect 32416 6798 32444 8078
rect 32496 8016 32548 8022
rect 32496 7958 32548 7964
rect 32508 7290 32536 7958
rect 32588 7880 32640 7886
rect 32588 7822 32640 7828
rect 32600 7410 32628 7822
rect 32588 7404 32640 7410
rect 32588 7346 32640 7352
rect 32508 7262 32628 7290
rect 32496 7200 32548 7206
rect 32496 7142 32548 7148
rect 32036 6792 32088 6798
rect 32034 6760 32036 6769
rect 32404 6792 32456 6798
rect 32088 6760 32090 6769
rect 31772 6718 31984 6746
rect 31666 6695 31668 6704
rect 31720 6695 31722 6704
rect 31668 6666 31720 6672
rect 31852 6656 31904 6662
rect 31680 6582 31800 6610
rect 31852 6598 31904 6604
rect 31392 6452 31444 6458
rect 31392 6394 31444 6400
rect 31576 6452 31628 6458
rect 31576 6394 31628 6400
rect 31680 6338 31708 6582
rect 31312 6310 31708 6338
rect 31772 6322 31800 6582
rect 31760 6316 31812 6322
rect 31760 6258 31812 6264
rect 31758 6216 31814 6225
rect 31758 6151 31814 6160
rect 31300 6112 31352 6118
rect 31300 6054 31352 6060
rect 31208 5908 31260 5914
rect 31208 5850 31260 5856
rect 31114 5400 31170 5409
rect 31114 5335 31170 5344
rect 31128 4622 31156 5335
rect 31208 5160 31260 5166
rect 31208 5102 31260 5108
rect 31116 4616 31168 4622
rect 31116 4558 31168 4564
rect 31128 3942 31156 4558
rect 31116 3936 31168 3942
rect 31116 3878 31168 3884
rect 31128 3602 31156 3878
rect 31116 3596 31168 3602
rect 31116 3538 31168 3544
rect 31220 3126 31248 5102
rect 31312 4078 31340 6054
rect 31574 5128 31630 5137
rect 31574 5063 31630 5072
rect 31300 4072 31352 4078
rect 31300 4014 31352 4020
rect 31588 3534 31616 5063
rect 31668 4684 31720 4690
rect 31668 4626 31720 4632
rect 31680 4214 31708 4626
rect 31668 4208 31720 4214
rect 31668 4150 31720 4156
rect 31772 4010 31800 6151
rect 31864 4729 31892 6598
rect 31956 6458 31984 6718
rect 32404 6734 32456 6740
rect 32034 6695 32090 6704
rect 32036 6656 32088 6662
rect 32312 6656 32364 6662
rect 32036 6598 32088 6604
rect 32310 6624 32312 6633
rect 32364 6624 32366 6633
rect 31944 6452 31996 6458
rect 31944 6394 31996 6400
rect 32048 6118 32076 6598
rect 32310 6559 32366 6568
rect 32312 6248 32364 6254
rect 32364 6208 32444 6236
rect 32312 6190 32364 6196
rect 32036 6112 32088 6118
rect 32036 6054 32088 6060
rect 32312 6112 32364 6118
rect 32312 6054 32364 6060
rect 31950 6012 32258 6021
rect 31950 6010 31956 6012
rect 32012 6010 32036 6012
rect 32092 6010 32116 6012
rect 32172 6010 32196 6012
rect 32252 6010 32258 6012
rect 32012 5958 32014 6010
rect 32194 5958 32196 6010
rect 31950 5956 31956 5958
rect 32012 5956 32036 5958
rect 32092 5956 32116 5958
rect 32172 5956 32196 5958
rect 32252 5956 32258 5958
rect 31950 5947 32258 5956
rect 32036 5704 32088 5710
rect 32220 5704 32272 5710
rect 32036 5646 32088 5652
rect 32218 5672 32220 5681
rect 32272 5672 32274 5681
rect 32048 5302 32076 5646
rect 32218 5607 32274 5616
rect 32036 5296 32088 5302
rect 32036 5238 32088 5244
rect 31950 4924 32258 4933
rect 31950 4922 31956 4924
rect 32012 4922 32036 4924
rect 32092 4922 32116 4924
rect 32172 4922 32196 4924
rect 32252 4922 32258 4924
rect 32012 4870 32014 4922
rect 32194 4870 32196 4922
rect 31950 4868 31956 4870
rect 32012 4868 32036 4870
rect 32092 4868 32116 4870
rect 32172 4868 32196 4870
rect 32252 4868 32258 4870
rect 31950 4859 32258 4868
rect 31850 4720 31906 4729
rect 32034 4720 32090 4729
rect 31850 4655 31906 4664
rect 31956 4678 32034 4706
rect 31956 4026 31984 4678
rect 32034 4655 32090 4664
rect 32220 4616 32272 4622
rect 32220 4558 32272 4564
rect 31760 4004 31812 4010
rect 31760 3946 31812 3952
rect 31864 3998 31984 4026
rect 31576 3528 31628 3534
rect 31628 3488 31708 3516
rect 31576 3470 31628 3476
rect 31208 3120 31260 3126
rect 31208 3062 31260 3068
rect 31484 3120 31536 3126
rect 31484 3062 31536 3068
rect 30932 2644 30984 2650
rect 30932 2586 30984 2592
rect 31392 2644 31444 2650
rect 31392 2586 31444 2592
rect 31404 2378 31432 2586
rect 31496 2582 31524 3062
rect 31680 3058 31708 3488
rect 31576 3052 31628 3058
rect 31576 2994 31628 3000
rect 31668 3052 31720 3058
rect 31668 2994 31720 3000
rect 31484 2576 31536 2582
rect 31484 2518 31536 2524
rect 31588 2514 31616 2994
rect 31576 2508 31628 2514
rect 31576 2450 31628 2456
rect 31392 2372 31444 2378
rect 31392 2314 31444 2320
rect 31588 1698 31616 2450
rect 31680 2446 31708 2994
rect 31864 2774 31892 3998
rect 32232 3924 32260 4558
rect 32324 4026 32352 6054
rect 32416 5370 32444 6208
rect 32404 5364 32456 5370
rect 32404 5306 32456 5312
rect 32416 4622 32444 5306
rect 32508 4622 32536 7142
rect 32404 4616 32456 4622
rect 32404 4558 32456 4564
rect 32496 4616 32548 4622
rect 32496 4558 32548 4564
rect 32600 4554 32628 7262
rect 32588 4548 32640 4554
rect 32588 4490 32640 4496
rect 32404 4480 32456 4486
rect 32404 4422 32456 4428
rect 32416 4146 32444 4422
rect 32404 4140 32456 4146
rect 32404 4082 32456 4088
rect 32588 4072 32640 4078
rect 32324 3998 32536 4026
rect 32588 4014 32640 4020
rect 32232 3896 32352 3924
rect 31950 3836 32258 3845
rect 31950 3834 31956 3836
rect 32012 3834 32036 3836
rect 32092 3834 32116 3836
rect 32172 3834 32196 3836
rect 32252 3834 32258 3836
rect 32012 3782 32014 3834
rect 32194 3782 32196 3834
rect 31950 3780 31956 3782
rect 32012 3780 32036 3782
rect 32092 3780 32116 3782
rect 32172 3780 32196 3782
rect 32252 3780 32258 3782
rect 31950 3771 32258 3780
rect 32324 3720 32352 3896
rect 32140 3692 32352 3720
rect 31944 3528 31996 3534
rect 31944 3470 31996 3476
rect 31956 3126 31984 3470
rect 31944 3120 31996 3126
rect 32140 3097 32168 3692
rect 32312 3528 32364 3534
rect 32312 3470 32364 3476
rect 32220 3392 32272 3398
rect 32220 3334 32272 3340
rect 32232 3126 32260 3334
rect 32220 3120 32272 3126
rect 31944 3062 31996 3068
rect 32126 3088 32182 3097
rect 31956 2990 31984 3062
rect 32220 3062 32272 3068
rect 32126 3023 32182 3032
rect 32140 2990 32168 3023
rect 31944 2984 31996 2990
rect 31944 2926 31996 2932
rect 32128 2984 32180 2990
rect 32128 2926 32180 2932
rect 31772 2746 31892 2774
rect 31950 2748 32258 2757
rect 31950 2746 31956 2748
rect 32012 2746 32036 2748
rect 32092 2746 32116 2748
rect 32172 2746 32196 2748
rect 32252 2746 32258 2748
rect 31668 2440 31720 2446
rect 31668 2382 31720 2388
rect 31576 1692 31628 1698
rect 31576 1634 31628 1640
rect 30852 1414 30972 1442
rect 29828 944 29880 950
rect 29828 886 29880 892
rect 29826 776 29882 785
rect 29826 711 29882 720
rect 29552 536 29604 542
rect 29552 478 29604 484
rect 29840 56 29868 711
rect 30944 56 30972 1414
rect 22192 2 22244 8
rect 23202 0 23258 56
rect 24306 0 24362 56
rect 25410 0 25466 56
rect 26514 0 26570 56
rect 27618 0 27674 56
rect 28722 0 28778 56
rect 29826 0 29882 56
rect 30930 0 30986 56
rect 31772 42 31800 2746
rect 32012 2694 32014 2746
rect 32194 2694 32196 2746
rect 31950 2692 31956 2694
rect 32012 2692 32036 2694
rect 32092 2692 32116 2694
rect 32172 2692 32196 2694
rect 32252 2692 32258 2694
rect 31950 2683 32258 2692
rect 32324 2650 32352 3470
rect 32312 2644 32364 2650
rect 32312 2586 32364 2592
rect 32508 1494 32536 3998
rect 32600 3040 32628 4014
rect 32692 3108 32720 8214
rect 32770 8120 32826 8129
rect 32770 8055 32826 8064
rect 32784 8022 32812 8055
rect 32772 8016 32824 8022
rect 32772 7958 32824 7964
rect 32862 7984 32918 7993
rect 32862 7919 32918 7928
rect 32772 7812 32824 7818
rect 32772 7754 32824 7760
rect 32784 7410 32812 7754
rect 32772 7404 32824 7410
rect 32772 7346 32824 7352
rect 32876 7290 32904 7919
rect 32968 7818 32996 8463
rect 33048 8434 33100 8440
rect 33060 8090 33088 8434
rect 33230 8256 33286 8265
rect 33230 8191 33286 8200
rect 33048 8084 33100 8090
rect 33048 8026 33100 8032
rect 33244 7886 33272 8191
rect 33428 8090 33456 9551
rect 33416 8084 33468 8090
rect 33416 8026 33468 8032
rect 33520 7886 33548 9823
rect 33612 8362 33640 11194
rect 33782 9888 33838 9897
rect 33782 9823 33838 9832
rect 33796 9790 33824 9823
rect 33784 9784 33836 9790
rect 33690 9752 33746 9761
rect 33784 9726 33836 9732
rect 33690 9687 33746 9696
rect 33600 8356 33652 8362
rect 33600 8298 33652 8304
rect 33232 7880 33284 7886
rect 33232 7822 33284 7828
rect 33508 7880 33560 7886
rect 33508 7822 33560 7828
rect 33598 7848 33654 7857
rect 32956 7812 33008 7818
rect 33704 7818 33732 9687
rect 33784 8832 33836 8838
rect 33784 8774 33836 8780
rect 33796 8294 33824 8774
rect 33888 8566 33916 11194
rect 34058 10024 34114 10033
rect 34058 9959 34114 9968
rect 33968 9240 34020 9246
rect 33968 9182 34020 9188
rect 33876 8560 33928 8566
rect 33876 8502 33928 8508
rect 33876 8424 33928 8430
rect 33876 8366 33928 8372
rect 33784 8288 33836 8294
rect 33784 8230 33836 8236
rect 33598 7783 33654 7792
rect 33692 7812 33744 7818
rect 32956 7754 33008 7760
rect 33612 7750 33640 7783
rect 33692 7754 33744 7760
rect 33600 7744 33652 7750
rect 33600 7686 33652 7692
rect 33010 7644 33318 7653
rect 33010 7642 33016 7644
rect 33072 7642 33096 7644
rect 33152 7642 33176 7644
rect 33232 7642 33256 7644
rect 33312 7642 33318 7644
rect 33072 7590 33074 7642
rect 33254 7590 33256 7642
rect 33010 7588 33016 7590
rect 33072 7588 33096 7590
rect 33152 7588 33176 7590
rect 33232 7588 33256 7590
rect 33312 7588 33318 7590
rect 33010 7579 33318 7588
rect 32956 7540 33008 7546
rect 32956 7482 33008 7488
rect 33048 7540 33100 7546
rect 33048 7482 33100 7488
rect 32968 7449 32996 7482
rect 32954 7440 33010 7449
rect 32954 7375 33010 7384
rect 33060 7290 33088 7482
rect 33784 7336 33836 7342
rect 32876 7262 33088 7290
rect 33230 7304 33286 7313
rect 33230 7239 33232 7248
rect 33284 7239 33286 7248
rect 33704 7284 33784 7290
rect 33704 7278 33836 7284
rect 33704 7262 33824 7278
rect 33232 7210 33284 7216
rect 32954 6896 33010 6905
rect 32954 6831 33010 6840
rect 32968 6798 32996 6831
rect 32956 6792 33008 6798
rect 32956 6734 33008 6740
rect 32772 6724 32824 6730
rect 32772 6666 32824 6672
rect 32784 5409 32812 6666
rect 33010 6556 33318 6565
rect 33010 6554 33016 6556
rect 33072 6554 33096 6556
rect 33152 6554 33176 6556
rect 33232 6554 33256 6556
rect 33312 6554 33318 6556
rect 33072 6502 33074 6554
rect 33254 6502 33256 6554
rect 33010 6500 33016 6502
rect 33072 6500 33096 6502
rect 33152 6500 33176 6502
rect 33232 6500 33256 6502
rect 33312 6500 33318 6502
rect 33010 6491 33318 6500
rect 33416 6112 33468 6118
rect 33416 6054 33468 6060
rect 33230 5944 33286 5953
rect 33230 5879 33286 5888
rect 32956 5772 33008 5778
rect 32956 5714 33008 5720
rect 32862 5672 32918 5681
rect 32862 5607 32918 5616
rect 32770 5400 32826 5409
rect 32770 5335 32826 5344
rect 32876 4729 32904 5607
rect 32968 5574 32996 5714
rect 33244 5574 33272 5879
rect 33428 5710 33456 6054
rect 33416 5704 33468 5710
rect 33416 5646 33468 5652
rect 32956 5568 33008 5574
rect 32956 5510 33008 5516
rect 33232 5568 33284 5574
rect 33232 5510 33284 5516
rect 33010 5468 33318 5477
rect 33010 5466 33016 5468
rect 33072 5466 33096 5468
rect 33152 5466 33176 5468
rect 33232 5466 33256 5468
rect 33312 5466 33318 5468
rect 33072 5414 33074 5466
rect 33254 5414 33256 5466
rect 33010 5412 33016 5414
rect 33072 5412 33096 5414
rect 33152 5412 33176 5414
rect 33232 5412 33256 5414
rect 33312 5412 33318 5414
rect 33010 5403 33318 5412
rect 33508 5024 33560 5030
rect 33508 4966 33560 4972
rect 32862 4720 32918 4729
rect 33520 4690 33548 4966
rect 33600 4752 33652 4758
rect 33600 4694 33652 4700
rect 32862 4655 32918 4664
rect 33508 4684 33560 4690
rect 33508 4626 33560 4632
rect 33612 4570 33640 4694
rect 33520 4542 33640 4570
rect 32864 4480 32916 4486
rect 32864 4422 32916 4428
rect 32876 4146 32904 4422
rect 33010 4380 33318 4389
rect 33010 4378 33016 4380
rect 33072 4378 33096 4380
rect 33152 4378 33176 4380
rect 33232 4378 33256 4380
rect 33312 4378 33318 4380
rect 33072 4326 33074 4378
rect 33254 4326 33256 4378
rect 33010 4324 33016 4326
rect 33072 4324 33096 4326
rect 33152 4324 33176 4326
rect 33232 4324 33256 4326
rect 33312 4324 33318 4326
rect 33010 4315 33318 4324
rect 32954 4176 33010 4185
rect 32864 4140 32916 4146
rect 32954 4111 33010 4120
rect 33416 4140 33468 4146
rect 32864 4082 32916 4088
rect 32772 3936 32824 3942
rect 32772 3878 32824 3884
rect 32784 3233 32812 3878
rect 32864 3664 32916 3670
rect 32864 3606 32916 3612
rect 32770 3224 32826 3233
rect 32876 3194 32904 3606
rect 32968 3398 32996 4111
rect 33416 4082 33468 4088
rect 32956 3392 33008 3398
rect 32956 3334 33008 3340
rect 33010 3292 33318 3301
rect 33010 3290 33016 3292
rect 33072 3290 33096 3292
rect 33152 3290 33176 3292
rect 33232 3290 33256 3292
rect 33312 3290 33318 3292
rect 33072 3238 33074 3290
rect 33254 3238 33256 3290
rect 33010 3236 33016 3238
rect 33072 3236 33096 3238
rect 33152 3236 33176 3238
rect 33232 3236 33256 3238
rect 33312 3236 33318 3238
rect 33010 3227 33318 3236
rect 32770 3159 32826 3168
rect 32864 3188 32916 3194
rect 32864 3130 32916 3136
rect 33048 3120 33100 3126
rect 32692 3080 32812 3108
rect 32600 3012 32720 3040
rect 32586 2816 32642 2825
rect 32586 2751 32642 2760
rect 32600 1970 32628 2751
rect 32692 2446 32720 3012
rect 32784 2446 32812 3080
rect 32968 3080 33048 3108
rect 32864 3052 32916 3058
rect 32864 2994 32916 3000
rect 32876 2922 32904 2994
rect 32864 2916 32916 2922
rect 32864 2858 32916 2864
rect 32680 2440 32732 2446
rect 32680 2382 32732 2388
rect 32772 2440 32824 2446
rect 32772 2382 32824 2388
rect 32876 2310 32904 2858
rect 32968 2825 32996 3080
rect 33428 3097 33456 4082
rect 33048 3062 33100 3068
rect 33414 3088 33470 3097
rect 33414 3023 33416 3032
rect 33468 3023 33470 3032
rect 33416 2994 33468 3000
rect 33048 2848 33100 2854
rect 32954 2816 33010 2825
rect 33048 2790 33100 2796
rect 32954 2751 33010 2760
rect 33060 2514 33088 2790
rect 33048 2508 33100 2514
rect 33048 2450 33100 2456
rect 32864 2304 32916 2310
rect 32864 2246 32916 2252
rect 33416 2304 33468 2310
rect 33416 2246 33468 2252
rect 33010 2204 33318 2213
rect 33010 2202 33016 2204
rect 33072 2202 33096 2204
rect 33152 2202 33176 2204
rect 33232 2202 33256 2204
rect 33312 2202 33318 2204
rect 33072 2150 33074 2202
rect 33254 2150 33256 2202
rect 33010 2148 33016 2150
rect 33072 2148 33096 2150
rect 33152 2148 33176 2150
rect 33232 2148 33256 2150
rect 33312 2148 33318 2150
rect 33010 2139 33318 2148
rect 32588 1964 32640 1970
rect 32588 1906 32640 1912
rect 33428 1766 33456 2246
rect 33416 1760 33468 1766
rect 33416 1702 33468 1708
rect 32496 1488 32548 1494
rect 32496 1430 32548 1436
rect 33520 1057 33548 4542
rect 33704 4434 33732 7262
rect 33784 7200 33836 7206
rect 33784 7142 33836 7148
rect 33612 4406 33732 4434
rect 33506 1048 33562 1057
rect 33506 983 33562 992
rect 31956 56 32076 82
rect 33152 56 33272 82
rect 31956 54 32090 56
rect 31956 42 31984 54
rect 31772 14 31984 42
rect 32034 0 32090 54
rect 33138 54 33272 56
rect 33138 0 33194 54
rect 33244 42 33272 54
rect 33612 42 33640 4406
rect 33796 4078 33824 7142
rect 33888 5250 33916 8366
rect 33980 7410 34008 9182
rect 34072 8378 34100 9959
rect 34164 8498 34192 11194
rect 34244 9444 34296 9450
rect 34244 9386 34296 9392
rect 34152 8492 34204 8498
rect 34152 8434 34204 8440
rect 34072 8350 34192 8378
rect 34164 7478 34192 8350
rect 34152 7472 34204 7478
rect 34152 7414 34204 7420
rect 34256 7410 34284 9386
rect 34336 8900 34388 8906
rect 34336 8842 34388 8848
rect 34348 8498 34376 8842
rect 34336 8492 34388 8498
rect 34440 8480 34468 11194
rect 34610 9344 34666 9353
rect 34610 9279 34666 9288
rect 34520 8968 34572 8974
rect 34520 8910 34572 8916
rect 34532 8634 34560 8910
rect 34520 8628 34572 8634
rect 34520 8570 34572 8576
rect 34440 8452 34560 8480
rect 34336 8434 34388 8440
rect 34532 8090 34560 8452
rect 34520 8084 34572 8090
rect 34520 8026 34572 8032
rect 34624 7970 34652 9279
rect 34716 8362 34744 11194
rect 34992 9194 35020 11194
rect 34992 9166 35204 9194
rect 34980 9104 35032 9110
rect 34980 9046 35032 9052
rect 34796 9036 34848 9042
rect 34796 8978 34848 8984
rect 34704 8356 34756 8362
rect 34704 8298 34756 8304
rect 34440 7942 34652 7970
rect 34440 7546 34468 7942
rect 34428 7540 34480 7546
rect 34428 7482 34480 7488
rect 34612 7472 34664 7478
rect 34612 7414 34664 7420
rect 33968 7404 34020 7410
rect 33968 7346 34020 7352
rect 34244 7404 34296 7410
rect 34244 7346 34296 7352
rect 34520 7404 34572 7410
rect 34520 7346 34572 7352
rect 34532 7002 34560 7346
rect 34520 6996 34572 7002
rect 34520 6938 34572 6944
rect 34060 6656 34112 6662
rect 34060 6598 34112 6604
rect 34152 6656 34204 6662
rect 34152 6598 34204 6604
rect 34072 6458 34100 6598
rect 34060 6452 34112 6458
rect 34060 6394 34112 6400
rect 34164 5846 34192 6598
rect 34520 6316 34572 6322
rect 34520 6258 34572 6264
rect 34152 5840 34204 5846
rect 34152 5782 34204 5788
rect 34532 5710 34560 6258
rect 34624 5778 34652 7414
rect 34808 7206 34836 8978
rect 34888 8492 34940 8498
rect 34888 8434 34940 8440
rect 34796 7200 34848 7206
rect 34796 7142 34848 7148
rect 34796 6724 34848 6730
rect 34796 6666 34848 6672
rect 34808 5778 34836 6666
rect 34900 6458 34928 8434
rect 34888 6452 34940 6458
rect 34888 6394 34940 6400
rect 34888 6248 34940 6254
rect 34888 6190 34940 6196
rect 34612 5772 34664 5778
rect 34612 5714 34664 5720
rect 34796 5772 34848 5778
rect 34796 5714 34848 5720
rect 34520 5704 34572 5710
rect 34520 5646 34572 5652
rect 34808 5574 34836 5714
rect 34796 5568 34848 5574
rect 34796 5510 34848 5516
rect 33888 5222 34008 5250
rect 33876 5160 33928 5166
rect 33876 5102 33928 5108
rect 33784 4072 33836 4078
rect 33784 4014 33836 4020
rect 33692 3052 33744 3058
rect 33692 2994 33744 3000
rect 33704 2446 33732 2994
rect 33692 2440 33744 2446
rect 33692 2382 33744 2388
rect 33888 1018 33916 5102
rect 33980 3398 34008 5222
rect 34900 4146 34928 6190
rect 34992 4214 35020 9046
rect 35176 8430 35204 9166
rect 35164 8424 35216 8430
rect 35164 8366 35216 8372
rect 35268 8294 35296 11194
rect 35438 9208 35494 9217
rect 35438 9143 35494 9152
rect 35348 8968 35400 8974
rect 35348 8910 35400 8916
rect 35360 8498 35388 8910
rect 35348 8492 35400 8498
rect 35348 8434 35400 8440
rect 35256 8288 35308 8294
rect 35256 8230 35308 8236
rect 35452 6798 35480 9143
rect 35544 8090 35572 11194
rect 35624 9920 35676 9926
rect 35624 9862 35676 9868
rect 35532 8084 35584 8090
rect 35532 8026 35584 8032
rect 35440 6792 35492 6798
rect 35440 6734 35492 6740
rect 35348 6316 35400 6322
rect 35452 6304 35480 6734
rect 35636 6662 35664 9862
rect 35716 8832 35768 8838
rect 35716 8774 35768 8780
rect 35728 8498 35756 8774
rect 35820 8634 35848 11194
rect 35808 8628 35860 8634
rect 35808 8570 35860 8576
rect 35716 8492 35768 8498
rect 35716 8434 35768 8440
rect 35900 8492 35952 8498
rect 35900 8434 35952 8440
rect 35808 6996 35860 7002
rect 35808 6938 35860 6944
rect 35716 6928 35768 6934
rect 35716 6870 35768 6876
rect 35624 6656 35676 6662
rect 35624 6598 35676 6604
rect 35532 6452 35584 6458
rect 35532 6394 35584 6400
rect 35400 6276 35480 6304
rect 35348 6258 35400 6264
rect 35256 6112 35308 6118
rect 35256 6054 35308 6060
rect 35268 5556 35296 6054
rect 35544 5710 35572 6394
rect 35624 6316 35676 6322
rect 35624 6258 35676 6264
rect 35532 5704 35584 5710
rect 35532 5646 35584 5652
rect 35084 5528 35296 5556
rect 35532 5568 35584 5574
rect 34980 4208 35032 4214
rect 34980 4150 35032 4156
rect 34888 4140 34940 4146
rect 34888 4082 34940 4088
rect 33968 3392 34020 3398
rect 33968 3334 34020 3340
rect 34428 3392 34480 3398
rect 34428 3334 34480 3340
rect 34244 3120 34296 3126
rect 34244 3062 34296 3068
rect 33876 1012 33928 1018
rect 33876 954 33928 960
rect 34256 56 34284 3062
rect 34440 2938 34468 3334
rect 34336 2916 34388 2922
rect 34440 2910 34744 2938
rect 34336 2858 34388 2864
rect 34348 2802 34376 2858
rect 34716 2854 34744 2910
rect 34704 2848 34756 2854
rect 34348 2774 34560 2802
rect 34704 2790 34756 2796
rect 34532 2446 34560 2774
rect 34520 2440 34572 2446
rect 34520 2382 34572 2388
rect 34612 2440 34664 2446
rect 34612 2382 34664 2388
rect 34624 2038 34652 2382
rect 34612 2032 34664 2038
rect 34612 1974 34664 1980
rect 35084 1358 35112 5528
rect 35532 5510 35584 5516
rect 35254 5264 35310 5273
rect 35254 5199 35310 5208
rect 35268 3602 35296 5199
rect 35544 4622 35572 5510
rect 35440 4616 35492 4622
rect 35438 4584 35440 4593
rect 35532 4616 35584 4622
rect 35492 4584 35494 4593
rect 35532 4558 35584 4564
rect 35438 4519 35494 4528
rect 35348 4480 35400 4486
rect 35348 4422 35400 4428
rect 35256 3596 35308 3602
rect 35256 3538 35308 3544
rect 35072 1352 35124 1358
rect 35072 1294 35124 1300
rect 35360 56 35388 4422
rect 35452 4146 35480 4519
rect 35440 4140 35492 4146
rect 35440 4082 35492 4088
rect 35636 2774 35664 6258
rect 35728 2922 35756 6870
rect 35820 4282 35848 6938
rect 35912 6866 35940 8434
rect 36096 8090 36124 11194
rect 36372 8362 36400 11194
rect 36544 8900 36596 8906
rect 36544 8842 36596 8848
rect 36360 8356 36412 8362
rect 36360 8298 36412 8304
rect 36084 8084 36136 8090
rect 36084 8026 36136 8032
rect 36360 7880 36412 7886
rect 36360 7822 36412 7828
rect 36452 7880 36504 7886
rect 36452 7822 36504 7828
rect 35992 7200 36044 7206
rect 35992 7142 36044 7148
rect 35900 6860 35952 6866
rect 35900 6802 35952 6808
rect 36004 4826 36032 7142
rect 36084 6792 36136 6798
rect 36084 6734 36136 6740
rect 36176 6792 36228 6798
rect 36176 6734 36228 6740
rect 36096 6458 36124 6734
rect 36084 6452 36136 6458
rect 36084 6394 36136 6400
rect 36188 6322 36216 6734
rect 36176 6316 36228 6322
rect 36176 6258 36228 6264
rect 36268 6248 36320 6254
rect 36268 6190 36320 6196
rect 35992 4820 36044 4826
rect 35992 4762 36044 4768
rect 35808 4276 35860 4282
rect 35808 4218 35860 4224
rect 36280 4146 36308 6190
rect 36372 5846 36400 7822
rect 36464 7546 36492 7822
rect 36452 7540 36504 7546
rect 36452 7482 36504 7488
rect 36360 5840 36412 5846
rect 36360 5782 36412 5788
rect 36556 5370 36584 8842
rect 36648 8090 36676 11194
rect 36924 8634 36952 11194
rect 36912 8628 36964 8634
rect 36912 8570 36964 8576
rect 36728 8492 36780 8498
rect 36728 8434 36780 8440
rect 36820 8492 36872 8498
rect 36820 8434 36872 8440
rect 36636 8084 36688 8090
rect 36636 8026 36688 8032
rect 36740 6662 36768 8434
rect 36728 6656 36780 6662
rect 36728 6598 36780 6604
rect 36636 6384 36688 6390
rect 36636 6326 36688 6332
rect 36648 5914 36676 6326
rect 36832 5914 36860 8434
rect 37200 8362 37228 11194
rect 37372 8832 37424 8838
rect 37372 8774 37424 8780
rect 37280 8492 37332 8498
rect 37280 8434 37332 8440
rect 37188 8356 37240 8362
rect 37188 8298 37240 8304
rect 37004 7880 37056 7886
rect 37004 7822 37056 7828
rect 36912 6452 36964 6458
rect 36912 6394 36964 6400
rect 36636 5908 36688 5914
rect 36636 5850 36688 5856
rect 36820 5908 36872 5914
rect 36820 5850 36872 5856
rect 36544 5364 36596 5370
rect 36544 5306 36596 5312
rect 36452 4548 36504 4554
rect 36452 4490 36504 4496
rect 36268 4140 36320 4146
rect 36268 4082 36320 4088
rect 35992 3936 36044 3942
rect 35992 3878 36044 3884
rect 36004 3534 36032 3878
rect 35992 3528 36044 3534
rect 35992 3470 36044 3476
rect 35808 3392 35860 3398
rect 35808 3334 35860 3340
rect 35716 2916 35768 2922
rect 35716 2858 35768 2864
rect 35636 2746 35756 2774
rect 35728 785 35756 2746
rect 35820 921 35848 3334
rect 36280 3194 36308 4082
rect 36268 3188 36320 3194
rect 36268 3130 36320 3136
rect 35806 912 35862 921
rect 35806 847 35862 856
rect 35714 776 35770 785
rect 35714 711 35770 720
rect 36464 56 36492 4490
rect 36636 4140 36688 4146
rect 36636 4082 36688 4088
rect 36648 2961 36676 4082
rect 36634 2952 36690 2961
rect 36634 2887 36690 2896
rect 36924 1834 36952 6394
rect 37016 4826 37044 7822
rect 37292 6934 37320 8434
rect 37384 7970 37412 8774
rect 37476 8566 37504 11194
rect 37464 8560 37516 8566
rect 37464 8502 37516 8508
rect 37648 8492 37700 8498
rect 37648 8434 37700 8440
rect 37384 7942 37504 7970
rect 37372 7880 37424 7886
rect 37372 7822 37424 7828
rect 37280 6928 37332 6934
rect 37280 6870 37332 6876
rect 37096 6316 37148 6322
rect 37096 6258 37148 6264
rect 37004 4820 37056 4826
rect 37004 4762 37056 4768
rect 37108 2009 37136 6258
rect 37278 5808 37334 5817
rect 37278 5743 37280 5752
rect 37332 5743 37334 5752
rect 37280 5714 37332 5720
rect 37278 5672 37334 5681
rect 37278 5607 37280 5616
rect 37332 5607 37334 5616
rect 37280 5578 37332 5584
rect 37278 4040 37334 4049
rect 37278 3975 37334 3984
rect 37292 3602 37320 3975
rect 37280 3596 37332 3602
rect 37280 3538 37332 3544
rect 37384 3194 37412 7822
rect 37476 4010 37504 7942
rect 37556 7812 37608 7818
rect 37556 7754 37608 7760
rect 37568 6186 37596 7754
rect 37556 6180 37608 6186
rect 37556 6122 37608 6128
rect 37556 5636 37608 5642
rect 37556 5578 37608 5584
rect 37464 4004 37516 4010
rect 37464 3946 37516 3952
rect 37372 3188 37424 3194
rect 37372 3130 37424 3136
rect 37464 2372 37516 2378
rect 37464 2314 37516 2320
rect 37476 2106 37504 2314
rect 37464 2100 37516 2106
rect 37464 2042 37516 2048
rect 37094 2000 37150 2009
rect 37094 1935 37150 1944
rect 36912 1828 36964 1834
rect 36912 1770 36964 1776
rect 37568 56 37596 5578
rect 37660 4826 37688 8434
rect 37752 8090 37780 11194
rect 39762 9888 39818 9897
rect 39762 9823 39818 9832
rect 39670 9616 39726 9625
rect 39670 9551 39726 9560
rect 38934 9344 38990 9353
rect 38568 9308 38620 9314
rect 38934 9279 38990 9288
rect 38568 9250 38620 9256
rect 38384 8968 38436 8974
rect 38384 8910 38436 8916
rect 37832 8424 37884 8430
rect 37832 8366 37884 8372
rect 37740 8084 37792 8090
rect 37740 8026 37792 8032
rect 37740 7812 37792 7818
rect 37740 7754 37792 7760
rect 37752 5386 37780 7754
rect 37844 5914 37872 8366
rect 37950 8188 38258 8197
rect 37950 8186 37956 8188
rect 38012 8186 38036 8188
rect 38092 8186 38116 8188
rect 38172 8186 38196 8188
rect 38252 8186 38258 8188
rect 38012 8134 38014 8186
rect 38194 8134 38196 8186
rect 37950 8132 37956 8134
rect 38012 8132 38036 8134
rect 38092 8132 38116 8134
rect 38172 8132 38196 8134
rect 38252 8132 38258 8134
rect 37950 8123 38258 8132
rect 38292 7404 38344 7410
rect 38292 7346 38344 7352
rect 37950 7100 38258 7109
rect 37950 7098 37956 7100
rect 38012 7098 38036 7100
rect 38092 7098 38116 7100
rect 38172 7098 38196 7100
rect 38252 7098 38258 7100
rect 38012 7046 38014 7098
rect 38194 7046 38196 7098
rect 37950 7044 37956 7046
rect 38012 7044 38036 7046
rect 38092 7044 38116 7046
rect 38172 7044 38196 7046
rect 38252 7044 38258 7046
rect 37950 7035 38258 7044
rect 38016 6656 38068 6662
rect 38016 6598 38068 6604
rect 38028 6361 38056 6598
rect 38014 6352 38070 6361
rect 38014 6287 38070 6296
rect 37950 6012 38258 6021
rect 37950 6010 37956 6012
rect 38012 6010 38036 6012
rect 38092 6010 38116 6012
rect 38172 6010 38196 6012
rect 38252 6010 38258 6012
rect 38012 5958 38014 6010
rect 38194 5958 38196 6010
rect 37950 5956 37956 5958
rect 38012 5956 38036 5958
rect 38092 5956 38116 5958
rect 38172 5956 38196 5958
rect 38252 5956 38258 5958
rect 37950 5947 38258 5956
rect 37832 5908 37884 5914
rect 37832 5850 37884 5856
rect 37752 5358 37872 5386
rect 37740 5228 37792 5234
rect 37740 5170 37792 5176
rect 37648 4820 37700 4826
rect 37648 4762 37700 4768
rect 37752 134 37780 5170
rect 37844 2514 37872 5358
rect 38200 5228 38252 5234
rect 38200 5170 38252 5176
rect 38212 5030 38240 5170
rect 38200 5024 38252 5030
rect 38200 4966 38252 4972
rect 37950 4924 38258 4933
rect 37950 4922 37956 4924
rect 38012 4922 38036 4924
rect 38092 4922 38116 4924
rect 38172 4922 38196 4924
rect 38252 4922 38258 4924
rect 38012 4870 38014 4922
rect 38194 4870 38196 4922
rect 37950 4868 37956 4870
rect 38012 4868 38036 4870
rect 38092 4868 38116 4870
rect 38172 4868 38196 4870
rect 38252 4868 38258 4870
rect 37950 4859 38258 4868
rect 37950 3836 38258 3845
rect 37950 3834 37956 3836
rect 38012 3834 38036 3836
rect 38092 3834 38116 3836
rect 38172 3834 38196 3836
rect 38252 3834 38258 3836
rect 38012 3782 38014 3834
rect 38194 3782 38196 3834
rect 37950 3780 37956 3782
rect 38012 3780 38036 3782
rect 38092 3780 38116 3782
rect 38172 3780 38196 3782
rect 38252 3780 38258 3782
rect 37950 3771 38258 3780
rect 37950 2748 38258 2757
rect 37950 2746 37956 2748
rect 38012 2746 38036 2748
rect 38092 2746 38116 2748
rect 38172 2746 38196 2748
rect 38252 2746 38258 2748
rect 38012 2694 38014 2746
rect 38194 2694 38196 2746
rect 37950 2692 37956 2694
rect 38012 2692 38036 2694
rect 38092 2692 38116 2694
rect 38172 2692 38196 2694
rect 38252 2692 38258 2694
rect 37950 2683 38258 2692
rect 38304 2650 38332 7346
rect 38396 5370 38424 8910
rect 38580 8566 38608 9250
rect 38568 8560 38620 8566
rect 38568 8502 38620 8508
rect 38658 8528 38714 8537
rect 38658 8463 38714 8472
rect 38752 8492 38804 8498
rect 38672 8090 38700 8463
rect 38752 8434 38804 8440
rect 38844 8492 38896 8498
rect 38844 8434 38896 8440
rect 38660 8084 38712 8090
rect 38660 8026 38712 8032
rect 38568 7268 38620 7274
rect 38568 7210 38620 7216
rect 38580 6905 38608 7210
rect 38566 6896 38622 6905
rect 38566 6831 38622 6840
rect 38476 6792 38528 6798
rect 38476 6734 38528 6740
rect 38488 6458 38516 6734
rect 38660 6656 38712 6662
rect 38660 6598 38712 6604
rect 38476 6452 38528 6458
rect 38476 6394 38528 6400
rect 38672 6361 38700 6598
rect 38658 6352 38714 6361
rect 38658 6287 38714 6296
rect 38476 6248 38528 6254
rect 38476 6190 38528 6196
rect 38384 5364 38436 5370
rect 38384 5306 38436 5312
rect 38488 5250 38516 6190
rect 38568 5704 38620 5710
rect 38568 5646 38620 5652
rect 38396 5222 38516 5250
rect 38396 3738 38424 5222
rect 38476 5024 38528 5030
rect 38476 4966 38528 4972
rect 38384 3732 38436 3738
rect 38384 3674 38436 3680
rect 38488 3466 38516 4966
rect 38476 3460 38528 3466
rect 38476 3402 38528 3408
rect 38292 2644 38344 2650
rect 38292 2586 38344 2592
rect 37832 2508 37884 2514
rect 37832 2450 37884 2456
rect 38108 2440 38160 2446
rect 38108 2382 38160 2388
rect 37924 2304 37976 2310
rect 37924 2246 37976 2252
rect 37936 1737 37964 2246
rect 38120 1902 38148 2382
rect 38292 2304 38344 2310
rect 38292 2246 38344 2252
rect 38108 1896 38160 1902
rect 38108 1838 38160 1844
rect 37922 1728 37978 1737
rect 37922 1663 37978 1672
rect 38304 1465 38332 2246
rect 38290 1456 38346 1465
rect 38290 1391 38346 1400
rect 38580 202 38608 5646
rect 38764 5370 38792 8434
rect 38856 8401 38884 8434
rect 38842 8392 38898 8401
rect 38842 8327 38898 8336
rect 38948 7834 38976 9279
rect 39486 9072 39542 9081
rect 39486 9007 39542 9016
rect 39394 8936 39450 8945
rect 39394 8871 39450 8880
rect 39010 8732 39318 8741
rect 39010 8730 39016 8732
rect 39072 8730 39096 8732
rect 39152 8730 39176 8732
rect 39232 8730 39256 8732
rect 39312 8730 39318 8732
rect 39072 8678 39074 8730
rect 39254 8678 39256 8730
rect 39010 8676 39016 8678
rect 39072 8676 39096 8678
rect 39152 8676 39176 8678
rect 39232 8676 39256 8678
rect 39312 8676 39318 8678
rect 39010 8667 39318 8676
rect 39408 8514 39436 8871
rect 39316 8486 39436 8514
rect 39028 8356 39080 8362
rect 39028 8298 39080 8304
rect 39040 8265 39068 8298
rect 39026 8256 39082 8265
rect 39026 8191 39082 8200
rect 39316 7886 39344 8486
rect 39396 8356 39448 8362
rect 39396 8298 39448 8304
rect 39408 7993 39436 8298
rect 39394 7984 39450 7993
rect 39394 7919 39450 7928
rect 38856 7806 38976 7834
rect 39304 7880 39356 7886
rect 39304 7822 39356 7828
rect 38856 7546 38884 7806
rect 38936 7744 38988 7750
rect 39396 7744 39448 7750
rect 38936 7686 38988 7692
rect 39394 7712 39396 7721
rect 39448 7712 39450 7721
rect 38844 7540 38896 7546
rect 38844 7482 38896 7488
rect 38948 7449 38976 7686
rect 39010 7644 39318 7653
rect 39394 7647 39450 7656
rect 39010 7642 39016 7644
rect 39072 7642 39096 7644
rect 39152 7642 39176 7644
rect 39232 7642 39256 7644
rect 39312 7642 39318 7644
rect 39072 7590 39074 7642
rect 39254 7590 39256 7642
rect 39010 7588 39016 7590
rect 39072 7588 39096 7590
rect 39152 7588 39176 7590
rect 39232 7588 39256 7590
rect 39312 7588 39318 7590
rect 39010 7579 39318 7588
rect 38934 7440 38990 7449
rect 38934 7375 38990 7384
rect 39212 7404 39264 7410
rect 39212 7346 39264 7352
rect 39224 7002 39252 7346
rect 39396 7200 39448 7206
rect 39394 7168 39396 7177
rect 39448 7168 39450 7177
rect 39394 7103 39450 7112
rect 39212 6996 39264 7002
rect 39212 6938 39264 6944
rect 38844 6792 38896 6798
rect 38844 6734 38896 6740
rect 38856 6390 38884 6734
rect 39500 6662 39528 9007
rect 39578 8800 39634 8809
rect 39578 8735 39634 8744
rect 39592 7546 39620 8735
rect 39580 7540 39632 7546
rect 39580 7482 39632 7488
rect 39684 6730 39712 9551
rect 39776 7478 39804 9823
rect 39764 7472 39816 7478
rect 39764 7414 39816 7420
rect 39672 6724 39724 6730
rect 39672 6666 39724 6672
rect 39488 6656 39540 6662
rect 39394 6624 39450 6633
rect 39488 6598 39540 6604
rect 39010 6556 39318 6565
rect 39394 6559 39450 6568
rect 39010 6554 39016 6556
rect 39072 6554 39096 6556
rect 39152 6554 39176 6556
rect 39232 6554 39256 6556
rect 39312 6554 39318 6556
rect 39072 6502 39074 6554
rect 39254 6502 39256 6554
rect 39010 6500 39016 6502
rect 39072 6500 39096 6502
rect 39152 6500 39176 6502
rect 39232 6500 39256 6502
rect 39312 6500 39318 6502
rect 39010 6491 39318 6500
rect 39408 6458 39436 6559
rect 39396 6452 39448 6458
rect 39396 6394 39448 6400
rect 38844 6384 38896 6390
rect 38844 6326 38896 6332
rect 38844 6112 38896 6118
rect 38842 6080 38844 6089
rect 38896 6080 38898 6089
rect 38842 6015 38898 6024
rect 39396 5840 39448 5846
rect 39394 5808 39396 5817
rect 39448 5808 39450 5817
rect 39394 5743 39450 5752
rect 39212 5704 39264 5710
rect 39210 5672 39212 5681
rect 39264 5672 39266 5681
rect 39210 5607 39266 5616
rect 39764 5636 39816 5642
rect 39764 5578 39816 5584
rect 39010 5468 39318 5477
rect 39010 5466 39016 5468
rect 39072 5466 39096 5468
rect 39152 5466 39176 5468
rect 39232 5466 39256 5468
rect 39312 5466 39318 5468
rect 39072 5414 39074 5466
rect 39254 5414 39256 5466
rect 39010 5412 39016 5414
rect 39072 5412 39096 5414
rect 39152 5412 39176 5414
rect 39232 5412 39256 5414
rect 39312 5412 39318 5414
rect 39010 5403 39318 5412
rect 38752 5364 38804 5370
rect 38752 5306 38804 5312
rect 39396 5364 39448 5370
rect 39396 5306 39448 5312
rect 39408 5273 39436 5306
rect 39394 5264 39450 5273
rect 38660 5228 38712 5234
rect 39394 5199 39450 5208
rect 38660 5170 38712 5176
rect 38568 196 38620 202
rect 38568 138 38620 144
rect 37740 128 37792 134
rect 37740 70 37792 76
rect 38672 56 38700 5170
rect 39028 5024 39080 5030
rect 39026 4992 39028 5001
rect 39080 4992 39082 5001
rect 39026 4927 39082 4936
rect 39396 4752 39448 4758
rect 39394 4720 39396 4729
rect 39448 4720 39450 4729
rect 39394 4655 39450 4664
rect 39672 4480 39724 4486
rect 39672 4422 39724 4428
rect 39010 4380 39318 4389
rect 39010 4378 39016 4380
rect 39072 4378 39096 4380
rect 39152 4378 39176 4380
rect 39232 4378 39256 4380
rect 39312 4378 39318 4380
rect 39072 4326 39074 4378
rect 39254 4326 39256 4378
rect 39010 4324 39016 4326
rect 39072 4324 39096 4326
rect 39152 4324 39176 4326
rect 39232 4324 39256 4326
rect 39312 4324 39318 4326
rect 39010 4315 39318 4324
rect 39394 4176 39450 4185
rect 38844 4140 38896 4146
rect 39394 4111 39450 4120
rect 39580 4140 39632 4146
rect 38844 4082 38896 4088
rect 38856 3670 38884 4082
rect 39408 4010 39436 4111
rect 39580 4082 39632 4088
rect 39396 4004 39448 4010
rect 39396 3946 39448 3952
rect 39028 3936 39080 3942
rect 39026 3904 39028 3913
rect 39080 3904 39082 3913
rect 39026 3839 39082 3848
rect 38844 3664 38896 3670
rect 39396 3664 39448 3670
rect 38844 3606 38896 3612
rect 39394 3632 39396 3641
rect 39448 3632 39450 3641
rect 39394 3567 39450 3576
rect 39010 3292 39318 3301
rect 39010 3290 39016 3292
rect 39072 3290 39096 3292
rect 39152 3290 39176 3292
rect 39232 3290 39256 3292
rect 39312 3290 39318 3292
rect 39072 3238 39074 3290
rect 39254 3238 39256 3290
rect 39010 3236 39016 3238
rect 39072 3236 39096 3238
rect 39152 3236 39176 3238
rect 39232 3236 39256 3238
rect 39312 3236 39318 3238
rect 39010 3227 39318 3236
rect 39396 3188 39448 3194
rect 39396 3130 39448 3136
rect 39408 3097 39436 3130
rect 39394 3088 39450 3097
rect 38844 3052 38896 3058
rect 39394 3023 39450 3032
rect 38844 2994 38896 3000
rect 38856 2530 38884 2994
rect 39488 2984 39540 2990
rect 39488 2926 39540 2932
rect 39028 2848 39080 2854
rect 39026 2816 39028 2825
rect 39080 2816 39082 2825
rect 39026 2751 39082 2760
rect 39396 2576 39448 2582
rect 38764 2502 38884 2530
rect 39394 2544 39396 2553
rect 39448 2544 39450 2553
rect 38764 1873 38792 2502
rect 39394 2479 39450 2488
rect 38844 2440 38896 2446
rect 38844 2382 38896 2388
rect 38750 1864 38806 1873
rect 38750 1799 38806 1808
rect 38856 1222 38884 2382
rect 38936 2304 38988 2310
rect 38936 2246 38988 2252
rect 38948 2009 38976 2246
rect 39010 2204 39318 2213
rect 39010 2202 39016 2204
rect 39072 2202 39096 2204
rect 39152 2202 39176 2204
rect 39232 2202 39256 2204
rect 39312 2202 39318 2204
rect 39072 2150 39074 2202
rect 39254 2150 39256 2202
rect 39010 2148 39016 2150
rect 39072 2148 39096 2150
rect 39152 2148 39176 2150
rect 39232 2148 39256 2150
rect 39312 2148 39318 2150
rect 39010 2139 39318 2148
rect 38934 2000 38990 2009
rect 38934 1935 38990 1944
rect 38844 1216 38896 1222
rect 38844 1158 38896 1164
rect 39500 66 39528 2926
rect 39592 1290 39620 4082
rect 39580 1284 39632 1290
rect 39580 1226 39632 1232
rect 39684 1193 39712 4422
rect 39776 4298 39804 5578
rect 39948 5568 40000 5574
rect 39946 5536 39948 5545
rect 40000 5536 40002 5545
rect 39946 5471 40002 5480
rect 39856 4548 39908 4554
rect 39856 4490 39908 4496
rect 39868 4457 39896 4490
rect 39854 4448 39910 4457
rect 39854 4383 39910 4392
rect 39776 4270 39896 4298
rect 39764 2916 39816 2922
rect 39764 2858 39816 2864
rect 39670 1184 39726 1193
rect 39670 1119 39726 1128
rect 39488 60 39540 66
rect 33244 14 33640 42
rect 34242 0 34298 56
rect 35346 0 35402 56
rect 36450 0 36506 56
rect 37554 0 37610 56
rect 38658 0 38714 56
rect 39776 56 39804 2858
rect 39868 1329 39896 4270
rect 39948 3392 40000 3398
rect 39946 3360 39948 3369
rect 40000 3360 40002 3369
rect 39946 3295 40002 3304
rect 39948 2304 40000 2310
rect 39946 2272 39948 2281
rect 40000 2272 40002 2281
rect 39946 2207 40002 2216
rect 39854 1320 39910 1329
rect 39854 1255 39910 1264
rect 39488 2 39540 8
rect 39762 0 39818 56
<< via2 >>
rect 1306 9560 1362 9616
rect 110 9288 166 9344
rect 386 9016 442 9072
rect 202 8744 258 8800
rect 294 6296 350 6352
rect 846 8472 902 8528
rect 754 7656 810 7712
rect 754 7404 810 7440
rect 754 7384 756 7404
rect 756 7384 808 7404
rect 808 7384 810 7404
rect 754 7112 810 7168
rect 478 5752 534 5808
rect 386 4120 442 4176
rect 570 5208 626 5264
rect 1122 8200 1178 8256
rect 1214 7948 1270 7984
rect 1214 7928 1216 7948
rect 1216 7928 1268 7948
rect 1268 7928 1270 7948
rect 1030 6840 1086 6896
rect 938 6568 994 6624
rect 1214 6024 1270 6080
rect 1030 5480 1086 5536
rect 754 3848 810 3904
rect 754 3576 810 3632
rect 1306 4936 1362 4992
rect 1122 4700 1124 4720
rect 1124 4700 1176 4720
rect 1176 4700 1178 4720
rect 1122 4664 1178 4700
rect 1122 4392 1178 4448
rect 570 2760 626 2816
rect 386 1672 442 1728
rect 938 1400 994 1456
rect 1306 2216 1362 2272
rect 2318 9832 2374 9888
rect 1956 8186 2012 8188
rect 2036 8186 2092 8188
rect 2116 8186 2172 8188
rect 2196 8186 2252 8188
rect 1956 8134 2002 8186
rect 2002 8134 2012 8186
rect 2036 8134 2066 8186
rect 2066 8134 2078 8186
rect 2078 8134 2092 8186
rect 2116 8134 2130 8186
rect 2130 8134 2142 8186
rect 2142 8134 2172 8186
rect 2196 8134 2206 8186
rect 2206 8134 2252 8186
rect 1956 8132 2012 8134
rect 2036 8132 2092 8134
rect 2116 8132 2172 8134
rect 2196 8132 2252 8134
rect 1956 7098 2012 7100
rect 2036 7098 2092 7100
rect 2116 7098 2172 7100
rect 2196 7098 2252 7100
rect 1956 7046 2002 7098
rect 2002 7046 2012 7098
rect 2036 7046 2066 7098
rect 2066 7046 2078 7098
rect 2078 7046 2092 7098
rect 2116 7046 2130 7098
rect 2130 7046 2142 7098
rect 2142 7046 2172 7098
rect 2196 7046 2206 7098
rect 2206 7046 2252 7098
rect 1956 7044 2012 7046
rect 2036 7044 2092 7046
rect 2116 7044 2172 7046
rect 2196 7044 2252 7046
rect 2226 6296 2282 6352
rect 1766 5092 1822 5128
rect 1766 5072 1768 5092
rect 1768 5072 1820 5092
rect 1820 5072 1822 5092
rect 2134 6196 2136 6216
rect 2136 6196 2188 6216
rect 2188 6196 2190 6216
rect 2134 6160 2190 6196
rect 1956 6010 2012 6012
rect 2036 6010 2092 6012
rect 2116 6010 2172 6012
rect 2196 6010 2252 6012
rect 1956 5958 2002 6010
rect 2002 5958 2012 6010
rect 2036 5958 2066 6010
rect 2066 5958 2078 6010
rect 2078 5958 2092 6010
rect 2116 5958 2130 6010
rect 2130 5958 2142 6010
rect 2142 5958 2172 6010
rect 2196 5958 2206 6010
rect 2206 5958 2252 6010
rect 1956 5956 2012 5958
rect 2036 5956 2092 5958
rect 2116 5956 2172 5958
rect 2196 5956 2252 5958
rect 2502 9152 2558 9208
rect 2594 8064 2650 8120
rect 2594 7828 2596 7848
rect 2596 7828 2648 7848
rect 2648 7828 2650 7848
rect 2594 7792 2650 7828
rect 1956 4922 2012 4924
rect 2036 4922 2092 4924
rect 2116 4922 2172 4924
rect 2196 4922 2252 4924
rect 1956 4870 2002 4922
rect 2002 4870 2012 4922
rect 2036 4870 2066 4922
rect 2066 4870 2078 4922
rect 2078 4870 2092 4922
rect 2116 4870 2130 4922
rect 2130 4870 2142 4922
rect 2142 4870 2172 4922
rect 2196 4870 2206 4922
rect 2206 4870 2252 4922
rect 1956 4868 2012 4870
rect 2036 4868 2092 4870
rect 2116 4868 2172 4870
rect 2196 4868 2252 4870
rect 2502 6024 2558 6080
rect 2502 5908 2558 5944
rect 2502 5888 2504 5908
rect 2504 5888 2556 5908
rect 2556 5888 2558 5908
rect 2502 5652 2504 5672
rect 2504 5652 2556 5672
rect 2556 5652 2558 5672
rect 2502 5616 2558 5652
rect 2042 4548 2098 4584
rect 2042 4528 2044 4548
rect 2044 4528 2096 4548
rect 2096 4528 2098 4548
rect 2686 6296 2742 6352
rect 3016 8730 3072 8732
rect 3096 8730 3152 8732
rect 3176 8730 3232 8732
rect 3256 8730 3312 8732
rect 3016 8678 3062 8730
rect 3062 8678 3072 8730
rect 3096 8678 3126 8730
rect 3126 8678 3138 8730
rect 3138 8678 3152 8730
rect 3176 8678 3190 8730
rect 3190 8678 3202 8730
rect 3202 8678 3232 8730
rect 3256 8678 3266 8730
rect 3266 8678 3312 8730
rect 3016 8676 3072 8678
rect 3096 8676 3152 8678
rect 3176 8676 3232 8678
rect 3256 8676 3312 8678
rect 3016 7642 3072 7644
rect 3096 7642 3152 7644
rect 3176 7642 3232 7644
rect 3256 7642 3312 7644
rect 3016 7590 3062 7642
rect 3062 7590 3072 7642
rect 3096 7590 3126 7642
rect 3126 7590 3138 7642
rect 3138 7590 3152 7642
rect 3176 7590 3190 7642
rect 3190 7590 3202 7642
rect 3202 7590 3232 7642
rect 3256 7590 3266 7642
rect 3266 7590 3312 7642
rect 3016 7588 3072 7590
rect 3096 7588 3152 7590
rect 3176 7588 3232 7590
rect 3256 7588 3312 7590
rect 3514 9016 3570 9072
rect 3238 6976 3294 7032
rect 3238 6876 3240 6896
rect 3240 6876 3292 6896
rect 3292 6876 3294 6896
rect 3238 6840 3294 6876
rect 3238 6740 3240 6760
rect 3240 6740 3292 6760
rect 3292 6740 3294 6760
rect 3238 6704 3294 6740
rect 3016 6554 3072 6556
rect 3096 6554 3152 6556
rect 3176 6554 3232 6556
rect 3256 6554 3312 6556
rect 3016 6502 3062 6554
rect 3062 6502 3072 6554
rect 3096 6502 3126 6554
rect 3126 6502 3138 6554
rect 3138 6502 3152 6554
rect 3176 6502 3190 6554
rect 3190 6502 3202 6554
rect 3202 6502 3232 6554
rect 3256 6502 3266 6554
rect 3266 6502 3312 6554
rect 3016 6500 3072 6502
rect 3096 6500 3152 6502
rect 3176 6500 3232 6502
rect 3256 6500 3312 6502
rect 3146 5752 3202 5808
rect 4526 10240 4582 10296
rect 4434 9560 4490 9616
rect 3974 7656 4030 7712
rect 3514 5480 3570 5536
rect 3016 5466 3072 5468
rect 3096 5466 3152 5468
rect 3176 5466 3232 5468
rect 3256 5466 3312 5468
rect 3016 5414 3062 5466
rect 3062 5414 3072 5466
rect 3096 5414 3126 5466
rect 3126 5414 3138 5466
rect 3138 5414 3152 5466
rect 3176 5414 3190 5466
rect 3190 5414 3202 5466
rect 3202 5414 3232 5466
rect 3256 5414 3266 5466
rect 3266 5414 3312 5466
rect 3016 5412 3072 5414
rect 3096 5412 3152 5414
rect 3176 5412 3232 5414
rect 3256 5412 3312 5414
rect 3974 5888 4030 5944
rect 3016 4378 3072 4380
rect 3096 4378 3152 4380
rect 3176 4378 3232 4380
rect 3256 4378 3312 4380
rect 3016 4326 3062 4378
rect 3062 4326 3072 4378
rect 3096 4326 3126 4378
rect 3126 4326 3138 4378
rect 3138 4326 3152 4378
rect 3176 4326 3190 4378
rect 3190 4326 3202 4378
rect 3202 4326 3232 4378
rect 3256 4326 3266 4378
rect 3266 4326 3312 4378
rect 3016 4324 3072 4326
rect 3096 4324 3152 4326
rect 3176 4324 3232 4326
rect 3256 4324 3312 4326
rect 2778 4120 2834 4176
rect 1956 3834 2012 3836
rect 2036 3834 2092 3836
rect 2116 3834 2172 3836
rect 2196 3834 2252 3836
rect 1956 3782 2002 3834
rect 2002 3782 2012 3834
rect 2036 3782 2066 3834
rect 2066 3782 2078 3834
rect 2078 3782 2092 3834
rect 2116 3782 2130 3834
rect 2130 3782 2142 3834
rect 2142 3782 2172 3834
rect 2196 3782 2206 3834
rect 2206 3782 2252 3834
rect 1956 3780 2012 3782
rect 2036 3780 2092 3782
rect 2116 3780 2172 3782
rect 2196 3780 2252 3782
rect 1956 2746 2012 2748
rect 2036 2746 2092 2748
rect 2116 2746 2172 2748
rect 2196 2746 2252 2748
rect 1956 2694 2002 2746
rect 2002 2694 2012 2746
rect 2036 2694 2066 2746
rect 2066 2694 2078 2746
rect 2078 2694 2092 2746
rect 2116 2694 2130 2746
rect 2130 2694 2142 2746
rect 2142 2694 2172 2746
rect 2196 2694 2206 2746
rect 2206 2694 2252 2746
rect 1956 2692 2012 2694
rect 2036 2692 2092 2694
rect 2116 2692 2172 2694
rect 2196 2692 2252 2694
rect 1674 2352 1730 2408
rect 2318 1944 2374 2000
rect 2778 3984 2834 4040
rect 3054 3440 3110 3496
rect 2686 3304 2742 3360
rect 2686 3052 2742 3088
rect 2686 3032 2688 3052
rect 2688 3032 2740 3052
rect 2740 3032 2742 3052
rect 3016 3290 3072 3292
rect 3096 3290 3152 3292
rect 3176 3290 3232 3292
rect 3256 3290 3312 3292
rect 3016 3238 3062 3290
rect 3062 3238 3072 3290
rect 3096 3238 3126 3290
rect 3126 3238 3138 3290
rect 3138 3238 3152 3290
rect 3176 3238 3190 3290
rect 3190 3238 3202 3290
rect 3202 3238 3232 3290
rect 3256 3238 3266 3290
rect 3266 3238 3312 3290
rect 3016 3236 3072 3238
rect 3096 3236 3152 3238
rect 3176 3236 3232 3238
rect 3256 3236 3312 3238
rect 4434 7112 4490 7168
rect 4250 6740 4252 6760
rect 4252 6740 4304 6760
rect 4304 6740 4306 6760
rect 4250 6704 4306 6740
rect 4342 5752 4398 5808
rect 2594 2488 2650 2544
rect 3016 2202 3072 2204
rect 3096 2202 3152 2204
rect 3176 2202 3232 2204
rect 3256 2202 3312 2204
rect 3016 2150 3062 2202
rect 3062 2150 3072 2202
rect 3096 2150 3126 2202
rect 3126 2150 3138 2202
rect 3138 2150 3152 2202
rect 3176 2150 3190 2202
rect 3190 2150 3202 2202
rect 3202 2150 3232 2202
rect 3256 2150 3266 2202
rect 3266 2150 3312 2202
rect 3016 2148 3072 2150
rect 3096 2148 3152 2150
rect 3176 2148 3232 2150
rect 3256 2148 3312 2150
rect 2594 584 2650 640
rect 4342 3612 4344 3632
rect 4344 3612 4396 3632
rect 4396 3612 4398 3632
rect 4342 3576 4398 3612
rect 4066 2916 4122 2952
rect 4066 2896 4068 2916
rect 4068 2896 4120 2916
rect 4120 2896 4122 2916
rect 4710 10648 4766 10704
rect 4066 1808 4122 1864
rect 3974 720 4030 776
rect 4986 10512 5042 10568
rect 5262 10376 5318 10432
rect 4894 6568 4950 6624
rect 5170 7384 5226 7440
rect 5170 6432 5226 6488
rect 5446 6568 5502 6624
rect 5446 6432 5502 6488
rect 5630 6840 5686 6896
rect 5354 5752 5410 5808
rect 5354 3848 5410 3904
rect 4894 3032 4950 3088
rect 4894 2488 4950 2544
rect 4618 1264 4674 1320
rect 5814 8880 5870 8936
rect 5814 6432 5870 6488
rect 6366 7384 6422 7440
rect 6734 8744 6790 8800
rect 7010 7928 7066 7984
rect 6918 7792 6974 7848
rect 6366 5480 6422 5536
rect 6182 4120 6238 4176
rect 6826 6976 6882 7032
rect 7010 7248 7066 7304
rect 6826 6296 6882 6352
rect 6642 5208 6698 5264
rect 6642 3612 6644 3632
rect 6644 3612 6696 3632
rect 6696 3612 6698 3632
rect 6642 3576 6698 3612
rect 5630 448 5686 504
rect 7194 8336 7250 8392
rect 7010 5364 7066 5400
rect 7010 5344 7012 5364
rect 7012 5344 7064 5364
rect 7064 5344 7066 5364
rect 6826 3188 6882 3224
rect 6826 3168 6828 3188
rect 6828 3168 6880 3188
rect 6880 3168 6882 3188
rect 7286 6024 7342 6080
rect 7562 9832 7618 9888
rect 7654 9424 7710 9480
rect 7746 8200 7802 8256
rect 7654 8064 7710 8120
rect 7102 1944 7158 2000
rect 7470 3712 7526 3768
rect 8206 10240 8262 10296
rect 7930 9696 7986 9752
rect 8022 8472 8078 8528
rect 7956 8186 8012 8188
rect 8036 8186 8092 8188
rect 8116 8186 8172 8188
rect 8196 8186 8252 8188
rect 7956 8134 8002 8186
rect 8002 8134 8012 8186
rect 8036 8134 8066 8186
rect 8066 8134 8078 8186
rect 8078 8134 8092 8186
rect 8116 8134 8130 8186
rect 8130 8134 8142 8186
rect 8142 8134 8172 8186
rect 8196 8134 8206 8186
rect 8206 8134 8252 8186
rect 7956 8132 8012 8134
rect 8036 8132 8092 8134
rect 8116 8132 8172 8134
rect 8196 8132 8252 8134
rect 7930 7384 7986 7440
rect 8390 8236 8392 8256
rect 8392 8236 8444 8256
rect 8444 8236 8446 8256
rect 8390 8200 8446 8236
rect 9310 10376 9366 10432
rect 9402 10240 9458 10296
rect 9402 8744 9458 8800
rect 9016 8730 9072 8732
rect 9096 8730 9152 8732
rect 9176 8730 9232 8732
rect 9256 8730 9312 8732
rect 9016 8678 9062 8730
rect 9062 8678 9072 8730
rect 9096 8678 9126 8730
rect 9126 8678 9138 8730
rect 9138 8678 9152 8730
rect 9176 8678 9190 8730
rect 9190 8678 9202 8730
rect 9202 8678 9232 8730
rect 9256 8678 9266 8730
rect 9266 8678 9312 8730
rect 9016 8676 9072 8678
rect 9096 8676 9152 8678
rect 9176 8676 9232 8678
rect 9256 8676 9312 8678
rect 10046 10648 10102 10704
rect 9862 9832 9918 9888
rect 10046 9832 10102 9888
rect 8666 8200 8722 8256
rect 8574 7928 8630 7984
rect 8574 7656 8630 7712
rect 8666 7520 8722 7576
rect 9016 7642 9072 7644
rect 9096 7642 9152 7644
rect 9176 7642 9232 7644
rect 9256 7642 9312 7644
rect 9016 7590 9062 7642
rect 9062 7590 9072 7642
rect 9096 7590 9126 7642
rect 9126 7590 9138 7642
rect 9138 7590 9152 7642
rect 9176 7590 9190 7642
rect 9190 7590 9202 7642
rect 9202 7590 9232 7642
rect 9256 7590 9266 7642
rect 9266 7590 9312 7642
rect 9016 7588 9072 7590
rect 9096 7588 9152 7590
rect 9176 7588 9232 7590
rect 9256 7588 9312 7590
rect 8482 7248 8538 7304
rect 7956 7098 8012 7100
rect 8036 7098 8092 7100
rect 8116 7098 8172 7100
rect 8196 7098 8252 7100
rect 7956 7046 8002 7098
rect 8002 7046 8012 7098
rect 8036 7046 8066 7098
rect 8066 7046 8078 7098
rect 8078 7046 8092 7098
rect 8116 7046 8130 7098
rect 8130 7046 8142 7098
rect 8142 7046 8172 7098
rect 8196 7046 8206 7098
rect 8206 7046 8252 7098
rect 7956 7044 8012 7046
rect 8036 7044 8092 7046
rect 8116 7044 8172 7046
rect 8196 7044 8252 7046
rect 7956 6010 8012 6012
rect 8036 6010 8092 6012
rect 8116 6010 8172 6012
rect 8196 6010 8252 6012
rect 7956 5958 8002 6010
rect 8002 5958 8012 6010
rect 8036 5958 8066 6010
rect 8066 5958 8078 6010
rect 8078 5958 8092 6010
rect 8116 5958 8130 6010
rect 8130 5958 8142 6010
rect 8142 5958 8172 6010
rect 8196 5958 8206 6010
rect 8206 5958 8252 6010
rect 7956 5956 8012 5958
rect 8036 5956 8092 5958
rect 8116 5956 8172 5958
rect 8196 5956 8252 5958
rect 8482 6840 8538 6896
rect 8482 6568 8538 6624
rect 7956 4922 8012 4924
rect 8036 4922 8092 4924
rect 8116 4922 8172 4924
rect 8196 4922 8252 4924
rect 7956 4870 8002 4922
rect 8002 4870 8012 4922
rect 8036 4870 8066 4922
rect 8066 4870 8078 4922
rect 8078 4870 8092 4922
rect 8116 4870 8130 4922
rect 8130 4870 8142 4922
rect 8142 4870 8172 4922
rect 8196 4870 8206 4922
rect 8206 4870 8252 4922
rect 7956 4868 8012 4870
rect 8036 4868 8092 4870
rect 8116 4868 8172 4870
rect 8196 4868 8252 4870
rect 7746 4700 7748 4720
rect 7748 4700 7800 4720
rect 7800 4700 7802 4720
rect 7746 4664 7802 4700
rect 8390 5344 8446 5400
rect 8482 4800 8538 4856
rect 8758 6452 8814 6488
rect 8758 6432 8760 6452
rect 8760 6432 8812 6452
rect 8812 6432 8814 6452
rect 7956 3834 8012 3836
rect 8036 3834 8092 3836
rect 8116 3834 8172 3836
rect 8196 3834 8252 3836
rect 7956 3782 8002 3834
rect 8002 3782 8012 3834
rect 8036 3782 8066 3834
rect 8066 3782 8078 3834
rect 8078 3782 8092 3834
rect 8116 3782 8130 3834
rect 8130 3782 8142 3834
rect 8142 3782 8172 3834
rect 8196 3782 8206 3834
rect 8206 3782 8252 3834
rect 7956 3780 8012 3782
rect 8036 3780 8092 3782
rect 8116 3780 8172 3782
rect 8196 3780 8252 3782
rect 9016 6554 9072 6556
rect 9096 6554 9152 6556
rect 9176 6554 9232 6556
rect 9256 6554 9312 6556
rect 9016 6502 9062 6554
rect 9062 6502 9072 6554
rect 9096 6502 9126 6554
rect 9126 6502 9138 6554
rect 9138 6502 9152 6554
rect 9176 6502 9190 6554
rect 9190 6502 9202 6554
rect 9202 6502 9232 6554
rect 9256 6502 9266 6554
rect 9266 6502 9312 6554
rect 9016 6500 9072 6502
rect 9096 6500 9152 6502
rect 9176 6500 9232 6502
rect 9256 6500 9312 6502
rect 9586 6316 9642 6352
rect 9586 6296 9588 6316
rect 9588 6296 9640 6316
rect 9640 6296 9642 6316
rect 9126 6024 9182 6080
rect 9494 6024 9550 6080
rect 9016 5466 9072 5468
rect 9096 5466 9152 5468
rect 9176 5466 9232 5468
rect 9256 5466 9312 5468
rect 9016 5414 9062 5466
rect 9062 5414 9072 5466
rect 9096 5414 9126 5466
rect 9126 5414 9138 5466
rect 9138 5414 9152 5466
rect 9176 5414 9190 5466
rect 9190 5414 9202 5466
rect 9202 5414 9232 5466
rect 9256 5414 9266 5466
rect 9266 5414 9312 5466
rect 9016 5412 9072 5414
rect 9096 5412 9152 5414
rect 9176 5412 9232 5414
rect 9256 5412 9312 5414
rect 9494 4820 9550 4856
rect 9494 4800 9496 4820
rect 9496 4800 9548 4820
rect 9548 4800 9550 4820
rect 9016 4378 9072 4380
rect 9096 4378 9152 4380
rect 9176 4378 9232 4380
rect 9256 4378 9312 4380
rect 9016 4326 9062 4378
rect 9062 4326 9072 4378
rect 9096 4326 9126 4378
rect 9126 4326 9138 4378
rect 9138 4326 9152 4378
rect 9176 4326 9190 4378
rect 9190 4326 9202 4378
rect 9202 4326 9232 4378
rect 9256 4326 9266 4378
rect 9266 4326 9312 4378
rect 9016 4324 9072 4326
rect 9096 4324 9152 4326
rect 9176 4324 9232 4326
rect 9256 4324 9312 4326
rect 8850 3848 8906 3904
rect 7654 3304 7710 3360
rect 8482 3304 8538 3360
rect 7956 2746 8012 2748
rect 8036 2746 8092 2748
rect 8116 2746 8172 2748
rect 8196 2746 8252 2748
rect 7956 2694 8002 2746
rect 8002 2694 8012 2746
rect 8036 2694 8066 2746
rect 8066 2694 8078 2746
rect 8078 2694 8092 2746
rect 8116 2694 8130 2746
rect 8130 2694 8142 2746
rect 8142 2694 8172 2746
rect 8196 2694 8206 2746
rect 8206 2694 8252 2746
rect 7956 2692 8012 2694
rect 8036 2692 8092 2694
rect 8116 2692 8172 2694
rect 8196 2692 8252 2694
rect 9402 3848 9458 3904
rect 9310 3576 9366 3632
rect 9586 3884 9588 3904
rect 9588 3884 9640 3904
rect 9640 3884 9642 3904
rect 9586 3848 9642 3884
rect 10138 9016 10194 9072
rect 10322 7520 10378 7576
rect 9954 4392 10010 4448
rect 10690 10512 10746 10568
rect 10874 10512 10930 10568
rect 10506 9324 10508 9344
rect 10508 9324 10560 9344
rect 10560 9324 10562 9344
rect 10506 9288 10562 9324
rect 10598 8608 10654 8664
rect 11242 10240 11298 10296
rect 10966 8880 11022 8936
rect 10230 4800 10286 4856
rect 10506 4936 10562 4992
rect 9770 3576 9826 3632
rect 9954 3440 10010 3496
rect 9016 3290 9072 3292
rect 9096 3290 9152 3292
rect 9176 3290 9232 3292
rect 9256 3290 9312 3292
rect 9016 3238 9062 3290
rect 9062 3238 9072 3290
rect 9096 3238 9126 3290
rect 9126 3238 9138 3290
rect 9138 3238 9152 3290
rect 9176 3238 9190 3290
rect 9190 3238 9202 3290
rect 9202 3238 9232 3290
rect 9256 3238 9266 3290
rect 9266 3238 9312 3290
rect 9016 3236 9072 3238
rect 9096 3236 9152 3238
rect 9176 3236 9232 3238
rect 9256 3236 9312 3238
rect 8850 3168 8906 3224
rect 9402 3168 9458 3224
rect 8666 2624 8722 2680
rect 9016 2202 9072 2204
rect 9096 2202 9152 2204
rect 9176 2202 9232 2204
rect 9256 2202 9312 2204
rect 9016 2150 9062 2202
rect 9062 2150 9072 2202
rect 9096 2150 9126 2202
rect 9126 2150 9138 2202
rect 9138 2150 9152 2202
rect 9176 2150 9190 2202
rect 9190 2150 9202 2202
rect 9202 2150 9232 2202
rect 9256 2150 9266 2202
rect 9266 2150 9312 2202
rect 9016 2148 9072 2150
rect 9096 2148 9152 2150
rect 9176 2148 9232 2150
rect 9256 2148 9312 2150
rect 9586 1536 9642 1592
rect 10874 8200 10930 8256
rect 10322 2216 10378 2272
rect 10598 2760 10654 2816
rect 10506 2080 10562 2136
rect 10782 4256 10838 4312
rect 11242 6840 11298 6896
rect 11426 6024 11482 6080
rect 12530 8064 12586 8120
rect 12346 6976 12402 7032
rect 11242 4392 11298 4448
rect 10874 2760 10930 2816
rect 11058 2796 11060 2816
rect 11060 2796 11112 2816
rect 11112 2796 11114 2816
rect 11058 2760 11114 2796
rect 11150 2624 11206 2680
rect 11426 4392 11482 4448
rect 12714 7656 12770 7712
rect 12622 4800 12678 4856
rect 12530 4120 12586 4176
rect 12254 3032 12310 3088
rect 12162 2624 12218 2680
rect 11886 2488 11942 2544
rect 11150 1536 11206 1592
rect 12714 3440 12770 3496
rect 13450 10240 13506 10296
rect 13174 9696 13230 9752
rect 12898 6160 12954 6216
rect 13174 7112 13230 7168
rect 13174 6568 13230 6624
rect 13542 8336 13598 8392
rect 13634 7928 13690 7984
rect 13358 6160 13414 6216
rect 13358 5616 13414 5672
rect 13266 5344 13322 5400
rect 13726 7692 13728 7712
rect 13728 7692 13780 7712
rect 13780 7692 13782 7712
rect 13726 7656 13782 7692
rect 13956 8186 14012 8188
rect 14036 8186 14092 8188
rect 14116 8186 14172 8188
rect 14196 8186 14252 8188
rect 13956 8134 14002 8186
rect 14002 8134 14012 8186
rect 14036 8134 14066 8186
rect 14066 8134 14078 8186
rect 14078 8134 14092 8186
rect 14116 8134 14130 8186
rect 14130 8134 14142 8186
rect 14142 8134 14172 8186
rect 14196 8134 14206 8186
rect 14206 8134 14252 8186
rect 13956 8132 14012 8134
rect 14036 8132 14092 8134
rect 14116 8132 14172 8134
rect 14196 8132 14252 8134
rect 14830 9696 14886 9752
rect 14370 8608 14426 8664
rect 14738 8608 14794 8664
rect 13634 6876 13636 6896
rect 13636 6876 13688 6896
rect 13688 6876 13690 6896
rect 13634 6840 13690 6876
rect 13956 7098 14012 7100
rect 14036 7098 14092 7100
rect 14116 7098 14172 7100
rect 14196 7098 14252 7100
rect 13956 7046 14002 7098
rect 14002 7046 14012 7098
rect 14036 7046 14066 7098
rect 14066 7046 14078 7098
rect 14078 7046 14092 7098
rect 14116 7046 14130 7098
rect 14130 7046 14142 7098
rect 14142 7046 14172 7098
rect 14196 7046 14206 7098
rect 14206 7046 14252 7098
rect 13956 7044 14012 7046
rect 14036 7044 14092 7046
rect 14116 7044 14172 7046
rect 14196 7044 14252 7046
rect 13956 6010 14012 6012
rect 14036 6010 14092 6012
rect 14116 6010 14172 6012
rect 14196 6010 14252 6012
rect 13956 5958 14002 6010
rect 14002 5958 14012 6010
rect 14036 5958 14066 6010
rect 14066 5958 14078 6010
rect 14078 5958 14092 6010
rect 14116 5958 14130 6010
rect 14130 5958 14142 6010
rect 14142 5958 14172 6010
rect 14196 5958 14206 6010
rect 14206 5958 14252 6010
rect 13956 5956 14012 5958
rect 14036 5956 14092 5958
rect 14116 5956 14172 5958
rect 14196 5956 14252 5958
rect 13956 4922 14012 4924
rect 14036 4922 14092 4924
rect 14116 4922 14172 4924
rect 14196 4922 14252 4924
rect 13956 4870 14002 4922
rect 14002 4870 14012 4922
rect 14036 4870 14066 4922
rect 14066 4870 14078 4922
rect 14078 4870 14092 4922
rect 14116 4870 14130 4922
rect 14130 4870 14142 4922
rect 14142 4870 14172 4922
rect 14196 4870 14206 4922
rect 14206 4870 14252 4922
rect 13956 4868 14012 4870
rect 14036 4868 14092 4870
rect 14116 4868 14172 4870
rect 14196 4868 14252 4870
rect 15198 9016 15254 9072
rect 15016 8730 15072 8732
rect 15096 8730 15152 8732
rect 15176 8730 15232 8732
rect 15256 8730 15312 8732
rect 15016 8678 15062 8730
rect 15062 8678 15072 8730
rect 15096 8678 15126 8730
rect 15126 8678 15138 8730
rect 15138 8678 15152 8730
rect 15176 8678 15190 8730
rect 15190 8678 15202 8730
rect 15202 8678 15232 8730
rect 15256 8678 15266 8730
rect 15266 8678 15312 8730
rect 15016 8676 15072 8678
rect 15096 8676 15152 8678
rect 15176 8676 15232 8678
rect 15256 8676 15312 8678
rect 15566 9288 15622 9344
rect 15750 9424 15806 9480
rect 16118 10240 16174 10296
rect 14738 8200 14794 8256
rect 14554 7928 14610 7984
rect 14554 7384 14610 7440
rect 14462 6024 14518 6080
rect 14554 5616 14610 5672
rect 13174 3168 13230 3224
rect 12898 3052 12954 3088
rect 12898 3032 12900 3052
rect 12900 3032 12952 3052
rect 12952 3032 12954 3052
rect 13634 3440 13690 3496
rect 13956 3834 14012 3836
rect 14036 3834 14092 3836
rect 14116 3834 14172 3836
rect 14196 3834 14252 3836
rect 13956 3782 14002 3834
rect 14002 3782 14012 3834
rect 14036 3782 14066 3834
rect 14066 3782 14078 3834
rect 14078 3782 14092 3834
rect 14116 3782 14130 3834
rect 14130 3782 14142 3834
rect 14142 3782 14172 3834
rect 14196 3782 14206 3834
rect 14206 3782 14252 3834
rect 13956 3780 14012 3782
rect 14036 3780 14092 3782
rect 14116 3780 14172 3782
rect 14196 3780 14252 3782
rect 14002 3440 14058 3496
rect 13542 2760 13598 2816
rect 14002 3032 14058 3088
rect 14830 8064 14886 8120
rect 14830 7656 14886 7712
rect 15658 8064 15714 8120
rect 15016 7642 15072 7644
rect 15096 7642 15152 7644
rect 15176 7642 15232 7644
rect 15256 7642 15312 7644
rect 15016 7590 15062 7642
rect 15062 7590 15072 7642
rect 15096 7590 15126 7642
rect 15126 7590 15138 7642
rect 15138 7590 15152 7642
rect 15176 7590 15190 7642
rect 15190 7590 15202 7642
rect 15202 7590 15232 7642
rect 15256 7590 15266 7642
rect 15266 7590 15312 7642
rect 15016 7588 15072 7590
rect 15096 7588 15152 7590
rect 15176 7588 15232 7590
rect 15256 7588 15312 7590
rect 15016 6554 15072 6556
rect 15096 6554 15152 6556
rect 15176 6554 15232 6556
rect 15256 6554 15312 6556
rect 15016 6502 15062 6554
rect 15062 6502 15072 6554
rect 15096 6502 15126 6554
rect 15126 6502 15138 6554
rect 15138 6502 15152 6554
rect 15176 6502 15190 6554
rect 15190 6502 15202 6554
rect 15202 6502 15232 6554
rect 15256 6502 15266 6554
rect 15266 6502 15312 6554
rect 15016 6500 15072 6502
rect 15096 6500 15152 6502
rect 15176 6500 15232 6502
rect 15256 6500 15312 6502
rect 14830 5888 14886 5944
rect 14830 4936 14886 4992
rect 15016 5466 15072 5468
rect 15096 5466 15152 5468
rect 15176 5466 15232 5468
rect 15256 5466 15312 5468
rect 15016 5414 15062 5466
rect 15062 5414 15072 5466
rect 15096 5414 15126 5466
rect 15126 5414 15138 5466
rect 15138 5414 15152 5466
rect 15176 5414 15190 5466
rect 15190 5414 15202 5466
rect 15202 5414 15232 5466
rect 15256 5414 15266 5466
rect 15266 5414 15312 5466
rect 15016 5412 15072 5414
rect 15096 5412 15152 5414
rect 15176 5412 15232 5414
rect 15256 5412 15312 5414
rect 16026 7656 16082 7712
rect 15934 7384 15990 7440
rect 15658 5652 15660 5672
rect 15660 5652 15712 5672
rect 15712 5652 15714 5672
rect 15658 5616 15714 5652
rect 15750 5480 15806 5536
rect 14738 4392 14794 4448
rect 15016 4378 15072 4380
rect 15096 4378 15152 4380
rect 15176 4378 15232 4380
rect 15256 4378 15312 4380
rect 15016 4326 15062 4378
rect 15062 4326 15072 4378
rect 15096 4326 15126 4378
rect 15126 4326 15138 4378
rect 15138 4326 15152 4378
rect 15176 4326 15190 4378
rect 15190 4326 15202 4378
rect 15202 4326 15232 4378
rect 15256 4326 15266 4378
rect 15266 4326 15312 4378
rect 15016 4324 15072 4326
rect 15096 4324 15152 4326
rect 15176 4324 15232 4326
rect 15256 4324 15312 4326
rect 15382 4120 15438 4176
rect 14830 3848 14886 3904
rect 14830 3168 14886 3224
rect 14370 2760 14426 2816
rect 13956 2746 14012 2748
rect 14036 2746 14092 2748
rect 14116 2746 14172 2748
rect 14196 2746 14252 2748
rect 13956 2694 14002 2746
rect 14002 2694 14012 2746
rect 14036 2694 14066 2746
rect 14066 2694 14078 2746
rect 14078 2694 14092 2746
rect 14116 2694 14130 2746
rect 14130 2694 14142 2746
rect 14142 2694 14172 2746
rect 14196 2694 14206 2746
rect 14206 2694 14252 2746
rect 13956 2692 14012 2694
rect 14036 2692 14092 2694
rect 14116 2692 14172 2694
rect 14196 2692 14252 2694
rect 15750 4936 15806 4992
rect 15016 3290 15072 3292
rect 15096 3290 15152 3292
rect 15176 3290 15232 3292
rect 15256 3290 15312 3292
rect 15016 3238 15062 3290
rect 15062 3238 15072 3290
rect 15096 3238 15126 3290
rect 15126 3238 15138 3290
rect 15138 3238 15152 3290
rect 15176 3238 15190 3290
rect 15190 3238 15202 3290
rect 15202 3238 15232 3290
rect 15256 3238 15266 3290
rect 15266 3238 15312 3290
rect 15016 3236 15072 3238
rect 15096 3236 15152 3238
rect 15176 3236 15232 3238
rect 15256 3236 15312 3238
rect 14554 2488 14610 2544
rect 14278 2216 14334 2272
rect 15658 4120 15714 4176
rect 15658 3712 15714 3768
rect 15016 2202 15072 2204
rect 15096 2202 15152 2204
rect 15176 2202 15232 2204
rect 15256 2202 15312 2204
rect 15016 2150 15062 2202
rect 15062 2150 15072 2202
rect 15096 2150 15126 2202
rect 15126 2150 15138 2202
rect 15138 2150 15152 2202
rect 15176 2150 15190 2202
rect 15190 2150 15202 2202
rect 15202 2150 15232 2202
rect 15256 2150 15266 2202
rect 15266 2150 15312 2202
rect 15016 2148 15072 2150
rect 15096 2148 15152 2150
rect 15176 2148 15232 2150
rect 15256 2148 15312 2150
rect 14646 2080 14702 2136
rect 16026 7148 16028 7168
rect 16028 7148 16080 7168
rect 16080 7148 16082 7168
rect 16026 7112 16082 7148
rect 15934 6976 15990 7032
rect 16026 6432 16082 6488
rect 16302 8064 16358 8120
rect 16670 7656 16726 7712
rect 16486 6296 16542 6352
rect 16670 6840 16726 6896
rect 16670 6568 16726 6624
rect 16026 4140 16082 4176
rect 16026 4120 16028 4140
rect 16028 4120 16080 4140
rect 16080 4120 16082 4140
rect 16210 3440 16266 3496
rect 16118 3304 16174 3360
rect 17038 8472 17094 8528
rect 17406 10240 17462 10296
rect 17406 9832 17462 9888
rect 17406 6840 17462 6896
rect 17682 10512 17738 10568
rect 17682 9832 17738 9888
rect 17958 8880 18014 8936
rect 16854 5208 16910 5264
rect 17130 5616 17186 5672
rect 17590 6432 17646 6488
rect 17498 6296 17554 6352
rect 17314 5208 17370 5264
rect 16486 2488 16542 2544
rect 18050 8336 18106 8392
rect 18326 8744 18382 8800
rect 17958 8064 18014 8120
rect 18142 8064 18198 8120
rect 17958 7692 17960 7712
rect 17960 7692 18012 7712
rect 18012 7692 18014 7712
rect 17958 7656 18014 7692
rect 17866 6568 17922 6624
rect 17498 4120 17554 4176
rect 17498 3168 17554 3224
rect 17498 1400 17554 1456
rect 18326 6568 18382 6624
rect 18142 6296 18198 6352
rect 18142 6024 18198 6080
rect 18142 5208 18198 5264
rect 17866 1672 17922 1728
rect 18694 8608 18750 8664
rect 18510 7112 18566 7168
rect 18510 6876 18512 6896
rect 18512 6876 18564 6896
rect 18564 6876 18566 6896
rect 18510 6840 18566 6876
rect 18510 6704 18566 6760
rect 18602 6568 18658 6624
rect 18602 6024 18658 6080
rect 18234 3712 18290 3768
rect 18878 8064 18934 8120
rect 19062 8064 19118 8120
rect 18786 6976 18842 7032
rect 18694 5208 18750 5264
rect 19062 6876 19064 6896
rect 19064 6876 19116 6896
rect 19116 6876 19118 6896
rect 19062 6840 19118 6876
rect 19062 6432 19118 6488
rect 19522 9696 19578 9752
rect 19430 8200 19486 8256
rect 19246 6060 19248 6080
rect 19248 6060 19300 6080
rect 19300 6060 19302 6080
rect 19246 6024 19302 6060
rect 19430 5888 19486 5944
rect 19338 5208 19394 5264
rect 18694 3440 18750 3496
rect 18878 3440 18934 3496
rect 18786 3168 18842 3224
rect 18694 2896 18750 2952
rect 18510 2624 18566 2680
rect 19154 3304 19210 3360
rect 19956 8186 20012 8188
rect 20036 8186 20092 8188
rect 20116 8186 20172 8188
rect 20196 8186 20252 8188
rect 19956 8134 20002 8186
rect 20002 8134 20012 8186
rect 20036 8134 20066 8186
rect 20066 8134 20078 8186
rect 20078 8134 20092 8186
rect 20116 8134 20130 8186
rect 20130 8134 20142 8186
rect 20142 8134 20172 8186
rect 20196 8134 20206 8186
rect 20206 8134 20252 8186
rect 19956 8132 20012 8134
rect 20036 8132 20092 8134
rect 20116 8132 20172 8134
rect 20196 8132 20252 8134
rect 19246 2352 19302 2408
rect 19430 2896 19486 2952
rect 19338 1944 19394 2000
rect 19956 7098 20012 7100
rect 20036 7098 20092 7100
rect 20116 7098 20172 7100
rect 20196 7098 20252 7100
rect 19956 7046 20002 7098
rect 20002 7046 20012 7098
rect 20036 7046 20066 7098
rect 20066 7046 20078 7098
rect 20078 7046 20092 7098
rect 20116 7046 20130 7098
rect 20130 7046 20142 7098
rect 20142 7046 20172 7098
rect 20196 7046 20206 7098
rect 20206 7046 20252 7098
rect 19956 7044 20012 7046
rect 20036 7044 20092 7046
rect 20116 7044 20172 7046
rect 20196 7044 20252 7046
rect 20442 6840 20498 6896
rect 20350 6024 20406 6080
rect 19956 6010 20012 6012
rect 20036 6010 20092 6012
rect 20116 6010 20172 6012
rect 20196 6010 20252 6012
rect 19956 5958 20002 6010
rect 20002 5958 20012 6010
rect 20036 5958 20066 6010
rect 20066 5958 20078 6010
rect 20078 5958 20092 6010
rect 20116 5958 20130 6010
rect 20130 5958 20142 6010
rect 20142 5958 20172 6010
rect 20196 5958 20206 6010
rect 20206 5958 20252 6010
rect 19956 5956 20012 5958
rect 20036 5956 20092 5958
rect 20116 5956 20172 5958
rect 20196 5956 20252 5958
rect 19956 4922 20012 4924
rect 20036 4922 20092 4924
rect 20116 4922 20172 4924
rect 20196 4922 20252 4924
rect 19956 4870 20002 4922
rect 20002 4870 20012 4922
rect 20036 4870 20066 4922
rect 20066 4870 20078 4922
rect 20078 4870 20092 4922
rect 20116 4870 20130 4922
rect 20130 4870 20142 4922
rect 20142 4870 20172 4922
rect 20196 4870 20206 4922
rect 20206 4870 20252 4922
rect 19956 4868 20012 4870
rect 20036 4868 20092 4870
rect 20116 4868 20172 4870
rect 20196 4868 20252 4870
rect 21016 8730 21072 8732
rect 21096 8730 21152 8732
rect 21176 8730 21232 8732
rect 21256 8730 21312 8732
rect 21016 8678 21062 8730
rect 21062 8678 21072 8730
rect 21096 8678 21126 8730
rect 21126 8678 21138 8730
rect 21138 8678 21152 8730
rect 21176 8678 21190 8730
rect 21190 8678 21202 8730
rect 21202 8678 21232 8730
rect 21256 8678 21266 8730
rect 21266 8678 21312 8730
rect 21016 8676 21072 8678
rect 21096 8676 21152 8678
rect 21176 8676 21232 8678
rect 21256 8676 21312 8678
rect 20810 7656 20866 7712
rect 20718 7520 20774 7576
rect 20718 7248 20774 7304
rect 20810 7112 20866 7168
rect 20626 5888 20682 5944
rect 20626 5616 20682 5672
rect 19956 3834 20012 3836
rect 20036 3834 20092 3836
rect 20116 3834 20172 3836
rect 20196 3834 20252 3836
rect 19956 3782 20002 3834
rect 20002 3782 20012 3834
rect 20036 3782 20066 3834
rect 20066 3782 20078 3834
rect 20078 3782 20092 3834
rect 20116 3782 20130 3834
rect 20130 3782 20142 3834
rect 20142 3782 20172 3834
rect 20196 3782 20206 3834
rect 20206 3782 20252 3834
rect 19956 3780 20012 3782
rect 20036 3780 20092 3782
rect 20116 3780 20172 3782
rect 20196 3780 20252 3782
rect 20350 2760 20406 2816
rect 19956 2746 20012 2748
rect 20036 2746 20092 2748
rect 20116 2746 20172 2748
rect 20196 2746 20252 2748
rect 19956 2694 20002 2746
rect 20002 2694 20012 2746
rect 20036 2694 20066 2746
rect 20066 2694 20078 2746
rect 20078 2694 20092 2746
rect 20116 2694 20130 2746
rect 20130 2694 20142 2746
rect 20142 2694 20172 2746
rect 20196 2694 20206 2746
rect 20206 2694 20252 2746
rect 19956 2692 20012 2694
rect 20036 2692 20092 2694
rect 20116 2692 20172 2694
rect 20196 2692 20252 2694
rect 19798 1808 19854 1864
rect 20994 7928 21050 7984
rect 21016 7642 21072 7644
rect 21096 7642 21152 7644
rect 21176 7642 21232 7644
rect 21256 7642 21312 7644
rect 21016 7590 21062 7642
rect 21062 7590 21072 7642
rect 21096 7590 21126 7642
rect 21126 7590 21138 7642
rect 21138 7590 21152 7642
rect 21176 7590 21190 7642
rect 21190 7590 21202 7642
rect 21202 7590 21232 7642
rect 21256 7590 21266 7642
rect 21266 7590 21312 7642
rect 21016 7588 21072 7590
rect 21096 7588 21152 7590
rect 21176 7588 21232 7590
rect 21256 7588 21312 7590
rect 21454 7520 21510 7576
rect 21016 6554 21072 6556
rect 21096 6554 21152 6556
rect 21176 6554 21232 6556
rect 21256 6554 21312 6556
rect 21016 6502 21062 6554
rect 21062 6502 21072 6554
rect 21096 6502 21126 6554
rect 21126 6502 21138 6554
rect 21138 6502 21152 6554
rect 21176 6502 21190 6554
rect 21190 6502 21202 6554
rect 21202 6502 21232 6554
rect 21256 6502 21266 6554
rect 21266 6502 21312 6554
rect 21016 6500 21072 6502
rect 21096 6500 21152 6502
rect 21176 6500 21232 6502
rect 21256 6500 21312 6502
rect 21822 9152 21878 9208
rect 21016 5466 21072 5468
rect 21096 5466 21152 5468
rect 21176 5466 21232 5468
rect 21256 5466 21312 5468
rect 21016 5414 21062 5466
rect 21062 5414 21072 5466
rect 21096 5414 21126 5466
rect 21126 5414 21138 5466
rect 21138 5414 21152 5466
rect 21176 5414 21190 5466
rect 21190 5414 21202 5466
rect 21202 5414 21232 5466
rect 21256 5414 21266 5466
rect 21266 5414 21312 5466
rect 21016 5412 21072 5414
rect 21096 5412 21152 5414
rect 21176 5412 21232 5414
rect 21256 5412 21312 5414
rect 21270 4972 21272 4992
rect 21272 4972 21324 4992
rect 21324 4972 21326 4992
rect 21270 4936 21326 4972
rect 21178 4800 21234 4856
rect 21016 4378 21072 4380
rect 21096 4378 21152 4380
rect 21176 4378 21232 4380
rect 21256 4378 21312 4380
rect 21016 4326 21062 4378
rect 21062 4326 21072 4378
rect 21096 4326 21126 4378
rect 21126 4326 21138 4378
rect 21138 4326 21152 4378
rect 21176 4326 21190 4378
rect 21190 4326 21202 4378
rect 21202 4326 21232 4378
rect 21256 4326 21266 4378
rect 21266 4326 21312 4378
rect 21016 4324 21072 4326
rect 21096 4324 21152 4326
rect 21176 4324 21232 4326
rect 21256 4324 21312 4326
rect 20994 3732 21050 3768
rect 20994 3712 20996 3732
rect 20996 3712 21048 3732
rect 21048 3712 21050 3732
rect 21016 3290 21072 3292
rect 21096 3290 21152 3292
rect 21176 3290 21232 3292
rect 21256 3290 21312 3292
rect 21016 3238 21062 3290
rect 21062 3238 21072 3290
rect 21096 3238 21126 3290
rect 21126 3238 21138 3290
rect 21138 3238 21152 3290
rect 21176 3238 21190 3290
rect 21190 3238 21202 3290
rect 21202 3238 21232 3290
rect 21256 3238 21266 3290
rect 21266 3238 21312 3290
rect 21016 3236 21072 3238
rect 21096 3236 21152 3238
rect 21176 3236 21232 3238
rect 21256 3236 21312 3238
rect 21086 2352 21142 2408
rect 22466 10376 22522 10432
rect 22466 9968 22522 10024
rect 22834 9832 22890 9888
rect 22558 9696 22614 9752
rect 22466 7656 22522 7712
rect 22374 4936 22430 4992
rect 22466 4392 22522 4448
rect 22374 4256 22430 4312
rect 21914 2896 21970 2952
rect 23386 10104 23442 10160
rect 23294 8472 23350 8528
rect 23110 8236 23112 8256
rect 23112 8236 23164 8256
rect 23164 8236 23166 8256
rect 23110 8200 23166 8236
rect 23570 7656 23626 7712
rect 23478 6840 23534 6896
rect 23018 5888 23074 5944
rect 23202 5616 23258 5672
rect 23386 5616 23442 5672
rect 23938 7656 23994 7712
rect 23570 4392 23626 4448
rect 21016 2202 21072 2204
rect 21096 2202 21152 2204
rect 21176 2202 21232 2204
rect 21256 2202 21312 2204
rect 21016 2150 21062 2202
rect 21062 2150 21072 2202
rect 21096 2150 21126 2202
rect 21126 2150 21138 2202
rect 21138 2150 21152 2202
rect 21176 2150 21190 2202
rect 21190 2150 21202 2202
rect 21202 2150 21232 2202
rect 21256 2150 21266 2202
rect 21266 2150 21312 2202
rect 21016 2148 21072 2150
rect 21096 2148 21152 2150
rect 21176 2148 21232 2150
rect 21256 2148 21312 2150
rect 24122 8200 24178 8256
rect 24490 9968 24546 10024
rect 24214 7520 24270 7576
rect 24122 7112 24178 7168
rect 24122 6024 24178 6080
rect 24306 6704 24362 6760
rect 24490 8508 24492 8528
rect 24492 8508 24544 8528
rect 24544 8508 24546 8528
rect 24490 8472 24546 8508
rect 25134 9696 25190 9752
rect 25226 8472 25282 8528
rect 25042 6432 25098 6488
rect 23938 4684 23994 4720
rect 23938 4664 23940 4684
rect 23940 4664 23992 4684
rect 23992 4664 23994 4684
rect 23570 2352 23626 2408
rect 24674 3712 24730 3768
rect 24122 3188 24178 3224
rect 24122 3168 24124 3188
rect 24124 3168 24176 3188
rect 24176 3168 24178 3188
rect 25870 9696 25926 9752
rect 25778 8200 25834 8256
rect 25956 8186 26012 8188
rect 26036 8186 26092 8188
rect 26116 8186 26172 8188
rect 26196 8186 26252 8188
rect 25956 8134 26002 8186
rect 26002 8134 26012 8186
rect 26036 8134 26066 8186
rect 26066 8134 26078 8186
rect 26078 8134 26092 8186
rect 26116 8134 26130 8186
rect 26130 8134 26142 8186
rect 26142 8134 26172 8186
rect 26196 8134 26206 8186
rect 26206 8134 26252 8186
rect 25956 8132 26012 8134
rect 26036 8132 26092 8134
rect 26116 8132 26172 8134
rect 26196 8132 26252 8134
rect 25870 7656 25926 7712
rect 25778 6976 25834 7032
rect 25686 6704 25742 6760
rect 25318 3304 25374 3360
rect 25956 7098 26012 7100
rect 26036 7098 26092 7100
rect 26116 7098 26172 7100
rect 26196 7098 26252 7100
rect 25956 7046 26002 7098
rect 26002 7046 26012 7098
rect 26036 7046 26066 7098
rect 26066 7046 26078 7098
rect 26078 7046 26092 7098
rect 26116 7046 26130 7098
rect 26130 7046 26142 7098
rect 26142 7046 26172 7098
rect 26196 7046 26206 7098
rect 26206 7046 26252 7098
rect 25956 7044 26012 7046
rect 26036 7044 26092 7046
rect 26116 7044 26172 7046
rect 26196 7044 26252 7046
rect 26238 6740 26240 6760
rect 26240 6740 26292 6760
rect 26292 6740 26294 6760
rect 26238 6704 26294 6740
rect 26514 8608 26570 8664
rect 26422 7112 26478 7168
rect 26330 6024 26386 6080
rect 26974 10240 27030 10296
rect 27434 10512 27490 10568
rect 26790 8472 26846 8528
rect 27016 8730 27072 8732
rect 27096 8730 27152 8732
rect 27176 8730 27232 8732
rect 27256 8730 27312 8732
rect 27016 8678 27062 8730
rect 27062 8678 27072 8730
rect 27096 8678 27126 8730
rect 27126 8678 27138 8730
rect 27138 8678 27152 8730
rect 27176 8678 27190 8730
rect 27190 8678 27202 8730
rect 27202 8678 27232 8730
rect 27256 8678 27266 8730
rect 27266 8678 27312 8730
rect 27016 8676 27072 8678
rect 27096 8676 27152 8678
rect 27176 8676 27232 8678
rect 27256 8676 27312 8678
rect 27016 7642 27072 7644
rect 27096 7642 27152 7644
rect 27176 7642 27232 7644
rect 27256 7642 27312 7644
rect 27016 7590 27062 7642
rect 27062 7590 27072 7642
rect 27096 7590 27126 7642
rect 27126 7590 27138 7642
rect 27138 7590 27152 7642
rect 27176 7590 27190 7642
rect 27190 7590 27202 7642
rect 27202 7590 27232 7642
rect 27256 7590 27266 7642
rect 27266 7590 27312 7642
rect 27016 7588 27072 7590
rect 27096 7588 27152 7590
rect 27176 7588 27232 7590
rect 27256 7588 27312 7590
rect 26882 6976 26938 7032
rect 27158 6976 27214 7032
rect 27618 9696 27674 9752
rect 27434 6976 27490 7032
rect 27710 9152 27766 9208
rect 27710 8336 27766 8392
rect 27710 8236 27712 8256
rect 27712 8236 27764 8256
rect 27764 8236 27766 8256
rect 27710 8200 27766 8236
rect 27802 8064 27858 8120
rect 27158 6704 27214 6760
rect 27016 6554 27072 6556
rect 27096 6554 27152 6556
rect 27176 6554 27232 6556
rect 27256 6554 27312 6556
rect 27016 6502 27062 6554
rect 27062 6502 27072 6554
rect 27096 6502 27126 6554
rect 27126 6502 27138 6554
rect 27138 6502 27152 6554
rect 27176 6502 27190 6554
rect 27190 6502 27202 6554
rect 27202 6502 27232 6554
rect 27256 6502 27266 6554
rect 27266 6502 27312 6554
rect 27016 6500 27072 6502
rect 27096 6500 27152 6502
rect 27176 6500 27232 6502
rect 27256 6500 27312 6502
rect 26606 6316 26662 6352
rect 26606 6296 26608 6316
rect 26608 6296 26660 6316
rect 26660 6296 26662 6316
rect 25956 6010 26012 6012
rect 26036 6010 26092 6012
rect 26116 6010 26172 6012
rect 26196 6010 26252 6012
rect 25956 5958 26002 6010
rect 26002 5958 26012 6010
rect 26036 5958 26066 6010
rect 26066 5958 26078 6010
rect 26078 5958 26092 6010
rect 26116 5958 26130 6010
rect 26130 5958 26142 6010
rect 26142 5958 26172 6010
rect 26196 5958 26206 6010
rect 26206 5958 26252 6010
rect 25956 5956 26012 5958
rect 26036 5956 26092 5958
rect 26116 5956 26172 5958
rect 26196 5956 26252 5958
rect 25956 4922 26012 4924
rect 26036 4922 26092 4924
rect 26116 4922 26172 4924
rect 26196 4922 26252 4924
rect 25956 4870 26002 4922
rect 26002 4870 26012 4922
rect 26036 4870 26066 4922
rect 26066 4870 26078 4922
rect 26078 4870 26092 4922
rect 26116 4870 26130 4922
rect 26130 4870 26142 4922
rect 26142 4870 26172 4922
rect 26196 4870 26206 4922
rect 26206 4870 26252 4922
rect 25956 4868 26012 4870
rect 26036 4868 26092 4870
rect 26116 4868 26172 4870
rect 26196 4868 26252 4870
rect 26422 4256 26478 4312
rect 25778 3984 25834 4040
rect 26606 5480 26662 5536
rect 26790 6296 26846 6352
rect 26790 4972 26792 4992
rect 26792 4972 26844 4992
rect 26844 4972 26846 4992
rect 26606 4392 26662 4448
rect 25956 3834 26012 3836
rect 26036 3834 26092 3836
rect 26116 3834 26172 3836
rect 26196 3834 26252 3836
rect 25956 3782 26002 3834
rect 26002 3782 26012 3834
rect 26036 3782 26066 3834
rect 26066 3782 26078 3834
rect 26078 3782 26092 3834
rect 26116 3782 26130 3834
rect 26130 3782 26142 3834
rect 26142 3782 26172 3834
rect 26196 3782 26206 3834
rect 26206 3782 26252 3834
rect 25956 3780 26012 3782
rect 26036 3780 26092 3782
rect 26116 3780 26172 3782
rect 26196 3780 26252 3782
rect 26146 3576 26202 3632
rect 26514 3984 26570 4040
rect 26790 4936 26846 4972
rect 26606 3848 26662 3904
rect 26514 3712 26570 3768
rect 26422 3576 26478 3632
rect 26422 3304 26478 3360
rect 25962 2896 26018 2952
rect 26606 2896 26662 2952
rect 25778 2760 25834 2816
rect 25956 2746 26012 2748
rect 26036 2746 26092 2748
rect 26116 2746 26172 2748
rect 26196 2746 26252 2748
rect 25956 2694 26002 2746
rect 26002 2694 26012 2746
rect 26036 2694 26066 2746
rect 26066 2694 26078 2746
rect 26078 2694 26092 2746
rect 26116 2694 26130 2746
rect 26130 2694 26142 2746
rect 26142 2694 26172 2746
rect 26196 2694 26206 2746
rect 26206 2694 26252 2746
rect 25956 2692 26012 2694
rect 26036 2692 26092 2694
rect 26116 2692 26172 2694
rect 26196 2692 26252 2694
rect 27618 6316 27674 6352
rect 27618 6296 27620 6316
rect 27620 6296 27672 6316
rect 27672 6296 27674 6316
rect 27342 5752 27398 5808
rect 27016 5466 27072 5468
rect 27096 5466 27152 5468
rect 27176 5466 27232 5468
rect 27256 5466 27312 5468
rect 27016 5414 27062 5466
rect 27062 5414 27072 5466
rect 27096 5414 27126 5466
rect 27126 5414 27138 5466
rect 27138 5414 27152 5466
rect 27176 5414 27190 5466
rect 27190 5414 27202 5466
rect 27202 5414 27232 5466
rect 27256 5414 27266 5466
rect 27266 5414 27312 5466
rect 27016 5412 27072 5414
rect 27096 5412 27152 5414
rect 27176 5412 27232 5414
rect 27256 5412 27312 5414
rect 27016 4378 27072 4380
rect 27096 4378 27152 4380
rect 27176 4378 27232 4380
rect 27256 4378 27312 4380
rect 27016 4326 27062 4378
rect 27062 4326 27072 4378
rect 27096 4326 27126 4378
rect 27126 4326 27138 4378
rect 27138 4326 27152 4378
rect 27176 4326 27190 4378
rect 27190 4326 27202 4378
rect 27202 4326 27232 4378
rect 27256 4326 27266 4378
rect 27266 4326 27312 4378
rect 27016 4324 27072 4326
rect 27096 4324 27152 4326
rect 27176 4324 27232 4326
rect 27256 4324 27312 4326
rect 27016 3290 27072 3292
rect 27096 3290 27152 3292
rect 27176 3290 27232 3292
rect 27256 3290 27312 3292
rect 27016 3238 27062 3290
rect 27062 3238 27072 3290
rect 27096 3238 27126 3290
rect 27126 3238 27138 3290
rect 27138 3238 27152 3290
rect 27176 3238 27190 3290
rect 27190 3238 27202 3290
rect 27202 3238 27232 3290
rect 27256 3238 27266 3290
rect 27266 3238 27312 3290
rect 27016 3236 27072 3238
rect 27096 3236 27152 3238
rect 27176 3236 27232 3238
rect 27256 3236 27312 3238
rect 27250 2796 27252 2816
rect 27252 2796 27304 2816
rect 27304 2796 27306 2816
rect 27250 2760 27306 2796
rect 27016 2202 27072 2204
rect 27096 2202 27152 2204
rect 27176 2202 27232 2204
rect 27256 2202 27312 2204
rect 27016 2150 27062 2202
rect 27062 2150 27072 2202
rect 27096 2150 27126 2202
rect 27126 2150 27138 2202
rect 27138 2150 27152 2202
rect 27176 2150 27190 2202
rect 27190 2150 27202 2202
rect 27202 2150 27232 2202
rect 27256 2150 27266 2202
rect 27266 2150 27312 2202
rect 27016 2148 27072 2150
rect 27096 2148 27152 2150
rect 27176 2148 27232 2150
rect 27256 2148 27312 2150
rect 26514 1944 26570 2000
rect 27434 3168 27490 3224
rect 27618 2896 27674 2952
rect 27526 2760 27582 2816
rect 27342 1536 27398 1592
rect 28446 10104 28502 10160
rect 28354 9968 28410 10024
rect 28170 9832 28226 9888
rect 28078 8608 28134 8664
rect 28262 8628 28318 8664
rect 28262 8608 28264 8628
rect 28264 8608 28316 8628
rect 28316 8608 28318 8628
rect 28170 8200 28226 8256
rect 28538 7656 28594 7712
rect 28538 7112 28594 7168
rect 28722 8064 28778 8120
rect 28722 7964 28724 7984
rect 28724 7964 28776 7984
rect 28776 7964 28778 7984
rect 28722 7928 28778 7964
rect 28906 8628 28962 8664
rect 28906 8608 28908 8628
rect 28908 8608 28960 8628
rect 28960 8608 28962 8628
rect 29090 8608 29146 8664
rect 29458 10240 29514 10296
rect 28906 8200 28962 8256
rect 29182 6976 29238 7032
rect 27986 6432 28042 6488
rect 27894 4936 27950 4992
rect 28814 6296 28870 6352
rect 27986 4156 27988 4176
rect 27988 4156 28040 4176
rect 28040 4156 28042 4176
rect 27986 4120 28042 4156
rect 28722 6024 28778 6080
rect 28170 3712 28226 3768
rect 29366 7112 29422 7168
rect 29826 8608 29882 8664
rect 29734 7520 29790 7576
rect 29642 6704 29698 6760
rect 30286 7928 30342 7984
rect 30286 7656 30342 7712
rect 28906 3848 28962 3904
rect 28630 2352 28686 2408
rect 27710 720 27766 776
rect 29734 3032 29790 3088
rect 30010 6024 30066 6080
rect 30562 9968 30618 10024
rect 30470 8064 30526 8120
rect 29918 3440 29974 3496
rect 30194 3576 30250 3632
rect 30654 6160 30710 6216
rect 31114 9832 31170 9888
rect 31666 9696 31722 9752
rect 30930 8608 30986 8664
rect 30838 5752 30894 5808
rect 30562 4800 30618 4856
rect 31114 6704 31170 6760
rect 31022 6024 31078 6080
rect 32034 9152 32090 9208
rect 32034 8472 32090 8528
rect 31956 8186 32012 8188
rect 32036 8186 32092 8188
rect 32116 8186 32172 8188
rect 32196 8186 32252 8188
rect 31956 8134 32002 8186
rect 32002 8134 32012 8186
rect 32036 8134 32066 8186
rect 32066 8134 32078 8186
rect 32078 8134 32092 8186
rect 32116 8134 32130 8186
rect 32130 8134 32142 8186
rect 32142 8134 32172 8186
rect 32196 8134 32206 8186
rect 32206 8134 32252 8186
rect 31956 8132 32012 8134
rect 32036 8132 32092 8134
rect 32116 8132 32172 8134
rect 32196 8132 32252 8134
rect 32402 8472 32458 8528
rect 32402 8200 32458 8256
rect 33506 9832 33562 9888
rect 33414 9560 33470 9616
rect 33016 8730 33072 8732
rect 33096 8730 33152 8732
rect 33176 8730 33232 8732
rect 33256 8730 33312 8732
rect 33016 8678 33062 8730
rect 33062 8678 33072 8730
rect 33096 8678 33126 8730
rect 33126 8678 33138 8730
rect 33138 8678 33152 8730
rect 33176 8678 33190 8730
rect 33190 8678 33202 8730
rect 33202 8678 33232 8730
rect 33256 8678 33266 8730
rect 33266 8678 33312 8730
rect 33016 8676 33072 8678
rect 33096 8676 33152 8678
rect 33176 8676 33232 8678
rect 33256 8676 33312 8678
rect 32862 8628 32918 8664
rect 32862 8608 32864 8628
rect 32864 8608 32916 8628
rect 32916 8608 32918 8628
rect 32954 8472 33010 8528
rect 32218 7656 32274 7712
rect 31758 7112 31814 7168
rect 31956 7098 32012 7100
rect 32036 7098 32092 7100
rect 32116 7098 32172 7100
rect 32196 7098 32252 7100
rect 31956 7046 32002 7098
rect 32002 7046 32012 7098
rect 32036 7046 32066 7098
rect 32066 7046 32078 7098
rect 32078 7046 32092 7098
rect 32116 7046 32130 7098
rect 32130 7046 32142 7098
rect 32142 7046 32172 7098
rect 32196 7046 32206 7098
rect 32206 7046 32252 7098
rect 31956 7044 32012 7046
rect 32036 7044 32092 7046
rect 32116 7044 32172 7046
rect 32196 7044 32252 7046
rect 31758 6976 31814 7032
rect 31666 6724 31722 6760
rect 31666 6704 31668 6724
rect 31668 6704 31720 6724
rect 31720 6704 31722 6724
rect 31758 6160 31814 6216
rect 31114 5344 31170 5400
rect 31574 5072 31630 5128
rect 32034 6740 32036 6760
rect 32036 6740 32088 6760
rect 32088 6740 32090 6760
rect 32034 6704 32090 6740
rect 32310 6604 32312 6624
rect 32312 6604 32364 6624
rect 32364 6604 32366 6624
rect 32310 6568 32366 6604
rect 31956 6010 32012 6012
rect 32036 6010 32092 6012
rect 32116 6010 32172 6012
rect 32196 6010 32252 6012
rect 31956 5958 32002 6010
rect 32002 5958 32012 6010
rect 32036 5958 32066 6010
rect 32066 5958 32078 6010
rect 32078 5958 32092 6010
rect 32116 5958 32130 6010
rect 32130 5958 32142 6010
rect 32142 5958 32172 6010
rect 32196 5958 32206 6010
rect 32206 5958 32252 6010
rect 31956 5956 32012 5958
rect 32036 5956 32092 5958
rect 32116 5956 32172 5958
rect 32196 5956 32252 5958
rect 32218 5652 32220 5672
rect 32220 5652 32272 5672
rect 32272 5652 32274 5672
rect 32218 5616 32274 5652
rect 31956 4922 32012 4924
rect 32036 4922 32092 4924
rect 32116 4922 32172 4924
rect 32196 4922 32252 4924
rect 31956 4870 32002 4922
rect 32002 4870 32012 4922
rect 32036 4870 32066 4922
rect 32066 4870 32078 4922
rect 32078 4870 32092 4922
rect 32116 4870 32130 4922
rect 32130 4870 32142 4922
rect 32142 4870 32172 4922
rect 32196 4870 32206 4922
rect 32206 4870 32252 4922
rect 31956 4868 32012 4870
rect 32036 4868 32092 4870
rect 32116 4868 32172 4870
rect 32196 4868 32252 4870
rect 31850 4664 31906 4720
rect 32034 4664 32090 4720
rect 31956 3834 32012 3836
rect 32036 3834 32092 3836
rect 32116 3834 32172 3836
rect 32196 3834 32252 3836
rect 31956 3782 32002 3834
rect 32002 3782 32012 3834
rect 32036 3782 32066 3834
rect 32066 3782 32078 3834
rect 32078 3782 32092 3834
rect 32116 3782 32130 3834
rect 32130 3782 32142 3834
rect 32142 3782 32172 3834
rect 32196 3782 32206 3834
rect 32206 3782 32252 3834
rect 31956 3780 32012 3782
rect 32036 3780 32092 3782
rect 32116 3780 32172 3782
rect 32196 3780 32252 3782
rect 32126 3032 32182 3088
rect 31956 2746 32012 2748
rect 32036 2746 32092 2748
rect 32116 2746 32172 2748
rect 32196 2746 32252 2748
rect 29826 720 29882 776
rect 31956 2694 32002 2746
rect 32002 2694 32012 2746
rect 32036 2694 32066 2746
rect 32066 2694 32078 2746
rect 32078 2694 32092 2746
rect 32116 2694 32130 2746
rect 32130 2694 32142 2746
rect 32142 2694 32172 2746
rect 32196 2694 32206 2746
rect 32206 2694 32252 2746
rect 31956 2692 32012 2694
rect 32036 2692 32092 2694
rect 32116 2692 32172 2694
rect 32196 2692 32252 2694
rect 32770 8064 32826 8120
rect 32862 7928 32918 7984
rect 33230 8200 33286 8256
rect 33782 9832 33838 9888
rect 33690 9696 33746 9752
rect 33598 7792 33654 7848
rect 34058 9968 34114 10024
rect 33016 7642 33072 7644
rect 33096 7642 33152 7644
rect 33176 7642 33232 7644
rect 33256 7642 33312 7644
rect 33016 7590 33062 7642
rect 33062 7590 33072 7642
rect 33096 7590 33126 7642
rect 33126 7590 33138 7642
rect 33138 7590 33152 7642
rect 33176 7590 33190 7642
rect 33190 7590 33202 7642
rect 33202 7590 33232 7642
rect 33256 7590 33266 7642
rect 33266 7590 33312 7642
rect 33016 7588 33072 7590
rect 33096 7588 33152 7590
rect 33176 7588 33232 7590
rect 33256 7588 33312 7590
rect 32954 7384 33010 7440
rect 33230 7268 33286 7304
rect 33230 7248 33232 7268
rect 33232 7248 33284 7268
rect 33284 7248 33286 7268
rect 32954 6840 33010 6896
rect 33016 6554 33072 6556
rect 33096 6554 33152 6556
rect 33176 6554 33232 6556
rect 33256 6554 33312 6556
rect 33016 6502 33062 6554
rect 33062 6502 33072 6554
rect 33096 6502 33126 6554
rect 33126 6502 33138 6554
rect 33138 6502 33152 6554
rect 33176 6502 33190 6554
rect 33190 6502 33202 6554
rect 33202 6502 33232 6554
rect 33256 6502 33266 6554
rect 33266 6502 33312 6554
rect 33016 6500 33072 6502
rect 33096 6500 33152 6502
rect 33176 6500 33232 6502
rect 33256 6500 33312 6502
rect 33230 5888 33286 5944
rect 32862 5616 32918 5672
rect 32770 5344 32826 5400
rect 33016 5466 33072 5468
rect 33096 5466 33152 5468
rect 33176 5466 33232 5468
rect 33256 5466 33312 5468
rect 33016 5414 33062 5466
rect 33062 5414 33072 5466
rect 33096 5414 33126 5466
rect 33126 5414 33138 5466
rect 33138 5414 33152 5466
rect 33176 5414 33190 5466
rect 33190 5414 33202 5466
rect 33202 5414 33232 5466
rect 33256 5414 33266 5466
rect 33266 5414 33312 5466
rect 33016 5412 33072 5414
rect 33096 5412 33152 5414
rect 33176 5412 33232 5414
rect 33256 5412 33312 5414
rect 32862 4664 32918 4720
rect 33016 4378 33072 4380
rect 33096 4378 33152 4380
rect 33176 4378 33232 4380
rect 33256 4378 33312 4380
rect 33016 4326 33062 4378
rect 33062 4326 33072 4378
rect 33096 4326 33126 4378
rect 33126 4326 33138 4378
rect 33138 4326 33152 4378
rect 33176 4326 33190 4378
rect 33190 4326 33202 4378
rect 33202 4326 33232 4378
rect 33256 4326 33266 4378
rect 33266 4326 33312 4378
rect 33016 4324 33072 4326
rect 33096 4324 33152 4326
rect 33176 4324 33232 4326
rect 33256 4324 33312 4326
rect 32954 4120 33010 4176
rect 32770 3168 32826 3224
rect 33016 3290 33072 3292
rect 33096 3290 33152 3292
rect 33176 3290 33232 3292
rect 33256 3290 33312 3292
rect 33016 3238 33062 3290
rect 33062 3238 33072 3290
rect 33096 3238 33126 3290
rect 33126 3238 33138 3290
rect 33138 3238 33152 3290
rect 33176 3238 33190 3290
rect 33190 3238 33202 3290
rect 33202 3238 33232 3290
rect 33256 3238 33266 3290
rect 33266 3238 33312 3290
rect 33016 3236 33072 3238
rect 33096 3236 33152 3238
rect 33176 3236 33232 3238
rect 33256 3236 33312 3238
rect 32586 2760 32642 2816
rect 33414 3052 33470 3088
rect 33414 3032 33416 3052
rect 33416 3032 33468 3052
rect 33468 3032 33470 3052
rect 32954 2760 33010 2816
rect 33016 2202 33072 2204
rect 33096 2202 33152 2204
rect 33176 2202 33232 2204
rect 33256 2202 33312 2204
rect 33016 2150 33062 2202
rect 33062 2150 33072 2202
rect 33096 2150 33126 2202
rect 33126 2150 33138 2202
rect 33138 2150 33152 2202
rect 33176 2150 33190 2202
rect 33190 2150 33202 2202
rect 33202 2150 33232 2202
rect 33256 2150 33266 2202
rect 33266 2150 33312 2202
rect 33016 2148 33072 2150
rect 33096 2148 33152 2150
rect 33176 2148 33232 2150
rect 33256 2148 33312 2150
rect 33506 992 33562 1048
rect 34610 9288 34666 9344
rect 35438 9152 35494 9208
rect 35254 5208 35310 5264
rect 35438 4564 35440 4584
rect 35440 4564 35492 4584
rect 35492 4564 35494 4584
rect 35438 4528 35494 4564
rect 35806 856 35862 912
rect 35714 720 35770 776
rect 36634 2896 36690 2952
rect 37278 5772 37334 5808
rect 37278 5752 37280 5772
rect 37280 5752 37332 5772
rect 37332 5752 37334 5772
rect 37278 5636 37334 5672
rect 37278 5616 37280 5636
rect 37280 5616 37332 5636
rect 37332 5616 37334 5636
rect 37278 3984 37334 4040
rect 37094 1944 37150 2000
rect 39762 9832 39818 9888
rect 39670 9560 39726 9616
rect 38934 9288 38990 9344
rect 37956 8186 38012 8188
rect 38036 8186 38092 8188
rect 38116 8186 38172 8188
rect 38196 8186 38252 8188
rect 37956 8134 38002 8186
rect 38002 8134 38012 8186
rect 38036 8134 38066 8186
rect 38066 8134 38078 8186
rect 38078 8134 38092 8186
rect 38116 8134 38130 8186
rect 38130 8134 38142 8186
rect 38142 8134 38172 8186
rect 38196 8134 38206 8186
rect 38206 8134 38252 8186
rect 37956 8132 38012 8134
rect 38036 8132 38092 8134
rect 38116 8132 38172 8134
rect 38196 8132 38252 8134
rect 37956 7098 38012 7100
rect 38036 7098 38092 7100
rect 38116 7098 38172 7100
rect 38196 7098 38252 7100
rect 37956 7046 38002 7098
rect 38002 7046 38012 7098
rect 38036 7046 38066 7098
rect 38066 7046 38078 7098
rect 38078 7046 38092 7098
rect 38116 7046 38130 7098
rect 38130 7046 38142 7098
rect 38142 7046 38172 7098
rect 38196 7046 38206 7098
rect 38206 7046 38252 7098
rect 37956 7044 38012 7046
rect 38036 7044 38092 7046
rect 38116 7044 38172 7046
rect 38196 7044 38252 7046
rect 38014 6296 38070 6352
rect 37956 6010 38012 6012
rect 38036 6010 38092 6012
rect 38116 6010 38172 6012
rect 38196 6010 38252 6012
rect 37956 5958 38002 6010
rect 38002 5958 38012 6010
rect 38036 5958 38066 6010
rect 38066 5958 38078 6010
rect 38078 5958 38092 6010
rect 38116 5958 38130 6010
rect 38130 5958 38142 6010
rect 38142 5958 38172 6010
rect 38196 5958 38206 6010
rect 38206 5958 38252 6010
rect 37956 5956 38012 5958
rect 38036 5956 38092 5958
rect 38116 5956 38172 5958
rect 38196 5956 38252 5958
rect 37956 4922 38012 4924
rect 38036 4922 38092 4924
rect 38116 4922 38172 4924
rect 38196 4922 38252 4924
rect 37956 4870 38002 4922
rect 38002 4870 38012 4922
rect 38036 4870 38066 4922
rect 38066 4870 38078 4922
rect 38078 4870 38092 4922
rect 38116 4870 38130 4922
rect 38130 4870 38142 4922
rect 38142 4870 38172 4922
rect 38196 4870 38206 4922
rect 38206 4870 38252 4922
rect 37956 4868 38012 4870
rect 38036 4868 38092 4870
rect 38116 4868 38172 4870
rect 38196 4868 38252 4870
rect 37956 3834 38012 3836
rect 38036 3834 38092 3836
rect 38116 3834 38172 3836
rect 38196 3834 38252 3836
rect 37956 3782 38002 3834
rect 38002 3782 38012 3834
rect 38036 3782 38066 3834
rect 38066 3782 38078 3834
rect 38078 3782 38092 3834
rect 38116 3782 38130 3834
rect 38130 3782 38142 3834
rect 38142 3782 38172 3834
rect 38196 3782 38206 3834
rect 38206 3782 38252 3834
rect 37956 3780 38012 3782
rect 38036 3780 38092 3782
rect 38116 3780 38172 3782
rect 38196 3780 38252 3782
rect 37956 2746 38012 2748
rect 38036 2746 38092 2748
rect 38116 2746 38172 2748
rect 38196 2746 38252 2748
rect 37956 2694 38002 2746
rect 38002 2694 38012 2746
rect 38036 2694 38066 2746
rect 38066 2694 38078 2746
rect 38078 2694 38092 2746
rect 38116 2694 38130 2746
rect 38130 2694 38142 2746
rect 38142 2694 38172 2746
rect 38196 2694 38206 2746
rect 38206 2694 38252 2746
rect 37956 2692 38012 2694
rect 38036 2692 38092 2694
rect 38116 2692 38172 2694
rect 38196 2692 38252 2694
rect 38658 8472 38714 8528
rect 38566 6840 38622 6896
rect 38658 6296 38714 6352
rect 37922 1672 37978 1728
rect 38290 1400 38346 1456
rect 38842 8336 38898 8392
rect 39486 9016 39542 9072
rect 39394 8880 39450 8936
rect 39016 8730 39072 8732
rect 39096 8730 39152 8732
rect 39176 8730 39232 8732
rect 39256 8730 39312 8732
rect 39016 8678 39062 8730
rect 39062 8678 39072 8730
rect 39096 8678 39126 8730
rect 39126 8678 39138 8730
rect 39138 8678 39152 8730
rect 39176 8678 39190 8730
rect 39190 8678 39202 8730
rect 39202 8678 39232 8730
rect 39256 8678 39266 8730
rect 39266 8678 39312 8730
rect 39016 8676 39072 8678
rect 39096 8676 39152 8678
rect 39176 8676 39232 8678
rect 39256 8676 39312 8678
rect 39026 8200 39082 8256
rect 39394 7928 39450 7984
rect 39394 7692 39396 7712
rect 39396 7692 39448 7712
rect 39448 7692 39450 7712
rect 39394 7656 39450 7692
rect 39016 7642 39072 7644
rect 39096 7642 39152 7644
rect 39176 7642 39232 7644
rect 39256 7642 39312 7644
rect 39016 7590 39062 7642
rect 39062 7590 39072 7642
rect 39096 7590 39126 7642
rect 39126 7590 39138 7642
rect 39138 7590 39152 7642
rect 39176 7590 39190 7642
rect 39190 7590 39202 7642
rect 39202 7590 39232 7642
rect 39256 7590 39266 7642
rect 39266 7590 39312 7642
rect 39016 7588 39072 7590
rect 39096 7588 39152 7590
rect 39176 7588 39232 7590
rect 39256 7588 39312 7590
rect 38934 7384 38990 7440
rect 39394 7148 39396 7168
rect 39396 7148 39448 7168
rect 39448 7148 39450 7168
rect 39394 7112 39450 7148
rect 39578 8744 39634 8800
rect 39394 6568 39450 6624
rect 39016 6554 39072 6556
rect 39096 6554 39152 6556
rect 39176 6554 39232 6556
rect 39256 6554 39312 6556
rect 39016 6502 39062 6554
rect 39062 6502 39072 6554
rect 39096 6502 39126 6554
rect 39126 6502 39138 6554
rect 39138 6502 39152 6554
rect 39176 6502 39190 6554
rect 39190 6502 39202 6554
rect 39202 6502 39232 6554
rect 39256 6502 39266 6554
rect 39266 6502 39312 6554
rect 39016 6500 39072 6502
rect 39096 6500 39152 6502
rect 39176 6500 39232 6502
rect 39256 6500 39312 6502
rect 38842 6060 38844 6080
rect 38844 6060 38896 6080
rect 38896 6060 38898 6080
rect 38842 6024 38898 6060
rect 39394 5788 39396 5808
rect 39396 5788 39448 5808
rect 39448 5788 39450 5808
rect 39394 5752 39450 5788
rect 39210 5652 39212 5672
rect 39212 5652 39264 5672
rect 39264 5652 39266 5672
rect 39210 5616 39266 5652
rect 39016 5466 39072 5468
rect 39096 5466 39152 5468
rect 39176 5466 39232 5468
rect 39256 5466 39312 5468
rect 39016 5414 39062 5466
rect 39062 5414 39072 5466
rect 39096 5414 39126 5466
rect 39126 5414 39138 5466
rect 39138 5414 39152 5466
rect 39176 5414 39190 5466
rect 39190 5414 39202 5466
rect 39202 5414 39232 5466
rect 39256 5414 39266 5466
rect 39266 5414 39312 5466
rect 39016 5412 39072 5414
rect 39096 5412 39152 5414
rect 39176 5412 39232 5414
rect 39256 5412 39312 5414
rect 39394 5208 39450 5264
rect 39026 4972 39028 4992
rect 39028 4972 39080 4992
rect 39080 4972 39082 4992
rect 39026 4936 39082 4972
rect 39394 4700 39396 4720
rect 39396 4700 39448 4720
rect 39448 4700 39450 4720
rect 39394 4664 39450 4700
rect 39016 4378 39072 4380
rect 39096 4378 39152 4380
rect 39176 4378 39232 4380
rect 39256 4378 39312 4380
rect 39016 4326 39062 4378
rect 39062 4326 39072 4378
rect 39096 4326 39126 4378
rect 39126 4326 39138 4378
rect 39138 4326 39152 4378
rect 39176 4326 39190 4378
rect 39190 4326 39202 4378
rect 39202 4326 39232 4378
rect 39256 4326 39266 4378
rect 39266 4326 39312 4378
rect 39016 4324 39072 4326
rect 39096 4324 39152 4326
rect 39176 4324 39232 4326
rect 39256 4324 39312 4326
rect 39394 4120 39450 4176
rect 39026 3884 39028 3904
rect 39028 3884 39080 3904
rect 39080 3884 39082 3904
rect 39026 3848 39082 3884
rect 39394 3612 39396 3632
rect 39396 3612 39448 3632
rect 39448 3612 39450 3632
rect 39394 3576 39450 3612
rect 39016 3290 39072 3292
rect 39096 3290 39152 3292
rect 39176 3290 39232 3292
rect 39256 3290 39312 3292
rect 39016 3238 39062 3290
rect 39062 3238 39072 3290
rect 39096 3238 39126 3290
rect 39126 3238 39138 3290
rect 39138 3238 39152 3290
rect 39176 3238 39190 3290
rect 39190 3238 39202 3290
rect 39202 3238 39232 3290
rect 39256 3238 39266 3290
rect 39266 3238 39312 3290
rect 39016 3236 39072 3238
rect 39096 3236 39152 3238
rect 39176 3236 39232 3238
rect 39256 3236 39312 3238
rect 39394 3032 39450 3088
rect 39026 2796 39028 2816
rect 39028 2796 39080 2816
rect 39080 2796 39082 2816
rect 39026 2760 39082 2796
rect 39394 2524 39396 2544
rect 39396 2524 39448 2544
rect 39448 2524 39450 2544
rect 39394 2488 39450 2524
rect 38750 1808 38806 1864
rect 39016 2202 39072 2204
rect 39096 2202 39152 2204
rect 39176 2202 39232 2204
rect 39256 2202 39312 2204
rect 39016 2150 39062 2202
rect 39062 2150 39072 2202
rect 39096 2150 39126 2202
rect 39126 2150 39138 2202
rect 39138 2150 39152 2202
rect 39176 2150 39190 2202
rect 39190 2150 39202 2202
rect 39202 2150 39232 2202
rect 39256 2150 39266 2202
rect 39266 2150 39312 2202
rect 39016 2148 39072 2150
rect 39096 2148 39152 2150
rect 39176 2148 39232 2150
rect 39256 2148 39312 2150
rect 38934 1944 38990 2000
rect 39946 5516 39948 5536
rect 39948 5516 40000 5536
rect 40000 5516 40002 5536
rect 39946 5480 40002 5516
rect 39854 4392 39910 4448
rect 39670 1128 39726 1184
rect 39946 3340 39948 3360
rect 39948 3340 40000 3360
rect 40000 3340 40002 3360
rect 39946 3304 40002 3340
rect 39946 2252 39948 2272
rect 39948 2252 40000 2272
rect 40000 2252 40002 2272
rect 39946 2216 40002 2252
rect 39854 1264 39910 1320
<< metal3 >>
rect 4705 10706 4771 10709
rect 10041 10706 10107 10709
rect 4705 10704 10107 10706
rect 4705 10648 4710 10704
rect 4766 10648 10046 10704
rect 10102 10648 10107 10704
rect 4705 10646 10107 10648
rect 4705 10643 4771 10646
rect 10041 10643 10107 10646
rect 4981 10570 5047 10573
rect 10685 10570 10751 10573
rect 4981 10568 10751 10570
rect 4981 10512 4986 10568
rect 5042 10512 10690 10568
rect 10746 10512 10751 10568
rect 4981 10510 10751 10512
rect 4981 10507 5047 10510
rect 10685 10507 10751 10510
rect 10869 10570 10935 10573
rect 17677 10570 17743 10573
rect 27429 10570 27495 10573
rect 10869 10568 17743 10570
rect 10869 10512 10874 10568
rect 10930 10512 17682 10568
rect 17738 10512 17743 10568
rect 10869 10510 17743 10512
rect 10869 10507 10935 10510
rect 17677 10507 17743 10510
rect 22050 10568 27495 10570
rect 22050 10512 27434 10568
rect 27490 10512 27495 10568
rect 22050 10510 27495 10512
rect 5257 10434 5323 10437
rect 9305 10434 9371 10437
rect 22050 10434 22110 10510
rect 27429 10507 27495 10510
rect 5257 10432 9371 10434
rect 5257 10376 5262 10432
rect 5318 10376 9310 10432
rect 9366 10376 9371 10432
rect 5257 10374 9371 10376
rect 5257 10371 5323 10374
rect 9305 10371 9371 10374
rect 17174 10374 22110 10434
rect 22461 10434 22527 10437
rect 26734 10434 26740 10436
rect 22461 10432 26740 10434
rect 22461 10376 22466 10432
rect 22522 10376 26740 10432
rect 22461 10374 26740 10376
rect 4521 10298 4587 10301
rect 8201 10298 8267 10301
rect 4521 10296 8267 10298
rect 4521 10240 4526 10296
rect 4582 10240 8206 10296
rect 8262 10240 8267 10296
rect 4521 10238 8267 10240
rect 4521 10235 4587 10238
rect 8201 10235 8267 10238
rect 9397 10298 9463 10301
rect 11237 10298 11303 10301
rect 9397 10296 11303 10298
rect 9397 10240 9402 10296
rect 9458 10240 11242 10296
rect 11298 10240 11303 10296
rect 9397 10238 11303 10240
rect 9397 10235 9463 10238
rect 11237 10235 11303 10238
rect 13445 10298 13511 10301
rect 16113 10298 16179 10301
rect 13445 10296 16179 10298
rect 13445 10240 13450 10296
rect 13506 10240 16118 10296
rect 16174 10240 16179 10296
rect 13445 10238 16179 10240
rect 13445 10235 13511 10238
rect 16113 10235 16179 10238
rect 2630 10100 2636 10164
rect 2700 10162 2706 10164
rect 17174 10162 17234 10374
rect 22461 10371 22527 10374
rect 26734 10372 26740 10374
rect 26804 10372 26810 10436
rect 17401 10298 17467 10301
rect 24894 10298 24900 10300
rect 17401 10296 24900 10298
rect 17401 10240 17406 10296
rect 17462 10240 24900 10296
rect 17401 10238 24900 10240
rect 17401 10235 17467 10238
rect 24894 10236 24900 10238
rect 24964 10236 24970 10300
rect 26969 10298 27035 10301
rect 29453 10298 29519 10301
rect 26969 10296 29519 10298
rect 26969 10240 26974 10296
rect 27030 10240 29458 10296
rect 29514 10240 29519 10296
rect 26969 10238 29519 10240
rect 26969 10235 27035 10238
rect 29453 10235 29519 10238
rect 2700 10102 17234 10162
rect 23381 10162 23447 10165
rect 28441 10162 28507 10165
rect 23381 10160 28507 10162
rect 23381 10104 23386 10160
rect 23442 10104 28446 10160
rect 28502 10104 28507 10160
rect 23381 10102 28507 10104
rect 2700 10100 2706 10102
rect 23381 10099 23447 10102
rect 28441 10099 28507 10102
rect 7782 9964 7788 10028
rect 7852 10026 7858 10028
rect 22461 10026 22527 10029
rect 23422 10026 23428 10028
rect 7852 10024 22527 10026
rect 7852 9968 22466 10024
rect 22522 9968 22527 10024
rect 7852 9966 22527 9968
rect 7852 9964 7858 9966
rect 22461 9963 22527 9966
rect 22694 9966 23428 10026
rect 0 9890 120 9920
rect 2313 9890 2379 9893
rect 0 9888 2379 9890
rect 0 9832 2318 9888
rect 2374 9832 2379 9888
rect 0 9830 2379 9832
rect 0 9800 120 9830
rect 2313 9827 2379 9830
rect 7557 9890 7623 9893
rect 9857 9890 9923 9893
rect 7557 9888 9923 9890
rect 7557 9832 7562 9888
rect 7618 9832 9862 9888
rect 9918 9832 9923 9888
rect 7557 9830 9923 9832
rect 7557 9827 7623 9830
rect 9857 9827 9923 9830
rect 10041 9890 10107 9893
rect 17401 9890 17467 9893
rect 10041 9888 17467 9890
rect 10041 9832 10046 9888
rect 10102 9832 17406 9888
rect 17462 9832 17467 9888
rect 10041 9830 17467 9832
rect 10041 9827 10107 9830
rect 17401 9827 17467 9830
rect 17677 9890 17743 9893
rect 22694 9890 22754 9966
rect 23422 9964 23428 9966
rect 23492 9964 23498 10028
rect 24485 10026 24551 10029
rect 28349 10026 28415 10029
rect 24485 10024 28415 10026
rect 24485 9968 24490 10024
rect 24546 9968 28354 10024
rect 28410 9968 28415 10024
rect 24485 9966 28415 9968
rect 24485 9963 24551 9966
rect 28349 9963 28415 9966
rect 30557 10026 30623 10029
rect 34053 10026 34119 10029
rect 30557 10024 34119 10026
rect 30557 9968 30562 10024
rect 30618 9968 34058 10024
rect 34114 9968 34119 10024
rect 30557 9966 34119 9968
rect 30557 9963 30623 9966
rect 34053 9963 34119 9966
rect 17677 9888 22754 9890
rect 17677 9832 17682 9888
rect 17738 9832 22754 9888
rect 17677 9830 22754 9832
rect 22829 9890 22895 9893
rect 28165 9890 28231 9893
rect 22829 9888 28231 9890
rect 22829 9832 22834 9888
rect 22890 9832 28170 9888
rect 28226 9832 28231 9888
rect 22829 9830 28231 9832
rect 17677 9827 17743 9830
rect 22829 9827 22895 9830
rect 28165 9827 28231 9830
rect 31109 9890 31175 9893
rect 33501 9890 33567 9893
rect 33777 9892 33843 9893
rect 31109 9888 33567 9890
rect 31109 9832 31114 9888
rect 31170 9832 33506 9888
rect 33562 9832 33567 9888
rect 31109 9830 33567 9832
rect 31109 9827 31175 9830
rect 33501 9827 33567 9830
rect 33726 9828 33732 9892
rect 33796 9890 33843 9892
rect 39757 9890 39823 9893
rect 40880 9890 41000 9920
rect 33796 9888 33888 9890
rect 33838 9832 33888 9888
rect 33796 9830 33888 9832
rect 39757 9888 41000 9890
rect 39757 9832 39762 9888
rect 39818 9832 41000 9888
rect 39757 9830 41000 9832
rect 33796 9828 33843 9830
rect 33777 9827 33843 9828
rect 39757 9827 39823 9830
rect 40880 9800 41000 9830
rect 7925 9754 7991 9757
rect 13169 9754 13235 9757
rect 7925 9752 13235 9754
rect 7925 9696 7930 9752
rect 7986 9696 13174 9752
rect 13230 9696 13235 9752
rect 7925 9694 13235 9696
rect 7925 9691 7991 9694
rect 13169 9691 13235 9694
rect 14825 9754 14891 9757
rect 19517 9754 19583 9757
rect 14825 9752 19583 9754
rect 14825 9696 14830 9752
rect 14886 9696 19522 9752
rect 19578 9696 19583 9752
rect 14825 9694 19583 9696
rect 14825 9691 14891 9694
rect 19517 9691 19583 9694
rect 22553 9754 22619 9757
rect 25129 9754 25195 9757
rect 22553 9752 25195 9754
rect 22553 9696 22558 9752
rect 22614 9696 25134 9752
rect 25190 9696 25195 9752
rect 22553 9694 25195 9696
rect 22553 9691 22619 9694
rect 25129 9691 25195 9694
rect 25865 9754 25931 9757
rect 27613 9754 27679 9757
rect 25865 9752 27679 9754
rect 25865 9696 25870 9752
rect 25926 9696 27618 9752
rect 27674 9696 27679 9752
rect 25865 9694 27679 9696
rect 25865 9691 25931 9694
rect 27613 9691 27679 9694
rect 31661 9754 31727 9757
rect 33685 9754 33751 9757
rect 31661 9752 33751 9754
rect 31661 9696 31666 9752
rect 31722 9696 33690 9752
rect 33746 9696 33751 9752
rect 31661 9694 33751 9696
rect 31661 9691 31727 9694
rect 33685 9691 33751 9694
rect 0 9618 120 9648
rect 1301 9618 1367 9621
rect 0 9616 1367 9618
rect 0 9560 1306 9616
rect 1362 9560 1367 9616
rect 0 9558 1367 9560
rect 0 9528 120 9558
rect 1301 9555 1367 9558
rect 4429 9618 4495 9621
rect 33409 9618 33475 9621
rect 4429 9616 33475 9618
rect 4429 9560 4434 9616
rect 4490 9560 33414 9616
rect 33470 9560 33475 9616
rect 4429 9558 33475 9560
rect 4429 9555 4495 9558
rect 33409 9555 33475 9558
rect 39665 9618 39731 9621
rect 40880 9618 41000 9648
rect 39665 9616 41000 9618
rect 39665 9560 39670 9616
rect 39726 9560 41000 9616
rect 39665 9558 41000 9560
rect 39665 9555 39731 9558
rect 40880 9528 41000 9558
rect 7649 9482 7715 9485
rect 15510 9482 15516 9484
rect 7649 9480 15516 9482
rect 7649 9424 7654 9480
rect 7710 9424 15516 9480
rect 7649 9422 15516 9424
rect 7649 9419 7715 9422
rect 15510 9420 15516 9422
rect 15580 9420 15586 9484
rect 15745 9482 15811 9485
rect 32438 9482 32444 9484
rect 15745 9480 32444 9482
rect 15745 9424 15750 9480
rect 15806 9424 32444 9480
rect 15745 9422 32444 9424
rect 15745 9419 15811 9422
rect 32438 9420 32444 9422
rect 32508 9420 32514 9484
rect 0 9349 120 9376
rect 0 9344 171 9349
rect 0 9288 110 9344
rect 166 9288 171 9344
rect 0 9283 171 9288
rect 7598 9284 7604 9348
rect 7668 9346 7674 9348
rect 10501 9346 10567 9349
rect 7668 9344 10567 9346
rect 7668 9288 10506 9344
rect 10562 9288 10567 9344
rect 7668 9286 10567 9288
rect 7668 9284 7674 9286
rect 10501 9283 10567 9286
rect 15561 9346 15627 9349
rect 34605 9346 34671 9349
rect 15561 9344 34671 9346
rect 15561 9288 15566 9344
rect 15622 9288 34610 9344
rect 34666 9288 34671 9344
rect 15561 9286 34671 9288
rect 15561 9283 15627 9286
rect 34605 9283 34671 9286
rect 38929 9346 38995 9349
rect 40880 9346 41000 9376
rect 38929 9344 41000 9346
rect 38929 9288 38934 9344
rect 38990 9288 41000 9344
rect 38929 9286 41000 9288
rect 38929 9283 38995 9286
rect 0 9256 120 9283
rect 40880 9256 41000 9286
rect 2497 9210 2563 9213
rect 21817 9210 21883 9213
rect 2497 9208 21883 9210
rect 2497 9152 2502 9208
rect 2558 9152 21822 9208
rect 21878 9152 21883 9208
rect 2497 9150 21883 9152
rect 2497 9147 2563 9150
rect 21817 9147 21883 9150
rect 24158 9148 24164 9212
rect 24228 9210 24234 9212
rect 27705 9210 27771 9213
rect 24228 9208 27771 9210
rect 24228 9152 27710 9208
rect 27766 9152 27771 9208
rect 24228 9150 27771 9152
rect 24228 9148 24234 9150
rect 27705 9147 27771 9150
rect 32029 9210 32095 9213
rect 35433 9210 35499 9213
rect 32029 9208 35499 9210
rect 32029 9152 32034 9208
rect 32090 9152 35438 9208
rect 35494 9152 35499 9208
rect 32029 9150 35499 9152
rect 32029 9147 32095 9150
rect 35433 9147 35499 9150
rect 0 9074 120 9104
rect 381 9074 447 9077
rect 0 9072 447 9074
rect 0 9016 386 9072
rect 442 9016 447 9072
rect 0 9014 447 9016
rect 0 8984 120 9014
rect 381 9011 447 9014
rect 3509 9074 3575 9077
rect 10133 9074 10199 9077
rect 3509 9072 10199 9074
rect 3509 9016 3514 9072
rect 3570 9016 10138 9072
rect 10194 9016 10199 9072
rect 3509 9014 10199 9016
rect 3509 9011 3575 9014
rect 10133 9011 10199 9014
rect 15193 9074 15259 9077
rect 32806 9074 32812 9076
rect 15193 9072 32812 9074
rect 15193 9016 15198 9072
rect 15254 9016 32812 9072
rect 15193 9014 32812 9016
rect 15193 9011 15259 9014
rect 32806 9012 32812 9014
rect 32876 9012 32882 9076
rect 39481 9074 39547 9077
rect 40880 9074 41000 9104
rect 39481 9072 41000 9074
rect 39481 9016 39486 9072
rect 39542 9016 41000 9072
rect 39481 9014 41000 9016
rect 39481 9011 39547 9014
rect 40880 8984 41000 9014
rect 5809 8938 5875 8941
rect 10961 8938 11027 8941
rect 17953 8938 18019 8941
rect 39389 8938 39455 8941
rect 5809 8936 11027 8938
rect 5809 8880 5814 8936
rect 5870 8880 10966 8936
rect 11022 8880 11027 8936
rect 5809 8878 11027 8880
rect 5809 8875 5875 8878
rect 10961 8875 11027 8878
rect 12390 8878 17418 8938
rect 0 8802 120 8832
rect 197 8802 263 8805
rect 0 8800 263 8802
rect 0 8744 202 8800
rect 258 8744 263 8800
rect 0 8742 263 8744
rect 0 8712 120 8742
rect 197 8739 263 8742
rect 6729 8802 6795 8805
rect 6729 8800 8816 8802
rect 6729 8744 6734 8800
rect 6790 8744 8816 8800
rect 6729 8742 8816 8744
rect 6729 8739 6795 8742
rect 3006 8736 3322 8737
rect 3006 8672 3012 8736
rect 3076 8672 3092 8736
rect 3156 8672 3172 8736
rect 3236 8672 3252 8736
rect 3316 8672 3322 8736
rect 3006 8671 3322 8672
rect 8756 8632 8816 8742
rect 9397 8800 9463 8805
rect 9397 8744 9402 8800
rect 9458 8744 9463 8800
rect 9397 8739 9463 8744
rect 9622 8740 9628 8804
rect 9692 8802 9698 8804
rect 12390 8802 12450 8878
rect 9692 8742 12450 8802
rect 17358 8802 17418 8878
rect 17953 8936 39455 8938
rect 17953 8880 17958 8936
rect 18014 8880 39394 8936
rect 39450 8880 39455 8936
rect 17953 8878 39455 8880
rect 17953 8875 18019 8878
rect 39389 8875 39455 8878
rect 18321 8802 18387 8805
rect 17358 8800 18387 8802
rect 17358 8744 18326 8800
rect 18382 8744 18387 8800
rect 17358 8742 18387 8744
rect 9692 8740 9698 8742
rect 18321 8739 18387 8742
rect 39573 8802 39639 8805
rect 40880 8802 41000 8832
rect 39573 8800 41000 8802
rect 39573 8744 39578 8800
rect 39634 8744 41000 8800
rect 39573 8742 41000 8744
rect 39573 8739 39639 8742
rect 9006 8736 9322 8737
rect 9006 8672 9012 8736
rect 9076 8672 9092 8736
rect 9156 8672 9172 8736
rect 9236 8672 9252 8736
rect 9316 8672 9322 8736
rect 9006 8671 9322 8672
rect 8756 8572 8954 8632
rect 0 8530 120 8560
rect 841 8530 907 8533
rect 0 8528 907 8530
rect 0 8472 846 8528
rect 902 8472 907 8528
rect 0 8470 907 8472
rect 0 8440 120 8470
rect 841 8467 907 8470
rect 7046 8468 7052 8532
rect 7116 8530 7122 8532
rect 8017 8530 8083 8533
rect 7116 8528 8083 8530
rect 7116 8472 8022 8528
rect 8078 8472 8083 8528
rect 7116 8470 8083 8472
rect 8894 8530 8954 8572
rect 9400 8530 9460 8739
rect 15006 8736 15322 8737
rect 15006 8672 15012 8736
rect 15076 8672 15092 8736
rect 15156 8672 15172 8736
rect 15236 8672 15252 8736
rect 15316 8672 15322 8736
rect 15006 8671 15322 8672
rect 21006 8736 21322 8737
rect 21006 8672 21012 8736
rect 21076 8672 21092 8736
rect 21156 8672 21172 8736
rect 21236 8672 21252 8736
rect 21316 8672 21322 8736
rect 21006 8671 21322 8672
rect 27006 8736 27322 8737
rect 27006 8672 27012 8736
rect 27076 8672 27092 8736
rect 27156 8672 27172 8736
rect 27236 8672 27252 8736
rect 27316 8672 27322 8736
rect 27006 8671 27322 8672
rect 33006 8736 33322 8737
rect 33006 8672 33012 8736
rect 33076 8672 33092 8736
rect 33156 8672 33172 8736
rect 33236 8672 33252 8736
rect 33316 8672 33322 8736
rect 33006 8671 33322 8672
rect 39006 8736 39322 8737
rect 39006 8672 39012 8736
rect 39076 8672 39092 8736
rect 39156 8672 39172 8736
rect 39236 8672 39252 8736
rect 39316 8672 39322 8736
rect 40880 8712 41000 8742
rect 39006 8671 39322 8672
rect 10593 8666 10659 8669
rect 14365 8666 14431 8669
rect 14733 8666 14799 8669
rect 18689 8668 18755 8669
rect 10593 8664 14799 8666
rect 10593 8608 10598 8664
rect 10654 8608 14370 8664
rect 14426 8608 14738 8664
rect 14794 8608 14799 8664
rect 10593 8606 14799 8608
rect 10593 8603 10659 8606
rect 14365 8603 14431 8606
rect 14733 8603 14799 8606
rect 18638 8604 18644 8668
rect 18708 8666 18755 8668
rect 26509 8666 26575 8669
rect 28073 8668 28139 8669
rect 28022 8666 28028 8668
rect 18708 8664 18800 8666
rect 18750 8608 18800 8664
rect 18708 8606 18800 8608
rect 23062 8664 26575 8666
rect 23062 8608 26514 8664
rect 26570 8608 26575 8664
rect 23062 8606 26575 8608
rect 27982 8606 28028 8666
rect 28092 8664 28139 8668
rect 28134 8608 28139 8664
rect 18708 8604 18755 8606
rect 18689 8603 18755 8604
rect 16798 8530 16804 8532
rect 8894 8470 9460 8530
rect 9630 8470 16804 8530
rect 7116 8468 7122 8470
rect 8017 8467 8083 8470
rect 7189 8394 7255 8397
rect 9630 8394 9690 8470
rect 16798 8468 16804 8470
rect 16868 8468 16874 8532
rect 17033 8530 17099 8533
rect 23062 8530 23122 8606
rect 26509 8603 26575 8606
rect 28022 8604 28028 8606
rect 28092 8604 28139 8608
rect 28073 8603 28139 8604
rect 28257 8666 28323 8669
rect 28901 8666 28967 8669
rect 28257 8664 28967 8666
rect 28257 8608 28262 8664
rect 28318 8608 28906 8664
rect 28962 8608 28967 8664
rect 28257 8606 28967 8608
rect 28257 8603 28323 8606
rect 28901 8603 28967 8606
rect 29085 8666 29151 8669
rect 29821 8666 29887 8669
rect 29085 8664 29887 8666
rect 29085 8608 29090 8664
rect 29146 8608 29826 8664
rect 29882 8608 29887 8664
rect 29085 8606 29887 8608
rect 29085 8603 29151 8606
rect 29821 8603 29887 8606
rect 30925 8666 30991 8669
rect 32857 8666 32923 8669
rect 30925 8664 32923 8666
rect 30925 8608 30930 8664
rect 30986 8608 32862 8664
rect 32918 8608 32923 8664
rect 30925 8606 32923 8608
rect 30925 8603 30991 8606
rect 32857 8603 32923 8606
rect 17033 8528 23122 8530
rect 17033 8472 17038 8528
rect 17094 8472 23122 8528
rect 17033 8470 23122 8472
rect 23289 8530 23355 8533
rect 24485 8530 24551 8533
rect 23289 8528 24551 8530
rect 23289 8472 23294 8528
rect 23350 8472 24490 8528
rect 24546 8472 24551 8528
rect 23289 8470 24551 8472
rect 17033 8467 17099 8470
rect 23289 8467 23355 8470
rect 24485 8467 24551 8470
rect 25221 8532 25287 8533
rect 25221 8528 25268 8532
rect 25332 8530 25338 8532
rect 25221 8472 25226 8528
rect 25221 8468 25268 8472
rect 25332 8470 25378 8530
rect 25332 8468 25338 8470
rect 26550 8468 26556 8532
rect 26620 8530 26626 8532
rect 26785 8530 26851 8533
rect 32029 8530 32095 8533
rect 26620 8528 26851 8530
rect 26620 8472 26790 8528
rect 26846 8472 26851 8528
rect 26620 8470 26851 8472
rect 26620 8468 26626 8470
rect 25221 8467 25287 8468
rect 26785 8467 26851 8470
rect 27110 8528 32095 8530
rect 27110 8472 32034 8528
rect 32090 8472 32095 8528
rect 27110 8470 32095 8472
rect 7189 8392 9690 8394
rect 7189 8336 7194 8392
rect 7250 8336 9690 8392
rect 7189 8334 9690 8336
rect 13537 8394 13603 8397
rect 17902 8394 17908 8396
rect 13537 8392 17908 8394
rect 13537 8336 13542 8392
rect 13598 8336 17908 8392
rect 13537 8334 17908 8336
rect 7189 8331 7255 8334
rect 13537 8331 13603 8334
rect 17902 8332 17908 8334
rect 17972 8332 17978 8396
rect 18045 8394 18111 8397
rect 18045 8392 26802 8394
rect 18045 8336 18050 8392
rect 18106 8336 26802 8392
rect 18045 8334 26802 8336
rect 18045 8331 18111 8334
rect 0 8258 120 8288
rect 1117 8258 1183 8261
rect 7741 8260 7807 8261
rect 7741 8258 7788 8260
rect 0 8256 1183 8258
rect 0 8200 1122 8256
rect 1178 8200 1183 8256
rect 0 8198 1183 8200
rect 7696 8256 7788 8258
rect 7696 8200 7746 8256
rect 7696 8198 7788 8200
rect 0 8168 120 8198
rect 1117 8195 1183 8198
rect 7741 8196 7788 8198
rect 7852 8196 7858 8260
rect 8385 8258 8451 8261
rect 8518 8258 8524 8260
rect 8385 8256 8524 8258
rect 8385 8200 8390 8256
rect 8446 8200 8524 8256
rect 8385 8198 8524 8200
rect 7741 8195 7807 8196
rect 8385 8195 8451 8198
rect 8518 8196 8524 8198
rect 8588 8196 8594 8260
rect 8661 8258 8727 8261
rect 10869 8258 10935 8261
rect 8661 8256 10935 8258
rect 8661 8200 8666 8256
rect 8722 8200 10874 8256
rect 10930 8200 10935 8256
rect 8661 8198 10935 8200
rect 8661 8195 8727 8198
rect 10869 8195 10935 8198
rect 14733 8258 14799 8261
rect 19425 8258 19491 8261
rect 14733 8256 19491 8258
rect 14733 8200 14738 8256
rect 14794 8200 19430 8256
rect 19486 8200 19491 8256
rect 14733 8198 19491 8200
rect 14733 8195 14799 8198
rect 19425 8195 19491 8198
rect 23105 8258 23171 8261
rect 24117 8258 24183 8261
rect 23105 8256 24183 8258
rect 23105 8200 23110 8256
rect 23166 8200 24122 8256
rect 24178 8200 24183 8256
rect 23105 8198 24183 8200
rect 23105 8195 23171 8198
rect 24117 8195 24183 8198
rect 25446 8196 25452 8260
rect 25516 8258 25522 8260
rect 25773 8258 25839 8261
rect 25516 8256 25839 8258
rect 25516 8200 25778 8256
rect 25834 8200 25839 8256
rect 25516 8198 25839 8200
rect 26742 8258 26802 8334
rect 27110 8258 27170 8470
rect 32029 8467 32095 8470
rect 32397 8530 32463 8533
rect 32949 8530 33015 8533
rect 32397 8528 33015 8530
rect 32397 8472 32402 8528
rect 32458 8472 32954 8528
rect 33010 8472 33015 8528
rect 32397 8470 33015 8472
rect 32397 8467 32463 8470
rect 32949 8467 33015 8470
rect 38653 8530 38719 8533
rect 40880 8530 41000 8560
rect 38653 8528 41000 8530
rect 38653 8472 38658 8528
rect 38714 8472 41000 8528
rect 38653 8470 41000 8472
rect 38653 8467 38719 8470
rect 40880 8440 41000 8470
rect 27705 8394 27771 8397
rect 38837 8394 38903 8397
rect 27705 8392 38903 8394
rect 27705 8336 27710 8392
rect 27766 8336 38842 8392
rect 38898 8336 38903 8392
rect 27705 8334 38903 8336
rect 27705 8331 27771 8334
rect 38837 8331 38903 8334
rect 26742 8198 27170 8258
rect 27705 8258 27771 8261
rect 28165 8258 28231 8261
rect 28901 8258 28967 8261
rect 27705 8256 28044 8258
rect 27705 8200 27710 8256
rect 27766 8200 28044 8256
rect 27705 8198 28044 8200
rect 25516 8196 25522 8198
rect 25773 8195 25839 8198
rect 27705 8195 27771 8198
rect 1946 8192 2262 8193
rect 1946 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2262 8192
rect 1946 8127 2262 8128
rect 7946 8192 8262 8193
rect 7946 8128 7952 8192
rect 8016 8128 8032 8192
rect 8096 8128 8112 8192
rect 8176 8128 8192 8192
rect 8256 8128 8262 8192
rect 7946 8127 8262 8128
rect 13946 8192 14262 8193
rect 13946 8128 13952 8192
rect 14016 8128 14032 8192
rect 14096 8128 14112 8192
rect 14176 8128 14192 8192
rect 14256 8128 14262 8192
rect 13946 8127 14262 8128
rect 19946 8192 20262 8193
rect 19946 8128 19952 8192
rect 20016 8128 20032 8192
rect 20096 8128 20112 8192
rect 20176 8128 20192 8192
rect 20256 8128 20262 8192
rect 19946 8127 20262 8128
rect 25946 8192 26262 8193
rect 25946 8128 25952 8192
rect 26016 8128 26032 8192
rect 26096 8128 26112 8192
rect 26176 8128 26192 8192
rect 26256 8128 26262 8192
rect 25946 8127 26262 8128
rect 2589 8122 2655 8125
rect 7649 8122 7715 8125
rect 12525 8122 12591 8125
rect 2589 8120 7715 8122
rect 2589 8064 2594 8120
rect 2650 8064 7654 8120
rect 7710 8064 7715 8120
rect 2589 8062 7715 8064
rect 2589 8059 2655 8062
rect 7649 8059 7715 8062
rect 8342 8120 12591 8122
rect 8342 8064 12530 8120
rect 12586 8064 12591 8120
rect 8342 8062 12591 8064
rect 0 7986 120 8016
rect 1209 7986 1275 7989
rect 0 7984 1275 7986
rect 0 7928 1214 7984
rect 1270 7928 1275 7984
rect 0 7926 1275 7928
rect 0 7896 120 7926
rect 1209 7923 1275 7926
rect 7005 7986 7071 7989
rect 8342 7986 8402 8062
rect 12525 8059 12591 8062
rect 14825 8122 14891 8125
rect 15653 8122 15719 8125
rect 14825 8120 15719 8122
rect 14825 8064 14830 8120
rect 14886 8064 15658 8120
rect 15714 8064 15719 8120
rect 14825 8062 15719 8064
rect 14825 8059 14891 8062
rect 15653 8059 15719 8062
rect 16297 8122 16363 8125
rect 17953 8122 18019 8125
rect 16297 8120 18019 8122
rect 16297 8064 16302 8120
rect 16358 8064 17958 8120
rect 18014 8064 18019 8120
rect 16297 8062 18019 8064
rect 16297 8059 16363 8062
rect 17953 8059 18019 8062
rect 18137 8122 18203 8125
rect 18454 8122 18460 8124
rect 18137 8120 18460 8122
rect 18137 8064 18142 8120
rect 18198 8064 18460 8120
rect 18137 8062 18460 8064
rect 18137 8059 18203 8062
rect 18454 8060 18460 8062
rect 18524 8060 18530 8124
rect 18873 8122 18939 8125
rect 19057 8124 19123 8125
rect 19006 8122 19012 8124
rect 18873 8120 19012 8122
rect 19076 8122 19123 8124
rect 25630 8122 25636 8124
rect 19076 8120 19204 8122
rect 18873 8064 18878 8120
rect 18934 8064 19012 8120
rect 19118 8064 19204 8120
rect 18873 8062 19012 8064
rect 18873 8059 18939 8062
rect 19006 8060 19012 8062
rect 19076 8062 19204 8064
rect 20486 8062 25636 8122
rect 19076 8060 19123 8062
rect 19057 8059 19123 8060
rect 7005 7984 8402 7986
rect 7005 7928 7010 7984
rect 7066 7928 8402 7984
rect 7005 7926 8402 7928
rect 8569 7986 8635 7989
rect 13629 7986 13695 7989
rect 8569 7984 13695 7986
rect 8569 7928 8574 7984
rect 8630 7928 13634 7984
rect 13690 7928 13695 7984
rect 8569 7926 13695 7928
rect 7005 7923 7071 7926
rect 8569 7923 8635 7926
rect 13629 7923 13695 7926
rect 14549 7986 14615 7989
rect 20486 7986 20546 8062
rect 25630 8060 25636 8062
rect 25700 8060 25706 8124
rect 26366 8060 26372 8124
rect 26436 8122 26442 8124
rect 27797 8122 27863 8125
rect 26436 8120 27863 8122
rect 26436 8064 27802 8120
rect 27858 8064 27863 8120
rect 26436 8062 27863 8064
rect 27984 8122 28044 8198
rect 28165 8256 28967 8258
rect 28165 8200 28170 8256
rect 28226 8200 28906 8256
rect 28962 8200 28967 8256
rect 28165 8198 28967 8200
rect 28165 8195 28231 8198
rect 28901 8195 28967 8198
rect 32397 8258 32463 8261
rect 33225 8258 33291 8261
rect 32397 8256 33291 8258
rect 32397 8200 32402 8256
rect 32458 8200 33230 8256
rect 33286 8200 33291 8256
rect 32397 8198 33291 8200
rect 32397 8195 32463 8198
rect 33225 8195 33291 8198
rect 39021 8258 39087 8261
rect 40880 8258 41000 8288
rect 39021 8256 41000 8258
rect 39021 8200 39026 8256
rect 39082 8200 41000 8256
rect 39021 8198 41000 8200
rect 39021 8195 39087 8198
rect 31946 8192 32262 8193
rect 31946 8128 31952 8192
rect 32016 8128 32032 8192
rect 32096 8128 32112 8192
rect 32176 8128 32192 8192
rect 32256 8128 32262 8192
rect 31946 8127 32262 8128
rect 37946 8192 38262 8193
rect 37946 8128 37952 8192
rect 38016 8128 38032 8192
rect 38096 8128 38112 8192
rect 38176 8128 38192 8192
rect 38256 8128 38262 8192
rect 40880 8168 41000 8198
rect 37946 8127 38262 8128
rect 28717 8122 28783 8125
rect 27984 8120 28783 8122
rect 27984 8064 28722 8120
rect 28778 8064 28783 8120
rect 27984 8062 28783 8064
rect 26436 8060 26442 8062
rect 27797 8059 27863 8062
rect 28717 8059 28783 8062
rect 30465 8122 30531 8125
rect 30598 8122 30604 8124
rect 30465 8120 30604 8122
rect 30465 8064 30470 8120
rect 30526 8064 30604 8120
rect 30465 8062 30604 8064
rect 30465 8059 30531 8062
rect 30598 8060 30604 8062
rect 30668 8060 30674 8124
rect 32622 8060 32628 8124
rect 32692 8122 32698 8124
rect 32765 8122 32831 8125
rect 32692 8120 32831 8122
rect 32692 8064 32770 8120
rect 32826 8064 32831 8120
rect 32692 8062 32831 8064
rect 32692 8060 32698 8062
rect 32765 8059 32831 8062
rect 14549 7984 20546 7986
rect 14549 7928 14554 7984
rect 14610 7928 20546 7984
rect 14549 7926 20546 7928
rect 20989 7986 21055 7989
rect 28717 7986 28783 7989
rect 20989 7984 28783 7986
rect 20989 7928 20994 7984
rect 21050 7928 28722 7984
rect 28778 7928 28783 7984
rect 20989 7926 28783 7928
rect 14549 7923 14615 7926
rect 20989 7923 21055 7926
rect 28717 7923 28783 7926
rect 30281 7986 30347 7989
rect 32857 7986 32923 7989
rect 30281 7984 32923 7986
rect 30281 7928 30286 7984
rect 30342 7928 32862 7984
rect 32918 7928 32923 7984
rect 30281 7926 32923 7928
rect 30281 7923 30347 7926
rect 32857 7923 32923 7926
rect 39389 7986 39455 7989
rect 40880 7986 41000 8016
rect 39389 7984 41000 7986
rect 39389 7928 39394 7984
rect 39450 7928 41000 7984
rect 39389 7926 41000 7928
rect 39389 7923 39455 7926
rect 40880 7896 41000 7926
rect 2589 7850 2655 7853
rect 6913 7850 6979 7853
rect 2589 7848 3802 7850
rect 2589 7792 2594 7848
rect 2650 7792 3802 7848
rect 2589 7790 3802 7792
rect 2589 7787 2655 7790
rect 0 7714 120 7744
rect 749 7714 815 7717
rect 0 7712 815 7714
rect 0 7656 754 7712
rect 810 7656 815 7712
rect 0 7654 815 7656
rect 0 7624 120 7654
rect 749 7651 815 7654
rect 3006 7648 3322 7649
rect 3006 7584 3012 7648
rect 3076 7584 3092 7648
rect 3156 7584 3172 7648
rect 3236 7584 3252 7648
rect 3316 7584 3322 7648
rect 3006 7583 3322 7584
rect 3742 7578 3802 7790
rect 6913 7848 9506 7850
rect 6913 7792 6918 7848
rect 6974 7792 9506 7848
rect 6913 7790 9506 7792
rect 6913 7787 6979 7790
rect 3969 7714 4035 7717
rect 8569 7714 8635 7717
rect 3969 7712 8635 7714
rect 3969 7656 3974 7712
rect 4030 7656 8574 7712
rect 8630 7656 8635 7712
rect 3969 7654 8635 7656
rect 9446 7714 9506 7790
rect 10910 7788 10916 7852
rect 10980 7850 10986 7852
rect 33593 7850 33659 7853
rect 10980 7848 33659 7850
rect 10980 7792 33598 7848
rect 33654 7792 33659 7848
rect 10980 7790 33659 7792
rect 10980 7788 10986 7790
rect 33593 7787 33659 7790
rect 12709 7714 12775 7717
rect 13721 7714 13787 7717
rect 14825 7714 14891 7717
rect 9446 7654 12450 7714
rect 3969 7651 4035 7654
rect 8569 7651 8635 7654
rect 9006 7648 9322 7649
rect 9006 7584 9012 7648
rect 9076 7584 9092 7648
rect 9156 7584 9172 7648
rect 9236 7584 9252 7648
rect 9316 7584 9322 7648
rect 9006 7583 9322 7584
rect 8661 7578 8727 7581
rect 10317 7580 10383 7581
rect 10317 7578 10364 7580
rect 3742 7576 8727 7578
rect 3742 7520 8666 7576
rect 8722 7520 8727 7576
rect 3742 7518 8727 7520
rect 10272 7576 10364 7578
rect 10272 7520 10322 7576
rect 10272 7518 10364 7520
rect 8661 7515 8727 7518
rect 10317 7516 10364 7518
rect 10428 7516 10434 7580
rect 12390 7578 12450 7654
rect 12709 7712 14891 7714
rect 12709 7656 12714 7712
rect 12770 7656 13726 7712
rect 13782 7656 14830 7712
rect 14886 7656 14891 7712
rect 12709 7654 14891 7656
rect 12709 7651 12775 7654
rect 13721 7651 13787 7654
rect 14825 7651 14891 7654
rect 16021 7714 16087 7717
rect 16665 7714 16731 7717
rect 16021 7712 16731 7714
rect 16021 7656 16026 7712
rect 16082 7656 16670 7712
rect 16726 7656 16731 7712
rect 16021 7654 16731 7656
rect 16021 7651 16087 7654
rect 16665 7651 16731 7654
rect 17953 7714 18019 7717
rect 20805 7714 20871 7717
rect 17953 7712 20871 7714
rect 17953 7656 17958 7712
rect 18014 7656 20810 7712
rect 20866 7656 20871 7712
rect 17953 7654 20871 7656
rect 17953 7651 18019 7654
rect 20805 7651 20871 7654
rect 22461 7714 22527 7717
rect 23565 7714 23631 7717
rect 22461 7712 23631 7714
rect 22461 7656 22466 7712
rect 22522 7656 23570 7712
rect 23626 7656 23631 7712
rect 22461 7654 23631 7656
rect 22461 7651 22527 7654
rect 23565 7651 23631 7654
rect 23933 7714 23999 7717
rect 25865 7714 25931 7717
rect 23933 7712 25931 7714
rect 23933 7656 23938 7712
rect 23994 7656 25870 7712
rect 25926 7656 25931 7712
rect 23933 7654 25931 7656
rect 23933 7651 23999 7654
rect 25865 7651 25931 7654
rect 28533 7714 28599 7717
rect 30281 7714 30347 7717
rect 32213 7714 32279 7717
rect 28533 7712 30347 7714
rect 28533 7656 28538 7712
rect 28594 7656 30286 7712
rect 30342 7656 30347 7712
rect 28533 7654 30347 7656
rect 28533 7651 28599 7654
rect 30281 7651 30347 7654
rect 30606 7712 32279 7714
rect 30606 7656 32218 7712
rect 32274 7656 32279 7712
rect 30606 7654 32279 7656
rect 15006 7648 15322 7649
rect 15006 7584 15012 7648
rect 15076 7584 15092 7648
rect 15156 7584 15172 7648
rect 15236 7584 15252 7648
rect 15316 7584 15322 7648
rect 15006 7583 15322 7584
rect 21006 7648 21322 7649
rect 21006 7584 21012 7648
rect 21076 7584 21092 7648
rect 21156 7584 21172 7648
rect 21236 7584 21252 7648
rect 21316 7584 21322 7648
rect 21006 7583 21322 7584
rect 27006 7648 27322 7649
rect 27006 7584 27012 7648
rect 27076 7584 27092 7648
rect 27156 7584 27172 7648
rect 27236 7584 27252 7648
rect 27316 7584 27322 7648
rect 27006 7583 27322 7584
rect 20713 7578 20779 7581
rect 12390 7518 14842 7578
rect 10317 7515 10383 7516
rect 0 7442 120 7472
rect 749 7442 815 7445
rect 0 7440 815 7442
rect 0 7384 754 7440
rect 810 7384 815 7440
rect 0 7382 815 7384
rect 0 7352 120 7382
rect 749 7379 815 7382
rect 5165 7442 5231 7445
rect 6361 7442 6427 7445
rect 5165 7440 6427 7442
rect 5165 7384 5170 7440
rect 5226 7384 6366 7440
rect 6422 7384 6427 7440
rect 5165 7382 6427 7384
rect 5165 7379 5231 7382
rect 6361 7379 6427 7382
rect 7925 7442 7991 7445
rect 14549 7442 14615 7445
rect 7925 7440 14615 7442
rect 7925 7384 7930 7440
rect 7986 7384 14554 7440
rect 14610 7384 14615 7440
rect 7925 7382 14615 7384
rect 14782 7442 14842 7518
rect 15518 7576 20779 7578
rect 15518 7520 20718 7576
rect 20774 7520 20779 7576
rect 15518 7518 20779 7520
rect 15518 7442 15578 7518
rect 20713 7515 20779 7518
rect 21449 7578 21515 7581
rect 24209 7578 24275 7581
rect 21449 7576 24275 7578
rect 21449 7520 21454 7576
rect 21510 7520 24214 7576
rect 24270 7520 24275 7576
rect 21449 7518 24275 7520
rect 21449 7515 21515 7518
rect 24209 7515 24275 7518
rect 29729 7578 29795 7581
rect 30606 7578 30666 7654
rect 32213 7651 32279 7654
rect 39389 7714 39455 7717
rect 40880 7714 41000 7744
rect 39389 7712 41000 7714
rect 39389 7656 39394 7712
rect 39450 7656 41000 7712
rect 39389 7654 41000 7656
rect 39389 7651 39455 7654
rect 33006 7648 33322 7649
rect 33006 7584 33012 7648
rect 33076 7584 33092 7648
rect 33156 7584 33172 7648
rect 33236 7584 33252 7648
rect 33316 7584 33322 7648
rect 33006 7583 33322 7584
rect 39006 7648 39322 7649
rect 39006 7584 39012 7648
rect 39076 7584 39092 7648
rect 39156 7584 39172 7648
rect 39236 7584 39252 7648
rect 39316 7584 39322 7648
rect 40880 7624 41000 7654
rect 39006 7583 39322 7584
rect 29729 7576 30666 7578
rect 29729 7520 29734 7576
rect 29790 7520 30666 7576
rect 29729 7518 30666 7520
rect 29729 7515 29795 7518
rect 31334 7516 31340 7580
rect 31404 7578 31410 7580
rect 32622 7578 32628 7580
rect 31404 7518 32628 7578
rect 31404 7516 31410 7518
rect 32622 7516 32628 7518
rect 32692 7516 32698 7580
rect 14782 7382 15578 7442
rect 15929 7442 15995 7445
rect 32949 7442 33015 7445
rect 15929 7440 33015 7442
rect 15929 7384 15934 7440
rect 15990 7384 32954 7440
rect 33010 7384 33015 7440
rect 15929 7382 33015 7384
rect 7925 7379 7991 7382
rect 14549 7379 14615 7382
rect 15929 7379 15995 7382
rect 32949 7379 33015 7382
rect 38929 7442 38995 7445
rect 40880 7442 41000 7472
rect 38929 7440 41000 7442
rect 38929 7384 38934 7440
rect 38990 7384 41000 7440
rect 38929 7382 41000 7384
rect 38929 7379 38995 7382
rect 40880 7352 41000 7382
rect 7005 7306 7071 7309
rect 8477 7306 8543 7309
rect 7005 7304 8543 7306
rect 7005 7248 7010 7304
rect 7066 7248 8482 7304
rect 8538 7248 8543 7304
rect 7005 7246 8543 7248
rect 7005 7243 7071 7246
rect 8477 7243 8543 7246
rect 8702 7244 8708 7308
rect 8772 7306 8778 7308
rect 20713 7306 20779 7309
rect 33225 7306 33291 7309
rect 8772 7246 20546 7306
rect 8772 7244 8778 7246
rect 0 7170 120 7200
rect 749 7170 815 7173
rect 0 7168 815 7170
rect 0 7112 754 7168
rect 810 7112 815 7168
rect 0 7110 815 7112
rect 0 7080 120 7110
rect 749 7107 815 7110
rect 4429 7170 4495 7173
rect 4429 7168 7850 7170
rect 4429 7112 4434 7168
rect 4490 7112 7850 7168
rect 4429 7110 7850 7112
rect 4429 7107 4495 7110
rect 1946 7104 2262 7105
rect 1946 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2262 7104
rect 1946 7039 2262 7040
rect 3233 7034 3299 7037
rect 3918 7034 3924 7036
rect 3233 7032 3924 7034
rect 3233 6976 3238 7032
rect 3294 6976 3924 7032
rect 3233 6974 3924 6976
rect 3233 6971 3299 6974
rect 3918 6972 3924 6974
rect 3988 6972 3994 7036
rect 6678 6972 6684 7036
rect 6748 7034 6754 7036
rect 6821 7034 6887 7037
rect 6748 7032 6887 7034
rect 6748 6976 6826 7032
rect 6882 6976 6887 7032
rect 6748 6974 6887 6976
rect 6748 6972 6754 6974
rect 6821 6971 6887 6974
rect 0 6898 120 6928
rect 1025 6898 1091 6901
rect 0 6896 1091 6898
rect 0 6840 1030 6896
rect 1086 6840 1091 6896
rect 0 6838 1091 6840
rect 0 6808 120 6838
rect 1025 6835 1091 6838
rect 3233 6898 3299 6901
rect 5625 6898 5691 6901
rect 3233 6896 5691 6898
rect 3233 6840 3238 6896
rect 3294 6840 5630 6896
rect 5686 6840 5691 6896
rect 3233 6838 5691 6840
rect 7790 6898 7850 7110
rect 8518 7108 8524 7172
rect 8588 7170 8594 7172
rect 13169 7170 13235 7173
rect 8588 7168 13235 7170
rect 8588 7112 13174 7168
rect 13230 7112 13235 7168
rect 8588 7110 13235 7112
rect 8588 7108 8594 7110
rect 13169 7107 13235 7110
rect 14774 7108 14780 7172
rect 14844 7170 14850 7172
rect 16021 7170 16087 7173
rect 14844 7168 16087 7170
rect 14844 7112 16026 7168
rect 16082 7112 16087 7168
rect 14844 7110 16087 7112
rect 14844 7108 14850 7110
rect 16021 7107 16087 7110
rect 16246 7108 16252 7172
rect 16316 7170 16322 7172
rect 18505 7170 18571 7173
rect 16316 7168 18571 7170
rect 16316 7112 18510 7168
rect 18566 7112 18571 7168
rect 16316 7110 18571 7112
rect 16316 7108 16322 7110
rect 18505 7107 18571 7110
rect 7946 7104 8262 7105
rect 7946 7040 7952 7104
rect 8016 7040 8032 7104
rect 8096 7040 8112 7104
rect 8176 7040 8192 7104
rect 8256 7040 8262 7104
rect 7946 7039 8262 7040
rect 13946 7104 14262 7105
rect 13946 7040 13952 7104
rect 14016 7040 14032 7104
rect 14096 7040 14112 7104
rect 14176 7040 14192 7104
rect 14256 7040 14262 7104
rect 13946 7039 14262 7040
rect 19946 7104 20262 7105
rect 19946 7040 19952 7104
rect 20016 7040 20032 7104
rect 20096 7040 20112 7104
rect 20176 7040 20192 7104
rect 20256 7040 20262 7104
rect 19946 7039 20262 7040
rect 12341 7034 12407 7037
rect 15929 7036 15995 7037
rect 8342 7032 12407 7034
rect 8342 6976 12346 7032
rect 12402 6976 12407 7032
rect 8342 6974 12407 6976
rect 8342 6898 8402 6974
rect 12341 6971 12407 6974
rect 15878 6972 15884 7036
rect 15948 7034 15995 7036
rect 15948 7032 16040 7034
rect 15990 6976 16040 7032
rect 15948 6974 16040 6976
rect 15948 6972 15995 6974
rect 18638 6972 18644 7036
rect 18708 7034 18714 7036
rect 18781 7034 18847 7037
rect 18708 7032 18847 7034
rect 18708 6976 18786 7032
rect 18842 6976 18847 7032
rect 18708 6974 18847 6976
rect 20486 7034 20546 7246
rect 20713 7304 33291 7306
rect 20713 7248 20718 7304
rect 20774 7248 33230 7304
rect 33286 7248 33291 7304
rect 20713 7246 33291 7248
rect 20713 7243 20779 7246
rect 33225 7243 33291 7246
rect 20805 7170 20871 7173
rect 24117 7170 24183 7173
rect 20805 7168 24183 7170
rect 20805 7112 20810 7168
rect 20866 7112 24122 7168
rect 24178 7112 24183 7168
rect 20805 7110 24183 7112
rect 20805 7107 20871 7110
rect 24117 7107 24183 7110
rect 26417 7170 26483 7173
rect 28533 7170 28599 7173
rect 26417 7168 28599 7170
rect 26417 7112 26422 7168
rect 26478 7112 28538 7168
rect 28594 7112 28599 7168
rect 26417 7110 28599 7112
rect 26417 7107 26483 7110
rect 28533 7107 28599 7110
rect 29361 7170 29427 7173
rect 31753 7170 31819 7173
rect 29361 7168 31819 7170
rect 29361 7112 29366 7168
rect 29422 7112 31758 7168
rect 31814 7112 31819 7168
rect 29361 7110 31819 7112
rect 29361 7107 29427 7110
rect 31753 7107 31819 7110
rect 39389 7170 39455 7173
rect 40880 7170 41000 7200
rect 39389 7168 41000 7170
rect 39389 7112 39394 7168
rect 39450 7112 41000 7168
rect 39389 7110 41000 7112
rect 39389 7107 39455 7110
rect 25946 7104 26262 7105
rect 25946 7040 25952 7104
rect 26016 7040 26032 7104
rect 26096 7040 26112 7104
rect 26176 7040 26192 7104
rect 26256 7040 26262 7104
rect 25946 7039 26262 7040
rect 31946 7104 32262 7105
rect 31946 7040 31952 7104
rect 32016 7040 32032 7104
rect 32096 7040 32112 7104
rect 32176 7040 32192 7104
rect 32256 7040 32262 7104
rect 31946 7039 32262 7040
rect 37946 7104 38262 7105
rect 37946 7040 37952 7104
rect 38016 7040 38032 7104
rect 38096 7040 38112 7104
rect 38176 7040 38192 7104
rect 38256 7040 38262 7104
rect 40880 7080 41000 7110
rect 37946 7039 38262 7040
rect 25773 7034 25839 7037
rect 20486 7032 25839 7034
rect 20486 6976 25778 7032
rect 25834 6976 25839 7032
rect 20486 6974 25839 6976
rect 18708 6972 18714 6974
rect 15929 6971 15995 6972
rect 18781 6971 18847 6974
rect 25773 6971 25839 6974
rect 26734 6972 26740 7036
rect 26804 7034 26810 7036
rect 26877 7034 26943 7037
rect 26804 7032 26943 7034
rect 26804 6976 26882 7032
rect 26938 6976 26943 7032
rect 26804 6974 26943 6976
rect 26804 6972 26810 6974
rect 26877 6971 26943 6974
rect 27153 7034 27219 7037
rect 27429 7034 27495 7037
rect 29177 7034 29243 7037
rect 31753 7034 31819 7037
rect 27153 7032 29010 7034
rect 27153 6976 27158 7032
rect 27214 6976 27434 7032
rect 27490 6976 29010 7032
rect 27153 6974 29010 6976
rect 27153 6971 27219 6974
rect 27429 6971 27495 6974
rect 7790 6838 8402 6898
rect 8477 6898 8543 6901
rect 11237 6898 11303 6901
rect 8477 6896 11303 6898
rect 8477 6840 8482 6896
rect 8538 6840 11242 6896
rect 11298 6840 11303 6896
rect 8477 6838 11303 6840
rect 3233 6835 3299 6838
rect 5625 6835 5691 6838
rect 8477 6835 8543 6838
rect 11237 6835 11303 6838
rect 13629 6898 13695 6901
rect 16665 6898 16731 6901
rect 13629 6896 16731 6898
rect 13629 6840 13634 6896
rect 13690 6840 16670 6896
rect 16726 6840 16731 6896
rect 13629 6838 16731 6840
rect 13629 6835 13695 6838
rect 16665 6835 16731 6838
rect 17401 6898 17467 6901
rect 18505 6898 18571 6901
rect 17401 6896 18571 6898
rect 17401 6840 17406 6896
rect 17462 6840 18510 6896
rect 18566 6840 18571 6896
rect 17401 6838 18571 6840
rect 17401 6835 17467 6838
rect 18505 6835 18571 6838
rect 19057 6898 19123 6901
rect 20437 6898 20503 6901
rect 23473 6900 23539 6901
rect 19057 6896 20503 6898
rect 19057 6840 19062 6896
rect 19118 6840 20442 6896
rect 20498 6840 20503 6896
rect 19057 6838 20503 6840
rect 19057 6835 19123 6838
rect 20437 6835 20503 6838
rect 23422 6836 23428 6900
rect 23492 6898 23539 6900
rect 23492 6896 23584 6898
rect 23534 6840 23584 6896
rect 23492 6838 23584 6840
rect 23492 6836 23539 6838
rect 25630 6836 25636 6900
rect 25700 6898 25706 6900
rect 28950 6898 29010 6974
rect 29177 7032 31819 7034
rect 29177 6976 29182 7032
rect 29238 6976 31758 7032
rect 31814 6976 31819 7032
rect 29177 6974 31819 6976
rect 29177 6971 29243 6974
rect 31753 6971 31819 6974
rect 32949 6898 33015 6901
rect 25700 6838 27538 6898
rect 28950 6896 33015 6898
rect 28950 6840 32954 6896
rect 33010 6840 33015 6896
rect 28950 6838 33015 6840
rect 25700 6836 25706 6838
rect 23473 6835 23539 6836
rect 3233 6762 3299 6765
rect 4245 6762 4311 6765
rect 18505 6762 18571 6765
rect 24301 6762 24367 6765
rect 25681 6762 25747 6765
rect 3233 6760 4170 6762
rect 3233 6704 3238 6760
rect 3294 6704 4170 6760
rect 3233 6702 4170 6704
rect 3233 6699 3299 6702
rect 0 6626 120 6656
rect 933 6626 999 6629
rect 0 6624 999 6626
rect 0 6568 938 6624
rect 994 6568 999 6624
rect 0 6566 999 6568
rect 4110 6626 4170 6702
rect 4245 6760 18571 6762
rect 4245 6704 4250 6760
rect 4306 6704 18510 6760
rect 18566 6704 18571 6760
rect 4245 6702 18571 6704
rect 4245 6699 4311 6702
rect 18505 6699 18571 6702
rect 18830 6702 24226 6762
rect 4889 6626 4955 6629
rect 5441 6628 5507 6629
rect 5390 6626 5396 6628
rect 4110 6624 4955 6626
rect 4110 6568 4894 6624
rect 4950 6568 4955 6624
rect 4110 6566 4955 6568
rect 5350 6566 5396 6626
rect 5460 6624 5507 6628
rect 8477 6626 8543 6629
rect 13169 6626 13235 6629
rect 5502 6568 5507 6624
rect 0 6536 120 6566
rect 933 6563 999 6566
rect 4889 6563 4955 6566
rect 5390 6564 5396 6566
rect 5460 6564 5507 6568
rect 5441 6563 5507 6564
rect 5582 6624 8543 6626
rect 5582 6568 8482 6624
rect 8538 6568 8543 6624
rect 5582 6566 8543 6568
rect 3006 6560 3322 6561
rect 3006 6496 3012 6560
rect 3076 6496 3092 6560
rect 3156 6496 3172 6560
rect 3236 6496 3252 6560
rect 3316 6496 3322 6560
rect 3006 6495 3322 6496
rect 5165 6490 5231 6493
rect 5441 6490 5507 6493
rect 5165 6488 5507 6490
rect 5165 6432 5170 6488
rect 5226 6432 5446 6488
rect 5502 6432 5507 6488
rect 5165 6430 5507 6432
rect 5165 6427 5231 6430
rect 5441 6427 5507 6430
rect 0 6354 120 6384
rect 289 6354 355 6357
rect 0 6352 355 6354
rect 0 6296 294 6352
rect 350 6296 355 6352
rect 0 6294 355 6296
rect 0 6264 120 6294
rect 289 6291 355 6294
rect 2221 6354 2287 6357
rect 2446 6354 2452 6356
rect 2221 6352 2452 6354
rect 2221 6296 2226 6352
rect 2282 6296 2452 6352
rect 2221 6294 2452 6296
rect 2221 6291 2287 6294
rect 2446 6292 2452 6294
rect 2516 6292 2522 6356
rect 2681 6354 2747 6357
rect 5582 6354 5642 6566
rect 8477 6563 8543 6566
rect 12390 6624 13235 6626
rect 12390 6568 13174 6624
rect 13230 6568 13235 6624
rect 12390 6566 13235 6568
rect 9006 6560 9322 6561
rect 9006 6496 9012 6560
rect 9076 6496 9092 6560
rect 9156 6496 9172 6560
rect 9236 6496 9252 6560
rect 9316 6496 9322 6560
rect 9006 6495 9322 6496
rect 5809 6490 5875 6493
rect 8753 6490 8819 6493
rect 12390 6490 12450 6566
rect 13169 6563 13235 6566
rect 16665 6626 16731 6629
rect 17861 6626 17927 6629
rect 16665 6624 17927 6626
rect 16665 6568 16670 6624
rect 16726 6568 17866 6624
rect 17922 6568 17927 6624
rect 16665 6566 17927 6568
rect 16665 6563 16731 6566
rect 17861 6563 17927 6566
rect 18321 6626 18387 6629
rect 18597 6626 18663 6629
rect 18321 6624 18663 6626
rect 18321 6568 18326 6624
rect 18382 6568 18602 6624
rect 18658 6568 18663 6624
rect 18321 6566 18663 6568
rect 18321 6563 18387 6566
rect 18597 6563 18663 6566
rect 15006 6560 15322 6561
rect 15006 6496 15012 6560
rect 15076 6496 15092 6560
rect 15156 6496 15172 6560
rect 15236 6496 15252 6560
rect 15316 6496 15322 6560
rect 15006 6495 15322 6496
rect 5809 6488 8819 6490
rect 5809 6432 5814 6488
rect 5870 6432 8758 6488
rect 8814 6432 8819 6488
rect 5809 6430 8819 6432
rect 5809 6427 5875 6430
rect 8753 6427 8819 6430
rect 9446 6430 12450 6490
rect 16021 6492 16087 6493
rect 16021 6488 16068 6492
rect 16132 6490 16138 6492
rect 17585 6490 17651 6493
rect 18830 6490 18890 6702
rect 24166 6626 24226 6702
rect 24301 6760 25747 6762
rect 24301 6704 24306 6760
rect 24362 6704 25686 6760
rect 25742 6704 25747 6760
rect 24301 6702 25747 6704
rect 24301 6699 24367 6702
rect 25681 6699 25747 6702
rect 26233 6762 26299 6765
rect 27153 6762 27219 6765
rect 26233 6760 27219 6762
rect 26233 6704 26238 6760
rect 26294 6704 27158 6760
rect 27214 6704 27219 6760
rect 26233 6702 27219 6704
rect 26233 6699 26299 6702
rect 27153 6699 27219 6702
rect 27478 6626 27538 6838
rect 32949 6835 33015 6838
rect 38561 6898 38627 6901
rect 40880 6898 41000 6928
rect 38561 6896 41000 6898
rect 38561 6840 38566 6896
rect 38622 6840 41000 6896
rect 38561 6838 41000 6840
rect 38561 6835 38627 6838
rect 40880 6808 41000 6838
rect 29637 6762 29703 6765
rect 31109 6762 31175 6765
rect 29637 6760 31175 6762
rect 29637 6704 29642 6760
rect 29698 6704 31114 6760
rect 31170 6704 31175 6760
rect 29637 6702 31175 6704
rect 29637 6699 29703 6702
rect 31109 6699 31175 6702
rect 31661 6762 31727 6765
rect 32029 6762 32095 6765
rect 31661 6760 32095 6762
rect 31661 6704 31666 6760
rect 31722 6704 32034 6760
rect 32090 6704 32095 6760
rect 31661 6702 32095 6704
rect 31661 6699 31727 6702
rect 32029 6699 32095 6702
rect 32305 6626 32371 6629
rect 24166 6566 26848 6626
rect 27478 6624 32371 6626
rect 27478 6568 32310 6624
rect 32366 6568 32371 6624
rect 27478 6566 32371 6568
rect 21006 6560 21322 6561
rect 21006 6496 21012 6560
rect 21076 6496 21092 6560
rect 21156 6496 21172 6560
rect 21236 6496 21252 6560
rect 21316 6496 21322 6560
rect 21006 6495 21322 6496
rect 19057 6492 19123 6493
rect 16021 6432 16026 6488
rect 2681 6352 5642 6354
rect 2681 6296 2686 6352
rect 2742 6296 5642 6352
rect 2681 6294 5642 6296
rect 6821 6354 6887 6357
rect 9446 6354 9506 6430
rect 16021 6428 16068 6432
rect 16132 6430 16178 6490
rect 17585 6488 18890 6490
rect 17585 6432 17590 6488
rect 17646 6432 18890 6488
rect 17585 6430 18890 6432
rect 16132 6428 16138 6430
rect 16021 6427 16087 6428
rect 17585 6427 17651 6430
rect 19006 6428 19012 6492
rect 19076 6490 19123 6492
rect 19076 6488 19168 6490
rect 19118 6432 19168 6488
rect 19076 6430 19168 6432
rect 19076 6428 19123 6430
rect 24894 6428 24900 6492
rect 24964 6490 24970 6492
rect 25037 6490 25103 6493
rect 24964 6488 25103 6490
rect 24964 6432 25042 6488
rect 25098 6432 25103 6488
rect 24964 6430 25103 6432
rect 24964 6428 24970 6430
rect 19057 6427 19123 6428
rect 25037 6427 25103 6430
rect 26788 6357 26848 6566
rect 32305 6563 32371 6566
rect 39389 6626 39455 6629
rect 40880 6626 41000 6656
rect 39389 6624 41000 6626
rect 39389 6568 39394 6624
rect 39450 6568 41000 6624
rect 39389 6566 41000 6568
rect 39389 6563 39455 6566
rect 27006 6560 27322 6561
rect 27006 6496 27012 6560
rect 27076 6496 27092 6560
rect 27156 6496 27172 6560
rect 27236 6496 27252 6560
rect 27316 6496 27322 6560
rect 27006 6495 27322 6496
rect 33006 6560 33322 6561
rect 33006 6496 33012 6560
rect 33076 6496 33092 6560
rect 33156 6496 33172 6560
rect 33236 6496 33252 6560
rect 33316 6496 33322 6560
rect 33006 6495 33322 6496
rect 39006 6560 39322 6561
rect 39006 6496 39012 6560
rect 39076 6496 39092 6560
rect 39156 6496 39172 6560
rect 39236 6496 39252 6560
rect 39316 6496 39322 6560
rect 40880 6536 41000 6566
rect 39006 6495 39322 6496
rect 27981 6490 28047 6493
rect 31334 6490 31340 6492
rect 27981 6488 31340 6490
rect 27981 6432 27986 6488
rect 28042 6432 31340 6488
rect 27981 6430 31340 6432
rect 27981 6427 28047 6430
rect 31334 6428 31340 6430
rect 31404 6428 31410 6492
rect 6821 6352 9506 6354
rect 6821 6296 6826 6352
rect 6882 6296 9506 6352
rect 6821 6294 9506 6296
rect 9581 6354 9647 6357
rect 16481 6354 16547 6357
rect 9581 6352 16547 6354
rect 9581 6296 9586 6352
rect 9642 6296 16486 6352
rect 16542 6296 16547 6352
rect 9581 6294 16547 6296
rect 2681 6291 2747 6294
rect 6821 6291 6887 6294
rect 9581 6291 9647 6294
rect 16481 6291 16547 6294
rect 17493 6354 17559 6357
rect 18137 6354 18203 6357
rect 17493 6352 18203 6354
rect 17493 6296 17498 6352
rect 17554 6296 18142 6352
rect 18198 6296 18203 6352
rect 17493 6294 18203 6296
rect 17493 6291 17559 6294
rect 18137 6291 18203 6294
rect 18270 6292 18276 6356
rect 18340 6354 18346 6356
rect 26601 6354 26667 6357
rect 18340 6352 26667 6354
rect 18340 6296 26606 6352
rect 26662 6296 26667 6352
rect 18340 6294 26667 6296
rect 18340 6292 18346 6294
rect 26601 6291 26667 6294
rect 26785 6352 26851 6357
rect 26785 6296 26790 6352
rect 26846 6296 26851 6352
rect 26785 6291 26851 6296
rect 27613 6354 27679 6357
rect 28022 6354 28028 6356
rect 27613 6352 28028 6354
rect 27613 6296 27618 6352
rect 27674 6296 28028 6352
rect 27613 6294 28028 6296
rect 27613 6291 27679 6294
rect 28022 6292 28028 6294
rect 28092 6292 28098 6356
rect 28809 6354 28875 6357
rect 38009 6354 38075 6357
rect 28809 6352 38075 6354
rect 28809 6296 28814 6352
rect 28870 6296 38014 6352
rect 38070 6296 38075 6352
rect 28809 6294 38075 6296
rect 28809 6291 28875 6294
rect 38009 6291 38075 6294
rect 38653 6354 38719 6357
rect 40880 6354 41000 6384
rect 38653 6352 41000 6354
rect 38653 6296 38658 6352
rect 38714 6296 41000 6352
rect 38653 6294 41000 6296
rect 38653 6291 38719 6294
rect 40880 6264 41000 6294
rect 2129 6218 2195 6221
rect 12893 6218 12959 6221
rect 2129 6216 12959 6218
rect 2129 6160 2134 6216
rect 2190 6160 12898 6216
rect 12954 6160 12959 6216
rect 2129 6158 12959 6160
rect 2129 6155 2195 6158
rect 12893 6155 12959 6158
rect 13353 6218 13419 6221
rect 30649 6218 30715 6221
rect 13353 6216 30715 6218
rect 13353 6160 13358 6216
rect 13414 6160 30654 6216
rect 30710 6160 30715 6216
rect 13353 6158 30715 6160
rect 13353 6155 13419 6158
rect 30649 6155 30715 6158
rect 31753 6218 31819 6221
rect 32438 6218 32444 6220
rect 31753 6216 32444 6218
rect 31753 6160 31758 6216
rect 31814 6160 32444 6216
rect 31753 6158 32444 6160
rect 31753 6155 31819 6158
rect 32438 6156 32444 6158
rect 32508 6156 32514 6220
rect 0 6082 120 6112
rect 1209 6082 1275 6085
rect 0 6080 1275 6082
rect 0 6024 1214 6080
rect 1270 6024 1275 6080
rect 0 6022 1275 6024
rect 0 5992 120 6022
rect 1209 6019 1275 6022
rect 2497 6082 2563 6085
rect 7281 6082 7347 6085
rect 2497 6080 7347 6082
rect 2497 6024 2502 6080
rect 2558 6024 7286 6080
rect 7342 6024 7347 6080
rect 2497 6022 7347 6024
rect 2497 6019 2563 6022
rect 7281 6019 7347 6022
rect 9121 6082 9187 6085
rect 9489 6082 9555 6085
rect 11421 6082 11487 6085
rect 9121 6080 11487 6082
rect 9121 6024 9126 6080
rect 9182 6024 9494 6080
rect 9550 6024 11426 6080
rect 11482 6024 11487 6080
rect 9121 6022 11487 6024
rect 9121 6019 9187 6022
rect 9489 6019 9555 6022
rect 11421 6019 11487 6022
rect 14457 6082 14523 6085
rect 16246 6082 16252 6084
rect 14457 6080 16252 6082
rect 14457 6024 14462 6080
rect 14518 6024 16252 6080
rect 14457 6022 16252 6024
rect 14457 6019 14523 6022
rect 16246 6020 16252 6022
rect 16316 6020 16322 6084
rect 18137 6082 18203 6085
rect 18270 6082 18276 6084
rect 18137 6080 18276 6082
rect 18137 6024 18142 6080
rect 18198 6024 18276 6080
rect 18137 6022 18276 6024
rect 18137 6019 18203 6022
rect 18270 6020 18276 6022
rect 18340 6020 18346 6084
rect 18597 6082 18663 6085
rect 19241 6082 19307 6085
rect 18597 6080 19307 6082
rect 18597 6024 18602 6080
rect 18658 6024 19246 6080
rect 19302 6024 19307 6080
rect 18597 6022 19307 6024
rect 18597 6019 18663 6022
rect 19241 6019 19307 6022
rect 20345 6082 20411 6085
rect 24117 6082 24183 6085
rect 20345 6080 24183 6082
rect 20345 6024 20350 6080
rect 20406 6024 24122 6080
rect 24178 6024 24183 6080
rect 20345 6022 24183 6024
rect 20345 6019 20411 6022
rect 24117 6019 24183 6022
rect 26325 6082 26391 6085
rect 28717 6082 28783 6085
rect 26325 6080 28783 6082
rect 26325 6024 26330 6080
rect 26386 6024 28722 6080
rect 28778 6024 28783 6080
rect 26325 6022 28783 6024
rect 26325 6019 26391 6022
rect 28717 6019 28783 6022
rect 30005 6082 30071 6085
rect 31017 6082 31083 6085
rect 30005 6080 31083 6082
rect 30005 6024 30010 6080
rect 30066 6024 31022 6080
rect 31078 6024 31083 6080
rect 30005 6022 31083 6024
rect 30005 6019 30071 6022
rect 31017 6019 31083 6022
rect 38837 6082 38903 6085
rect 40880 6082 41000 6112
rect 38837 6080 41000 6082
rect 38837 6024 38842 6080
rect 38898 6024 41000 6080
rect 38837 6022 41000 6024
rect 38837 6019 38903 6022
rect 1946 6016 2262 6017
rect 1946 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2262 6016
rect 1946 5951 2262 5952
rect 7946 6016 8262 6017
rect 7946 5952 7952 6016
rect 8016 5952 8032 6016
rect 8096 5952 8112 6016
rect 8176 5952 8192 6016
rect 8256 5952 8262 6016
rect 7946 5951 8262 5952
rect 13946 6016 14262 6017
rect 13946 5952 13952 6016
rect 14016 5952 14032 6016
rect 14096 5952 14112 6016
rect 14176 5952 14192 6016
rect 14256 5952 14262 6016
rect 13946 5951 14262 5952
rect 19946 6016 20262 6017
rect 19946 5952 19952 6016
rect 20016 5952 20032 6016
rect 20096 5952 20112 6016
rect 20176 5952 20192 6016
rect 20256 5952 20262 6016
rect 19946 5951 20262 5952
rect 25946 6016 26262 6017
rect 25946 5952 25952 6016
rect 26016 5952 26032 6016
rect 26096 5952 26112 6016
rect 26176 5952 26192 6016
rect 26256 5952 26262 6016
rect 25946 5951 26262 5952
rect 31946 6016 32262 6017
rect 31946 5952 31952 6016
rect 32016 5952 32032 6016
rect 32096 5952 32112 6016
rect 32176 5952 32192 6016
rect 32256 5952 32262 6016
rect 31946 5951 32262 5952
rect 37946 6016 38262 6017
rect 37946 5952 37952 6016
rect 38016 5952 38032 6016
rect 38096 5952 38112 6016
rect 38176 5952 38192 6016
rect 38256 5952 38262 6016
rect 40880 5992 41000 6022
rect 37946 5951 38262 5952
rect 2497 5946 2563 5949
rect 2630 5946 2636 5948
rect 2497 5944 2636 5946
rect 2497 5888 2502 5944
rect 2558 5888 2636 5944
rect 2497 5886 2636 5888
rect 2497 5883 2563 5886
rect 2630 5884 2636 5886
rect 2700 5884 2706 5948
rect 3969 5946 4035 5949
rect 5574 5946 5580 5948
rect 3969 5944 5580 5946
rect 3969 5888 3974 5944
rect 4030 5888 5580 5944
rect 3969 5886 5580 5888
rect 3969 5883 4035 5886
rect 5574 5884 5580 5886
rect 5644 5884 5650 5948
rect 14590 5884 14596 5948
rect 14660 5946 14666 5948
rect 14825 5946 14891 5949
rect 19425 5946 19491 5949
rect 14660 5944 19491 5946
rect 14660 5888 14830 5944
rect 14886 5888 19430 5944
rect 19486 5888 19491 5944
rect 14660 5886 19491 5888
rect 14660 5884 14666 5886
rect 14825 5883 14891 5886
rect 19425 5883 19491 5886
rect 20621 5946 20687 5949
rect 23013 5946 23079 5949
rect 20621 5944 23079 5946
rect 20621 5888 20626 5944
rect 20682 5888 23018 5944
rect 23074 5888 23079 5944
rect 20621 5886 23079 5888
rect 20621 5883 20687 5886
rect 23013 5883 23079 5886
rect 33225 5946 33291 5949
rect 33726 5946 33732 5948
rect 33225 5944 33732 5946
rect 33225 5888 33230 5944
rect 33286 5888 33732 5944
rect 33225 5886 33732 5888
rect 33225 5883 33291 5886
rect 33726 5884 33732 5886
rect 33796 5884 33802 5948
rect 0 5810 120 5840
rect 473 5810 539 5813
rect 0 5808 539 5810
rect 0 5752 478 5808
rect 534 5752 539 5808
rect 0 5750 539 5752
rect 0 5720 120 5750
rect 473 5747 539 5750
rect 3141 5810 3207 5813
rect 4337 5810 4403 5813
rect 3141 5808 4403 5810
rect 3141 5752 3146 5808
rect 3202 5752 4342 5808
rect 4398 5752 4403 5808
rect 3141 5750 4403 5752
rect 3141 5747 3207 5750
rect 4337 5747 4403 5750
rect 5349 5810 5415 5813
rect 27337 5810 27403 5813
rect 5349 5808 27403 5810
rect 5349 5752 5354 5808
rect 5410 5752 27342 5808
rect 27398 5752 27403 5808
rect 5349 5750 27403 5752
rect 5349 5747 5415 5750
rect 27337 5747 27403 5750
rect 30833 5810 30899 5813
rect 37273 5810 37339 5813
rect 30833 5808 37339 5810
rect 30833 5752 30838 5808
rect 30894 5752 37278 5808
rect 37334 5752 37339 5808
rect 30833 5750 37339 5752
rect 30833 5747 30899 5750
rect 37273 5747 37339 5750
rect 39389 5810 39455 5813
rect 40880 5810 41000 5840
rect 39389 5808 41000 5810
rect 39389 5752 39394 5808
rect 39450 5752 41000 5808
rect 39389 5750 41000 5752
rect 39389 5747 39455 5750
rect 40880 5720 41000 5750
rect 2497 5674 2563 5677
rect 13353 5674 13419 5677
rect 2497 5672 13419 5674
rect 2497 5616 2502 5672
rect 2558 5616 13358 5672
rect 13414 5616 13419 5672
rect 2497 5614 13419 5616
rect 2497 5611 2563 5614
rect 13353 5611 13419 5614
rect 14549 5674 14615 5677
rect 15653 5674 15719 5677
rect 17125 5674 17191 5677
rect 20621 5674 20687 5677
rect 14549 5672 20687 5674
rect 14549 5616 14554 5672
rect 14610 5616 15658 5672
rect 15714 5616 17130 5672
rect 17186 5616 20626 5672
rect 20682 5616 20687 5672
rect 14549 5614 20687 5616
rect 14549 5611 14615 5614
rect 15653 5611 15719 5614
rect 17125 5611 17191 5614
rect 20621 5611 20687 5614
rect 20854 5614 21466 5674
rect 0 5538 120 5568
rect 1025 5538 1091 5541
rect 0 5536 1091 5538
rect 0 5480 1030 5536
rect 1086 5480 1091 5536
rect 0 5478 1091 5480
rect 0 5448 120 5478
rect 1025 5475 1091 5478
rect 3509 5538 3575 5541
rect 6361 5538 6427 5541
rect 8518 5538 8524 5540
rect 3509 5536 8524 5538
rect 3509 5480 3514 5536
rect 3570 5480 6366 5536
rect 6422 5480 8524 5536
rect 3509 5478 8524 5480
rect 3509 5475 3575 5478
rect 6361 5475 6427 5478
rect 8518 5476 8524 5478
rect 8588 5476 8594 5540
rect 15745 5538 15811 5541
rect 20854 5538 20914 5614
rect 15745 5536 20914 5538
rect 15745 5480 15750 5536
rect 15806 5480 20914 5536
rect 15745 5478 20914 5480
rect 21406 5538 21466 5614
rect 22134 5612 22140 5676
rect 22204 5674 22210 5676
rect 23197 5674 23263 5677
rect 22204 5672 23263 5674
rect 22204 5616 23202 5672
rect 23258 5616 23263 5672
rect 22204 5614 23263 5616
rect 22204 5612 22210 5614
rect 23197 5611 23263 5614
rect 23381 5674 23447 5677
rect 32213 5674 32279 5677
rect 23381 5672 32279 5674
rect 23381 5616 23386 5672
rect 23442 5616 32218 5672
rect 32274 5616 32279 5672
rect 23381 5614 32279 5616
rect 23381 5611 23447 5614
rect 32213 5611 32279 5614
rect 32857 5674 32923 5677
rect 37273 5674 37339 5677
rect 32857 5672 37339 5674
rect 32857 5616 32862 5672
rect 32918 5616 37278 5672
rect 37334 5616 37339 5672
rect 32857 5614 37339 5616
rect 32857 5611 32923 5614
rect 37273 5611 37339 5614
rect 37774 5612 37780 5676
rect 37844 5674 37850 5676
rect 39205 5674 39271 5677
rect 37844 5672 39271 5674
rect 37844 5616 39210 5672
rect 39266 5616 39271 5672
rect 37844 5614 39271 5616
rect 37844 5612 37850 5614
rect 39205 5611 39271 5614
rect 26601 5538 26667 5541
rect 21406 5536 26667 5538
rect 21406 5480 26606 5536
rect 26662 5480 26667 5536
rect 21406 5478 26667 5480
rect 15745 5475 15811 5478
rect 26601 5475 26667 5478
rect 39941 5538 40007 5541
rect 40880 5538 41000 5568
rect 39941 5536 41000 5538
rect 39941 5480 39946 5536
rect 40002 5480 41000 5536
rect 39941 5478 41000 5480
rect 39941 5475 40007 5478
rect 3006 5472 3322 5473
rect 3006 5408 3012 5472
rect 3076 5408 3092 5472
rect 3156 5408 3172 5472
rect 3236 5408 3252 5472
rect 3316 5408 3322 5472
rect 3006 5407 3322 5408
rect 9006 5472 9322 5473
rect 9006 5408 9012 5472
rect 9076 5408 9092 5472
rect 9156 5408 9172 5472
rect 9236 5408 9252 5472
rect 9316 5408 9322 5472
rect 9006 5407 9322 5408
rect 15006 5472 15322 5473
rect 15006 5408 15012 5472
rect 15076 5408 15092 5472
rect 15156 5408 15172 5472
rect 15236 5408 15252 5472
rect 15316 5408 15322 5472
rect 15006 5407 15322 5408
rect 21006 5472 21322 5473
rect 21006 5408 21012 5472
rect 21076 5408 21092 5472
rect 21156 5408 21172 5472
rect 21236 5408 21252 5472
rect 21316 5408 21322 5472
rect 21006 5407 21322 5408
rect 27006 5472 27322 5473
rect 27006 5408 27012 5472
rect 27076 5408 27092 5472
rect 27156 5408 27172 5472
rect 27236 5408 27252 5472
rect 27316 5408 27322 5472
rect 27006 5407 27322 5408
rect 33006 5472 33322 5473
rect 33006 5408 33012 5472
rect 33076 5408 33092 5472
rect 33156 5408 33172 5472
rect 33236 5408 33252 5472
rect 33316 5408 33322 5472
rect 33006 5407 33322 5408
rect 39006 5472 39322 5473
rect 39006 5408 39012 5472
rect 39076 5408 39092 5472
rect 39156 5408 39172 5472
rect 39236 5408 39252 5472
rect 39316 5408 39322 5472
rect 40880 5448 41000 5478
rect 39006 5407 39322 5408
rect 7005 5404 7071 5405
rect 7005 5402 7052 5404
rect 6960 5400 7052 5402
rect 6960 5344 7010 5400
rect 6960 5342 7052 5344
rect 7005 5340 7052 5342
rect 7116 5340 7122 5404
rect 8385 5402 8451 5405
rect 8702 5402 8708 5404
rect 8385 5400 8708 5402
rect 8385 5344 8390 5400
rect 8446 5344 8708 5400
rect 8385 5342 8708 5344
rect 7005 5339 7071 5340
rect 8385 5339 8451 5342
rect 8702 5340 8708 5342
rect 8772 5340 8778 5404
rect 13261 5402 13327 5405
rect 9446 5400 13327 5402
rect 9446 5344 13266 5400
rect 13322 5344 13327 5400
rect 9446 5342 13327 5344
rect 0 5266 120 5296
rect 565 5266 631 5269
rect 0 5264 631 5266
rect 0 5208 570 5264
rect 626 5208 631 5264
rect 0 5206 631 5208
rect 0 5176 120 5206
rect 565 5203 631 5206
rect 6637 5266 6703 5269
rect 9446 5266 9506 5342
rect 13261 5339 13327 5342
rect 31109 5402 31175 5405
rect 32765 5402 32831 5405
rect 31109 5400 32831 5402
rect 31109 5344 31114 5400
rect 31170 5344 32770 5400
rect 32826 5344 32831 5400
rect 31109 5342 32831 5344
rect 31109 5339 31175 5342
rect 32765 5339 32831 5342
rect 6637 5264 9506 5266
rect 6637 5208 6642 5264
rect 6698 5208 9506 5264
rect 6637 5206 9506 5208
rect 6637 5203 6703 5206
rect 9806 5204 9812 5268
rect 9876 5266 9882 5268
rect 16849 5266 16915 5269
rect 9876 5264 16915 5266
rect 9876 5208 16854 5264
rect 16910 5208 16915 5264
rect 9876 5206 16915 5208
rect 9876 5204 9882 5206
rect 16849 5203 16915 5206
rect 17309 5266 17375 5269
rect 18137 5266 18203 5269
rect 17309 5264 18203 5266
rect 17309 5208 17314 5264
rect 17370 5208 18142 5264
rect 18198 5208 18203 5264
rect 17309 5206 18203 5208
rect 17309 5203 17375 5206
rect 18137 5203 18203 5206
rect 18454 5204 18460 5268
rect 18524 5266 18530 5268
rect 18689 5266 18755 5269
rect 18524 5264 18755 5266
rect 18524 5208 18694 5264
rect 18750 5208 18755 5264
rect 18524 5206 18755 5208
rect 18524 5204 18530 5206
rect 18689 5203 18755 5206
rect 19333 5266 19399 5269
rect 35249 5266 35315 5269
rect 19333 5264 35315 5266
rect 19333 5208 19338 5264
rect 19394 5208 35254 5264
rect 35310 5208 35315 5264
rect 19333 5206 35315 5208
rect 19333 5203 19399 5206
rect 35249 5203 35315 5206
rect 39389 5266 39455 5269
rect 40880 5266 41000 5296
rect 39389 5264 41000 5266
rect 39389 5208 39394 5264
rect 39450 5208 41000 5264
rect 39389 5206 41000 5208
rect 39389 5203 39455 5206
rect 40880 5176 41000 5206
rect 1761 5130 1827 5133
rect 31569 5130 31635 5133
rect 1761 5128 31635 5130
rect 1761 5072 1766 5128
rect 1822 5072 31574 5128
rect 31630 5072 31635 5128
rect 1761 5070 31635 5072
rect 1761 5067 1827 5070
rect 31569 5067 31635 5070
rect 0 4994 120 5024
rect 1301 4994 1367 4997
rect 0 4992 1367 4994
rect 0 4936 1306 4992
rect 1362 4936 1367 4992
rect 0 4934 1367 4936
rect 0 4904 120 4934
rect 1301 4931 1367 4934
rect 8518 4932 8524 4996
rect 8588 4994 8594 4996
rect 10501 4994 10567 4997
rect 8588 4992 10567 4994
rect 8588 4936 10506 4992
rect 10562 4936 10567 4992
rect 8588 4934 10567 4936
rect 8588 4932 8594 4934
rect 10501 4931 10567 4934
rect 14825 4994 14891 4997
rect 15745 4994 15811 4997
rect 14825 4992 15811 4994
rect 14825 4936 14830 4992
rect 14886 4936 15750 4992
rect 15806 4936 15811 4992
rect 14825 4934 15811 4936
rect 14825 4931 14891 4934
rect 15745 4931 15811 4934
rect 21265 4994 21331 4997
rect 22369 4994 22435 4997
rect 21265 4992 22435 4994
rect 21265 4936 21270 4992
rect 21326 4936 22374 4992
rect 22430 4936 22435 4992
rect 21265 4934 22435 4936
rect 21265 4931 21331 4934
rect 22369 4931 22435 4934
rect 26785 4994 26851 4997
rect 27889 4994 27955 4997
rect 26785 4992 27955 4994
rect 26785 4936 26790 4992
rect 26846 4936 27894 4992
rect 27950 4936 27955 4992
rect 26785 4934 27955 4936
rect 26785 4931 26851 4934
rect 27889 4931 27955 4934
rect 39021 4994 39087 4997
rect 40880 4994 41000 5024
rect 39021 4992 41000 4994
rect 39021 4936 39026 4992
rect 39082 4936 41000 4992
rect 39021 4934 41000 4936
rect 39021 4931 39087 4934
rect 1946 4928 2262 4929
rect 1946 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2262 4928
rect 1946 4863 2262 4864
rect 7946 4928 8262 4929
rect 7946 4864 7952 4928
rect 8016 4864 8032 4928
rect 8096 4864 8112 4928
rect 8176 4864 8192 4928
rect 8256 4864 8262 4928
rect 7946 4863 8262 4864
rect 13946 4928 14262 4929
rect 13946 4864 13952 4928
rect 14016 4864 14032 4928
rect 14096 4864 14112 4928
rect 14176 4864 14192 4928
rect 14256 4864 14262 4928
rect 13946 4863 14262 4864
rect 19946 4928 20262 4929
rect 19946 4864 19952 4928
rect 20016 4864 20032 4928
rect 20096 4864 20112 4928
rect 20176 4864 20192 4928
rect 20256 4864 20262 4928
rect 19946 4863 20262 4864
rect 25946 4928 26262 4929
rect 25946 4864 25952 4928
rect 26016 4864 26032 4928
rect 26096 4864 26112 4928
rect 26176 4864 26192 4928
rect 26256 4864 26262 4928
rect 25946 4863 26262 4864
rect 31946 4928 32262 4929
rect 31946 4864 31952 4928
rect 32016 4864 32032 4928
rect 32096 4864 32112 4928
rect 32176 4864 32192 4928
rect 32256 4864 32262 4928
rect 31946 4863 32262 4864
rect 37946 4928 38262 4929
rect 37946 4864 37952 4928
rect 38016 4864 38032 4928
rect 38096 4864 38112 4928
rect 38176 4864 38192 4928
rect 38256 4864 38262 4928
rect 40880 4904 41000 4934
rect 37946 4863 38262 4864
rect 8477 4858 8543 4861
rect 9489 4858 9555 4861
rect 8477 4856 9555 4858
rect 8477 4800 8482 4856
rect 8538 4800 9494 4856
rect 9550 4800 9555 4856
rect 8477 4798 9555 4800
rect 8477 4795 8543 4798
rect 9489 4795 9555 4798
rect 10225 4858 10291 4861
rect 12617 4858 12683 4861
rect 10225 4856 12683 4858
rect 10225 4800 10230 4856
rect 10286 4800 12622 4856
rect 12678 4800 12683 4856
rect 10225 4798 12683 4800
rect 10225 4795 10291 4798
rect 12617 4795 12683 4798
rect 21173 4858 21239 4861
rect 30557 4860 30623 4861
rect 30557 4858 30604 4860
rect 21173 4856 24180 4858
rect 21173 4800 21178 4856
rect 21234 4800 24180 4856
rect 21173 4798 24180 4800
rect 30512 4856 30604 4858
rect 30512 4800 30562 4856
rect 30512 4798 30604 4800
rect 21173 4795 21239 4798
rect 0 4722 120 4752
rect 1117 4722 1183 4725
rect 0 4720 1183 4722
rect 0 4664 1122 4720
rect 1178 4664 1183 4720
rect 0 4662 1183 4664
rect 0 4632 120 4662
rect 1117 4659 1183 4662
rect 7741 4722 7807 4725
rect 23933 4722 23999 4725
rect 7741 4720 23999 4722
rect 7741 4664 7746 4720
rect 7802 4664 23938 4720
rect 23994 4664 23999 4720
rect 7741 4662 23999 4664
rect 24120 4722 24180 4798
rect 30557 4796 30604 4798
rect 30668 4796 30674 4860
rect 30557 4795 30623 4796
rect 31845 4722 31911 4725
rect 24120 4720 31911 4722
rect 24120 4664 31850 4720
rect 31906 4664 31911 4720
rect 24120 4662 31911 4664
rect 7741 4659 7807 4662
rect 23933 4659 23999 4662
rect 31845 4659 31911 4662
rect 32029 4722 32095 4725
rect 32857 4722 32923 4725
rect 32029 4720 32923 4722
rect 32029 4664 32034 4720
rect 32090 4664 32862 4720
rect 32918 4664 32923 4720
rect 32029 4662 32923 4664
rect 32029 4659 32095 4662
rect 32857 4659 32923 4662
rect 39389 4722 39455 4725
rect 40880 4722 41000 4752
rect 39389 4720 41000 4722
rect 39389 4664 39394 4720
rect 39450 4664 41000 4720
rect 39389 4662 41000 4664
rect 39389 4659 39455 4662
rect 40880 4632 41000 4662
rect 2037 4586 2103 4589
rect 35433 4586 35499 4589
rect 2037 4584 35499 4586
rect 2037 4528 2042 4584
rect 2098 4528 35438 4584
rect 35494 4528 35499 4584
rect 2037 4526 35499 4528
rect 2037 4523 2103 4526
rect 35433 4523 35499 4526
rect 0 4450 120 4480
rect 1117 4450 1183 4453
rect 0 4448 1183 4450
rect 0 4392 1122 4448
rect 1178 4392 1183 4448
rect 0 4390 1183 4392
rect 0 4360 120 4390
rect 1117 4387 1183 4390
rect 9949 4450 10015 4453
rect 11237 4450 11303 4453
rect 9949 4448 11303 4450
rect 9949 4392 9954 4448
rect 10010 4392 11242 4448
rect 11298 4392 11303 4448
rect 9949 4390 11303 4392
rect 9949 4387 10015 4390
rect 11237 4387 11303 4390
rect 11421 4450 11487 4453
rect 14733 4452 14799 4453
rect 14733 4450 14780 4452
rect 11421 4448 14780 4450
rect 14844 4450 14850 4452
rect 22461 4450 22527 4453
rect 23565 4450 23631 4453
rect 26601 4450 26667 4453
rect 11421 4392 11426 4448
rect 11482 4392 14738 4448
rect 11421 4390 14780 4392
rect 11421 4387 11487 4390
rect 14733 4388 14780 4390
rect 14844 4390 14926 4450
rect 22461 4448 26667 4450
rect 22461 4392 22466 4448
rect 22522 4392 23570 4448
rect 23626 4392 26606 4448
rect 26662 4392 26667 4448
rect 22461 4390 26667 4392
rect 14844 4388 14850 4390
rect 14733 4387 14799 4388
rect 22461 4387 22527 4390
rect 23565 4387 23631 4390
rect 26601 4387 26667 4390
rect 39849 4450 39915 4453
rect 40880 4450 41000 4480
rect 39849 4448 41000 4450
rect 39849 4392 39854 4448
rect 39910 4392 41000 4448
rect 39849 4390 41000 4392
rect 39849 4387 39915 4390
rect 3006 4384 3322 4385
rect 3006 4320 3012 4384
rect 3076 4320 3092 4384
rect 3156 4320 3172 4384
rect 3236 4320 3252 4384
rect 3316 4320 3322 4384
rect 3006 4319 3322 4320
rect 9006 4384 9322 4385
rect 9006 4320 9012 4384
rect 9076 4320 9092 4384
rect 9156 4320 9172 4384
rect 9236 4320 9252 4384
rect 9316 4320 9322 4384
rect 9006 4319 9322 4320
rect 15006 4384 15322 4385
rect 15006 4320 15012 4384
rect 15076 4320 15092 4384
rect 15156 4320 15172 4384
rect 15236 4320 15252 4384
rect 15316 4320 15322 4384
rect 15006 4319 15322 4320
rect 21006 4384 21322 4385
rect 21006 4320 21012 4384
rect 21076 4320 21092 4384
rect 21156 4320 21172 4384
rect 21236 4320 21252 4384
rect 21316 4320 21322 4384
rect 21006 4319 21322 4320
rect 27006 4384 27322 4385
rect 27006 4320 27012 4384
rect 27076 4320 27092 4384
rect 27156 4320 27172 4384
rect 27236 4320 27252 4384
rect 27316 4320 27322 4384
rect 27006 4319 27322 4320
rect 33006 4384 33322 4385
rect 33006 4320 33012 4384
rect 33076 4320 33092 4384
rect 33156 4320 33172 4384
rect 33236 4320 33252 4384
rect 33316 4320 33322 4384
rect 33006 4319 33322 4320
rect 39006 4384 39322 4385
rect 39006 4320 39012 4384
rect 39076 4320 39092 4384
rect 39156 4320 39172 4384
rect 39236 4320 39252 4384
rect 39316 4320 39322 4384
rect 40880 4360 41000 4390
rect 39006 4319 39322 4320
rect 10777 4314 10843 4317
rect 10910 4314 10916 4316
rect 5950 4254 7666 4314
rect 0 4178 120 4208
rect 381 4178 447 4181
rect 0 4176 447 4178
rect 0 4120 386 4176
rect 442 4120 447 4176
rect 0 4118 447 4120
rect 0 4088 120 4118
rect 381 4115 447 4118
rect 2773 4178 2839 4181
rect 5950 4178 6010 4254
rect 2773 4176 6010 4178
rect 2773 4120 2778 4176
rect 2834 4120 6010 4176
rect 2773 4118 6010 4120
rect 6177 4178 6243 4181
rect 7046 4178 7052 4180
rect 6177 4176 7052 4178
rect 6177 4120 6182 4176
rect 6238 4120 7052 4176
rect 6177 4118 7052 4120
rect 2773 4115 2839 4118
rect 6177 4115 6243 4118
rect 7046 4116 7052 4118
rect 7116 4116 7122 4180
rect 7606 4178 7666 4254
rect 10777 4312 10916 4314
rect 10777 4256 10782 4312
rect 10838 4256 10916 4312
rect 10777 4254 10916 4256
rect 10777 4251 10843 4254
rect 10910 4252 10916 4254
rect 10980 4252 10986 4316
rect 22369 4314 22435 4317
rect 26417 4314 26483 4317
rect 22369 4312 26483 4314
rect 22369 4256 22374 4312
rect 22430 4256 26422 4312
rect 26478 4256 26483 4312
rect 22369 4254 26483 4256
rect 22369 4251 22435 4254
rect 26417 4251 26483 4254
rect 12525 4178 12591 4181
rect 7606 4176 12591 4178
rect 7606 4120 12530 4176
rect 12586 4120 12591 4176
rect 7606 4118 12591 4120
rect 12525 4115 12591 4118
rect 15377 4178 15443 4181
rect 15653 4178 15719 4181
rect 16021 4180 16087 4181
rect 16021 4178 16068 4180
rect 15377 4176 15719 4178
rect 15377 4120 15382 4176
rect 15438 4120 15658 4176
rect 15714 4120 15719 4176
rect 15377 4118 15719 4120
rect 15976 4176 16068 4178
rect 15976 4120 16026 4176
rect 15976 4118 16068 4120
rect 15377 4115 15443 4118
rect 15653 4115 15719 4118
rect 16021 4116 16068 4118
rect 16132 4116 16138 4180
rect 17493 4178 17559 4181
rect 27981 4178 28047 4181
rect 17493 4176 28047 4178
rect 17493 4120 17498 4176
rect 17554 4120 27986 4176
rect 28042 4120 28047 4176
rect 17493 4118 28047 4120
rect 16021 4115 16087 4116
rect 17493 4115 17559 4118
rect 27981 4115 28047 4118
rect 32806 4116 32812 4180
rect 32876 4178 32882 4180
rect 32949 4178 33015 4181
rect 32876 4176 33015 4178
rect 32876 4120 32954 4176
rect 33010 4120 33015 4176
rect 32876 4118 33015 4120
rect 32876 4116 32882 4118
rect 32949 4115 33015 4118
rect 39389 4178 39455 4181
rect 40880 4178 41000 4208
rect 39389 4176 41000 4178
rect 39389 4120 39394 4176
rect 39450 4120 41000 4176
rect 39389 4118 41000 4120
rect 39389 4115 39455 4118
rect 40880 4088 41000 4118
rect 2773 4042 2839 4045
rect 25773 4042 25839 4045
rect 2773 4040 25839 4042
rect 2773 3984 2778 4040
rect 2834 3984 25778 4040
rect 25834 3984 25839 4040
rect 2773 3982 25839 3984
rect 2773 3979 2839 3982
rect 25773 3979 25839 3982
rect 26509 4042 26575 4045
rect 37273 4042 37339 4045
rect 26509 4040 37339 4042
rect 26509 3984 26514 4040
rect 26570 3984 37278 4040
rect 37334 3984 37339 4040
rect 26509 3982 37339 3984
rect 26509 3979 26575 3982
rect 37273 3979 37339 3982
rect 0 3906 120 3936
rect 749 3906 815 3909
rect 0 3904 815 3906
rect 0 3848 754 3904
rect 810 3848 815 3904
rect 0 3846 815 3848
rect 0 3816 120 3846
rect 749 3843 815 3846
rect 5349 3908 5415 3909
rect 5349 3904 5396 3908
rect 5460 3906 5466 3908
rect 8845 3906 8911 3909
rect 9397 3906 9463 3909
rect 5349 3848 5354 3904
rect 5349 3844 5396 3848
rect 5460 3846 5506 3906
rect 8845 3904 9463 3906
rect 8845 3848 8850 3904
rect 8906 3848 9402 3904
rect 9458 3848 9463 3904
rect 8845 3846 9463 3848
rect 5460 3844 5466 3846
rect 5349 3843 5415 3844
rect 8845 3843 8911 3846
rect 9397 3843 9463 3846
rect 9581 3906 9647 3909
rect 9806 3906 9812 3908
rect 9581 3904 9812 3906
rect 9581 3848 9586 3904
rect 9642 3848 9812 3904
rect 9581 3846 9812 3848
rect 9581 3843 9647 3846
rect 9806 3844 9812 3846
rect 9876 3844 9882 3908
rect 14825 3906 14891 3909
rect 15878 3906 15884 3908
rect 14825 3904 15884 3906
rect 14825 3848 14830 3904
rect 14886 3848 15884 3904
rect 14825 3846 15884 3848
rect 14825 3843 14891 3846
rect 15878 3844 15884 3846
rect 15948 3844 15954 3908
rect 26601 3906 26667 3909
rect 28901 3906 28967 3909
rect 26601 3904 28967 3906
rect 26601 3848 26606 3904
rect 26662 3848 28906 3904
rect 28962 3848 28967 3904
rect 26601 3846 28967 3848
rect 26601 3843 26667 3846
rect 28901 3843 28967 3846
rect 39021 3906 39087 3909
rect 40880 3906 41000 3936
rect 39021 3904 41000 3906
rect 39021 3848 39026 3904
rect 39082 3848 41000 3904
rect 39021 3846 41000 3848
rect 39021 3843 39087 3846
rect 1946 3840 2262 3841
rect 1946 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2262 3840
rect 1946 3775 2262 3776
rect 7946 3840 8262 3841
rect 7946 3776 7952 3840
rect 8016 3776 8032 3840
rect 8096 3776 8112 3840
rect 8176 3776 8192 3840
rect 8256 3776 8262 3840
rect 7946 3775 8262 3776
rect 13946 3840 14262 3841
rect 13946 3776 13952 3840
rect 14016 3776 14032 3840
rect 14096 3776 14112 3840
rect 14176 3776 14192 3840
rect 14256 3776 14262 3840
rect 13946 3775 14262 3776
rect 19946 3840 20262 3841
rect 19946 3776 19952 3840
rect 20016 3776 20032 3840
rect 20096 3776 20112 3840
rect 20176 3776 20192 3840
rect 20256 3776 20262 3840
rect 19946 3775 20262 3776
rect 25946 3840 26262 3841
rect 25946 3776 25952 3840
rect 26016 3776 26032 3840
rect 26096 3776 26112 3840
rect 26176 3776 26192 3840
rect 26256 3776 26262 3840
rect 25946 3775 26262 3776
rect 31946 3840 32262 3841
rect 31946 3776 31952 3840
rect 32016 3776 32032 3840
rect 32096 3776 32112 3840
rect 32176 3776 32192 3840
rect 32256 3776 32262 3840
rect 31946 3775 32262 3776
rect 37946 3840 38262 3841
rect 37946 3776 37952 3840
rect 38016 3776 38032 3840
rect 38096 3776 38112 3840
rect 38176 3776 38192 3840
rect 38256 3776 38262 3840
rect 40880 3816 41000 3846
rect 37946 3775 38262 3776
rect 7465 3770 7531 3773
rect 7598 3770 7604 3772
rect 7465 3768 7604 3770
rect 7465 3712 7470 3768
rect 7526 3712 7604 3768
rect 7465 3710 7604 3712
rect 7465 3707 7531 3710
rect 7598 3708 7604 3710
rect 7668 3708 7674 3772
rect 15510 3708 15516 3772
rect 15580 3770 15586 3772
rect 15653 3770 15719 3773
rect 15580 3768 15719 3770
rect 15580 3712 15658 3768
rect 15714 3712 15719 3768
rect 15580 3710 15719 3712
rect 15580 3708 15586 3710
rect 15653 3707 15719 3710
rect 16798 3708 16804 3772
rect 16868 3770 16874 3772
rect 18229 3770 18295 3773
rect 16868 3768 18295 3770
rect 16868 3712 18234 3768
rect 18290 3712 18295 3768
rect 16868 3710 18295 3712
rect 16868 3708 16874 3710
rect 18229 3707 18295 3710
rect 20989 3770 21055 3773
rect 24669 3770 24735 3773
rect 20989 3768 24735 3770
rect 20989 3712 20994 3768
rect 21050 3712 24674 3768
rect 24730 3712 24735 3768
rect 20989 3710 24735 3712
rect 20989 3707 21055 3710
rect 24669 3707 24735 3710
rect 26509 3770 26575 3773
rect 28165 3770 28231 3773
rect 26509 3768 28231 3770
rect 26509 3712 26514 3768
rect 26570 3712 28170 3768
rect 28226 3712 28231 3768
rect 26509 3710 28231 3712
rect 26509 3707 26575 3710
rect 28165 3707 28231 3710
rect 0 3634 120 3664
rect 749 3634 815 3637
rect 0 3632 815 3634
rect 0 3576 754 3632
rect 810 3576 815 3632
rect 0 3574 815 3576
rect 0 3544 120 3574
rect 749 3571 815 3574
rect 4337 3634 4403 3637
rect 6637 3634 6703 3637
rect 4337 3632 6703 3634
rect 4337 3576 4342 3632
rect 4398 3576 6642 3632
rect 6698 3576 6703 3632
rect 4337 3574 6703 3576
rect 4337 3571 4403 3574
rect 6637 3571 6703 3574
rect 9305 3634 9371 3637
rect 9622 3634 9628 3636
rect 9305 3632 9628 3634
rect 9305 3576 9310 3632
rect 9366 3576 9628 3632
rect 9305 3574 9628 3576
rect 9305 3571 9371 3574
rect 9622 3572 9628 3574
rect 9692 3572 9698 3636
rect 9765 3634 9831 3637
rect 26141 3634 26207 3637
rect 9765 3632 26207 3634
rect 9765 3576 9770 3632
rect 9826 3576 26146 3632
rect 26202 3576 26207 3632
rect 9765 3574 26207 3576
rect 9765 3571 9831 3574
rect 26141 3571 26207 3574
rect 26417 3634 26483 3637
rect 30189 3634 30255 3637
rect 26417 3632 30255 3634
rect 26417 3576 26422 3632
rect 26478 3576 30194 3632
rect 30250 3576 30255 3632
rect 26417 3574 30255 3576
rect 26417 3571 26483 3574
rect 30189 3571 30255 3574
rect 39389 3634 39455 3637
rect 40880 3634 41000 3664
rect 39389 3632 41000 3634
rect 39389 3576 39394 3632
rect 39450 3576 41000 3632
rect 39389 3574 41000 3576
rect 39389 3571 39455 3574
rect 40880 3544 41000 3574
rect 3049 3498 3115 3501
rect 9949 3498 10015 3501
rect 12709 3498 12775 3501
rect 3049 3496 9506 3498
rect 3049 3440 3054 3496
rect 3110 3440 9506 3496
rect 3049 3438 9506 3440
rect 3049 3435 3115 3438
rect 0 3362 120 3392
rect 2681 3362 2747 3365
rect 0 3360 2747 3362
rect 0 3304 2686 3360
rect 2742 3304 2747 3360
rect 0 3302 2747 3304
rect 0 3272 120 3302
rect 2681 3299 2747 3302
rect 7649 3362 7715 3365
rect 8477 3362 8543 3365
rect 7649 3360 8543 3362
rect 7649 3304 7654 3360
rect 7710 3304 8482 3360
rect 8538 3304 8543 3360
rect 7649 3302 8543 3304
rect 9446 3362 9506 3438
rect 9949 3496 12775 3498
rect 9949 3440 9954 3496
rect 10010 3440 12714 3496
rect 12770 3440 12775 3496
rect 9949 3438 12775 3440
rect 9949 3435 10015 3438
rect 12709 3435 12775 3438
rect 13629 3498 13695 3501
rect 13997 3498 14063 3501
rect 16205 3498 16271 3501
rect 13629 3496 14063 3498
rect 13629 3440 13634 3496
rect 13690 3440 14002 3496
rect 14058 3440 14063 3496
rect 13629 3438 14063 3440
rect 13629 3435 13695 3438
rect 13997 3435 14063 3438
rect 14828 3496 16271 3498
rect 14828 3440 16210 3496
rect 16266 3440 16271 3496
rect 14828 3438 16271 3440
rect 14828 3362 14888 3438
rect 16205 3435 16271 3438
rect 17902 3436 17908 3500
rect 17972 3498 17978 3500
rect 18689 3498 18755 3501
rect 17972 3496 18755 3498
rect 17972 3440 18694 3496
rect 18750 3440 18755 3496
rect 17972 3438 18755 3440
rect 17972 3436 17978 3438
rect 18689 3435 18755 3438
rect 18873 3498 18939 3501
rect 29913 3498 29979 3501
rect 18873 3496 29979 3498
rect 18873 3440 18878 3496
rect 18934 3440 29918 3496
rect 29974 3440 29979 3496
rect 18873 3438 29979 3440
rect 18873 3435 18939 3438
rect 29913 3435 29979 3438
rect 9446 3302 14888 3362
rect 16113 3362 16179 3365
rect 19149 3362 19215 3365
rect 16113 3360 19215 3362
rect 16113 3304 16118 3360
rect 16174 3304 19154 3360
rect 19210 3304 19215 3360
rect 16113 3302 19215 3304
rect 7649 3299 7715 3302
rect 8477 3299 8543 3302
rect 16113 3299 16179 3302
rect 19149 3299 19215 3302
rect 25313 3362 25379 3365
rect 26417 3362 26483 3365
rect 25313 3360 26483 3362
rect 25313 3304 25318 3360
rect 25374 3304 26422 3360
rect 26478 3304 26483 3360
rect 25313 3302 26483 3304
rect 25313 3299 25379 3302
rect 26417 3299 26483 3302
rect 39941 3362 40007 3365
rect 40880 3362 41000 3392
rect 39941 3360 41000 3362
rect 39941 3304 39946 3360
rect 40002 3304 41000 3360
rect 39941 3302 41000 3304
rect 39941 3299 40007 3302
rect 3006 3296 3322 3297
rect 3006 3232 3012 3296
rect 3076 3232 3092 3296
rect 3156 3232 3172 3296
rect 3236 3232 3252 3296
rect 3316 3232 3322 3296
rect 3006 3231 3322 3232
rect 9006 3296 9322 3297
rect 9006 3232 9012 3296
rect 9076 3232 9092 3296
rect 9156 3232 9172 3296
rect 9236 3232 9252 3296
rect 9316 3232 9322 3296
rect 9006 3231 9322 3232
rect 15006 3296 15322 3297
rect 15006 3232 15012 3296
rect 15076 3232 15092 3296
rect 15156 3232 15172 3296
rect 15236 3232 15252 3296
rect 15316 3232 15322 3296
rect 15006 3231 15322 3232
rect 21006 3296 21322 3297
rect 21006 3232 21012 3296
rect 21076 3232 21092 3296
rect 21156 3232 21172 3296
rect 21236 3232 21252 3296
rect 21316 3232 21322 3296
rect 21006 3231 21322 3232
rect 27006 3296 27322 3297
rect 27006 3232 27012 3296
rect 27076 3232 27092 3296
rect 27156 3232 27172 3296
rect 27236 3232 27252 3296
rect 27316 3232 27322 3296
rect 27006 3231 27322 3232
rect 33006 3296 33322 3297
rect 33006 3232 33012 3296
rect 33076 3232 33092 3296
rect 33156 3232 33172 3296
rect 33236 3232 33252 3296
rect 33316 3232 33322 3296
rect 33006 3231 33322 3232
rect 39006 3296 39322 3297
rect 39006 3232 39012 3296
rect 39076 3232 39092 3296
rect 39156 3232 39172 3296
rect 39236 3232 39252 3296
rect 39316 3232 39322 3296
rect 40880 3272 41000 3302
rect 39006 3231 39322 3232
rect 6821 3226 6887 3229
rect 8845 3226 8911 3229
rect 6821 3224 8911 3226
rect 6821 3168 6826 3224
rect 6882 3168 8850 3224
rect 8906 3168 8911 3224
rect 6821 3166 8911 3168
rect 6821 3163 6887 3166
rect 8845 3163 8911 3166
rect 9397 3226 9463 3229
rect 13169 3226 13235 3229
rect 14825 3226 14891 3229
rect 9397 3224 12450 3226
rect 9397 3168 9402 3224
rect 9458 3168 12450 3224
rect 9397 3166 12450 3168
rect 9397 3163 9463 3166
rect 0 3090 120 3120
rect 2681 3090 2747 3093
rect 0 3088 2747 3090
rect 0 3032 2686 3088
rect 2742 3032 2747 3088
rect 0 3030 2747 3032
rect 0 3000 120 3030
rect 2681 3027 2747 3030
rect 4889 3090 4955 3093
rect 12249 3090 12315 3093
rect 4889 3088 12315 3090
rect 4889 3032 4894 3088
rect 4950 3032 12254 3088
rect 12310 3032 12315 3088
rect 4889 3030 12315 3032
rect 12390 3090 12450 3166
rect 13169 3224 14891 3226
rect 13169 3168 13174 3224
rect 13230 3168 14830 3224
rect 14886 3168 14891 3224
rect 13169 3166 14891 3168
rect 13169 3163 13235 3166
rect 14825 3163 14891 3166
rect 17493 3226 17559 3229
rect 18781 3226 18847 3229
rect 24117 3228 24183 3229
rect 24117 3226 24164 3228
rect 17493 3224 18847 3226
rect 17493 3168 17498 3224
rect 17554 3168 18786 3224
rect 18842 3168 18847 3224
rect 17493 3166 18847 3168
rect 24072 3224 24164 3226
rect 24072 3168 24122 3224
rect 24072 3166 24164 3168
rect 17493 3163 17559 3166
rect 18781 3163 18847 3166
rect 24117 3164 24164 3166
rect 24228 3164 24234 3228
rect 27429 3226 27495 3229
rect 32765 3226 32831 3229
rect 27429 3224 32831 3226
rect 27429 3168 27434 3224
rect 27490 3168 32770 3224
rect 32826 3168 32831 3224
rect 27429 3166 32831 3168
rect 24117 3163 24183 3164
rect 27429 3163 27495 3166
rect 32765 3163 32831 3166
rect 12893 3090 12959 3093
rect 13997 3090 14063 3093
rect 25446 3090 25452 3092
rect 12390 3088 25452 3090
rect 12390 3032 12898 3088
rect 12954 3032 14002 3088
rect 14058 3032 25452 3088
rect 12390 3030 25452 3032
rect 4889 3027 4955 3030
rect 12249 3027 12315 3030
rect 12893 3027 12959 3030
rect 13997 3027 14063 3030
rect 25446 3028 25452 3030
rect 25516 3090 25522 3092
rect 29729 3090 29795 3093
rect 25516 3088 29795 3090
rect 25516 3032 29734 3088
rect 29790 3032 29795 3088
rect 25516 3030 29795 3032
rect 25516 3028 25522 3030
rect 29729 3027 29795 3030
rect 32121 3090 32187 3093
rect 33409 3090 33475 3093
rect 32121 3088 33475 3090
rect 32121 3032 32126 3088
rect 32182 3032 33414 3088
rect 33470 3032 33475 3088
rect 32121 3030 33475 3032
rect 32121 3027 32187 3030
rect 33409 3027 33475 3030
rect 39389 3090 39455 3093
rect 40880 3090 41000 3120
rect 39389 3088 41000 3090
rect 39389 3032 39394 3088
rect 39450 3032 41000 3088
rect 39389 3030 41000 3032
rect 39389 3027 39455 3030
rect 40880 3000 41000 3030
rect 4061 2954 4127 2957
rect 18689 2954 18755 2957
rect 19425 2954 19491 2957
rect 21909 2954 21975 2957
rect 4061 2952 19491 2954
rect 4061 2896 4066 2952
rect 4122 2896 18694 2952
rect 18750 2896 19430 2952
rect 19486 2896 19491 2952
rect 4061 2894 19491 2896
rect 4061 2891 4127 2894
rect 18689 2891 18755 2894
rect 19425 2891 19491 2894
rect 19796 2952 21975 2954
rect 19796 2896 21914 2952
rect 21970 2896 21975 2952
rect 19796 2894 21975 2896
rect 0 2818 120 2848
rect 565 2818 631 2821
rect 0 2816 631 2818
rect 0 2760 570 2816
rect 626 2760 631 2816
rect 0 2758 631 2760
rect 0 2728 120 2758
rect 565 2755 631 2758
rect 10593 2818 10659 2821
rect 10869 2818 10935 2821
rect 10593 2816 10935 2818
rect 10593 2760 10598 2816
rect 10654 2760 10874 2816
rect 10930 2760 10935 2816
rect 10593 2758 10935 2760
rect 10593 2755 10659 2758
rect 10869 2755 10935 2758
rect 11053 2818 11119 2821
rect 13537 2818 13603 2821
rect 11053 2816 13603 2818
rect 11053 2760 11058 2816
rect 11114 2760 13542 2816
rect 13598 2760 13603 2816
rect 11053 2758 13603 2760
rect 11053 2755 11119 2758
rect 13537 2755 13603 2758
rect 14365 2818 14431 2821
rect 19796 2818 19856 2894
rect 21909 2891 21975 2894
rect 25957 2954 26023 2957
rect 26601 2956 26667 2957
rect 26366 2954 26372 2956
rect 25957 2952 26372 2954
rect 25957 2896 25962 2952
rect 26018 2896 26372 2952
rect 25957 2894 26372 2896
rect 25957 2891 26023 2894
rect 26366 2892 26372 2894
rect 26436 2892 26442 2956
rect 26550 2892 26556 2956
rect 26620 2954 26667 2956
rect 27613 2954 27679 2957
rect 36629 2954 36695 2957
rect 26620 2952 26712 2954
rect 26662 2896 26712 2952
rect 26620 2894 26712 2896
rect 27613 2952 36695 2954
rect 27613 2896 27618 2952
rect 27674 2896 36634 2952
rect 36690 2896 36695 2952
rect 27613 2894 36695 2896
rect 26620 2892 26667 2894
rect 26601 2891 26667 2892
rect 27613 2891 27679 2894
rect 36629 2891 36695 2894
rect 14365 2816 19856 2818
rect 14365 2760 14370 2816
rect 14426 2760 19856 2816
rect 14365 2758 19856 2760
rect 20345 2818 20411 2821
rect 25773 2818 25839 2821
rect 20345 2816 25839 2818
rect 20345 2760 20350 2816
rect 20406 2760 25778 2816
rect 25834 2760 25839 2816
rect 20345 2758 25839 2760
rect 14365 2755 14431 2758
rect 20345 2755 20411 2758
rect 25773 2755 25839 2758
rect 27245 2818 27311 2821
rect 27521 2818 27587 2821
rect 27245 2816 27587 2818
rect 27245 2760 27250 2816
rect 27306 2760 27526 2816
rect 27582 2760 27587 2816
rect 27245 2758 27587 2760
rect 27245 2755 27311 2758
rect 27521 2755 27587 2758
rect 32581 2818 32647 2821
rect 32949 2818 33015 2821
rect 32581 2816 33015 2818
rect 32581 2760 32586 2816
rect 32642 2760 32954 2816
rect 33010 2760 33015 2816
rect 32581 2758 33015 2760
rect 32581 2755 32647 2758
rect 32949 2755 33015 2758
rect 39021 2818 39087 2821
rect 40880 2818 41000 2848
rect 39021 2816 41000 2818
rect 39021 2760 39026 2816
rect 39082 2760 41000 2816
rect 39021 2758 41000 2760
rect 39021 2755 39087 2758
rect 1946 2752 2262 2753
rect 1946 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2262 2752
rect 1946 2687 2262 2688
rect 7946 2752 8262 2753
rect 7946 2688 7952 2752
rect 8016 2688 8032 2752
rect 8096 2688 8112 2752
rect 8176 2688 8192 2752
rect 8256 2688 8262 2752
rect 7946 2687 8262 2688
rect 13946 2752 14262 2753
rect 13946 2688 13952 2752
rect 14016 2688 14032 2752
rect 14096 2688 14112 2752
rect 14176 2688 14192 2752
rect 14256 2688 14262 2752
rect 13946 2687 14262 2688
rect 19946 2752 20262 2753
rect 19946 2688 19952 2752
rect 20016 2688 20032 2752
rect 20096 2688 20112 2752
rect 20176 2688 20192 2752
rect 20256 2688 20262 2752
rect 19946 2687 20262 2688
rect 25946 2752 26262 2753
rect 25946 2688 25952 2752
rect 26016 2688 26032 2752
rect 26096 2688 26112 2752
rect 26176 2688 26192 2752
rect 26256 2688 26262 2752
rect 25946 2687 26262 2688
rect 31946 2752 32262 2753
rect 31946 2688 31952 2752
rect 32016 2688 32032 2752
rect 32096 2688 32112 2752
rect 32176 2688 32192 2752
rect 32256 2688 32262 2752
rect 31946 2687 32262 2688
rect 37946 2752 38262 2753
rect 37946 2688 37952 2752
rect 38016 2688 38032 2752
rect 38096 2688 38112 2752
rect 38176 2688 38192 2752
rect 38256 2688 38262 2752
rect 40880 2728 41000 2758
rect 37946 2687 38262 2688
rect 8661 2682 8727 2685
rect 11145 2682 11211 2685
rect 12157 2682 12223 2685
rect 18505 2682 18571 2685
rect 8661 2680 11211 2682
rect 8661 2624 8666 2680
rect 8722 2624 11150 2680
rect 11206 2624 11211 2680
rect 8661 2622 11211 2624
rect 8661 2619 8727 2622
rect 11145 2619 11211 2622
rect 11286 2680 12223 2682
rect 11286 2624 12162 2680
rect 12218 2624 12223 2680
rect 11286 2622 12223 2624
rect 0 2546 120 2576
rect 2589 2546 2655 2549
rect 0 2544 2655 2546
rect 0 2488 2594 2544
rect 2650 2488 2655 2544
rect 0 2486 2655 2488
rect 0 2456 120 2486
rect 2589 2483 2655 2486
rect 4889 2546 4955 2549
rect 11286 2546 11346 2622
rect 12157 2619 12223 2622
rect 14414 2680 18571 2682
rect 14414 2624 18510 2680
rect 18566 2624 18571 2680
rect 14414 2622 18571 2624
rect 4889 2544 11346 2546
rect 4889 2488 4894 2544
rect 4950 2488 11346 2544
rect 4889 2486 11346 2488
rect 11881 2546 11947 2549
rect 14414 2546 14474 2622
rect 18505 2619 18571 2622
rect 11881 2544 14474 2546
rect 11881 2488 11886 2544
rect 11942 2488 14474 2544
rect 11881 2486 14474 2488
rect 14549 2548 14615 2549
rect 14549 2544 14596 2548
rect 14660 2546 14666 2548
rect 16481 2546 16547 2549
rect 37774 2546 37780 2548
rect 14549 2488 14554 2544
rect 4889 2483 4955 2486
rect 11881 2483 11947 2486
rect 14549 2484 14596 2488
rect 14660 2486 14706 2546
rect 16481 2544 37780 2546
rect 16481 2488 16486 2544
rect 16542 2488 37780 2544
rect 16481 2486 37780 2488
rect 14660 2484 14666 2486
rect 14549 2483 14615 2484
rect 16481 2483 16547 2486
rect 37774 2484 37780 2486
rect 37844 2484 37850 2548
rect 39389 2546 39455 2549
rect 40880 2546 41000 2576
rect 39389 2544 41000 2546
rect 39389 2488 39394 2544
rect 39450 2488 41000 2544
rect 39389 2486 41000 2488
rect 39389 2483 39455 2486
rect 40880 2456 41000 2486
rect 1669 2410 1735 2413
rect 19241 2410 19307 2413
rect 1669 2408 19307 2410
rect 1669 2352 1674 2408
rect 1730 2352 19246 2408
rect 19302 2352 19307 2408
rect 1669 2350 19307 2352
rect 1669 2347 1735 2350
rect 19241 2347 19307 2350
rect 21081 2410 21147 2413
rect 23565 2410 23631 2413
rect 28625 2410 28691 2413
rect 21081 2408 28691 2410
rect 21081 2352 21086 2408
rect 21142 2352 23570 2408
rect 23626 2352 28630 2408
rect 28686 2352 28691 2408
rect 21081 2350 28691 2352
rect 21081 2347 21147 2350
rect 23565 2347 23631 2350
rect 28625 2347 28691 2350
rect 0 2274 120 2304
rect 1301 2274 1367 2277
rect 10317 2276 10383 2277
rect 10317 2274 10364 2276
rect 0 2272 1367 2274
rect 0 2216 1306 2272
rect 1362 2216 1367 2272
rect 0 2214 1367 2216
rect 10276 2272 10364 2274
rect 10428 2274 10434 2276
rect 14273 2274 14339 2277
rect 10428 2272 14339 2274
rect 10276 2216 10322 2272
rect 10428 2216 14278 2272
rect 14334 2216 14339 2272
rect 10276 2214 10364 2216
rect 0 2184 120 2214
rect 1301 2211 1367 2214
rect 10317 2212 10364 2214
rect 10428 2214 14339 2216
rect 10428 2212 10434 2214
rect 10317 2211 10383 2212
rect 14273 2211 14339 2214
rect 39941 2274 40007 2277
rect 40880 2274 41000 2304
rect 39941 2272 41000 2274
rect 39941 2216 39946 2272
rect 40002 2216 41000 2272
rect 39941 2214 41000 2216
rect 39941 2211 40007 2214
rect 3006 2208 3322 2209
rect 3006 2144 3012 2208
rect 3076 2144 3092 2208
rect 3156 2144 3172 2208
rect 3236 2144 3252 2208
rect 3316 2144 3322 2208
rect 3006 2143 3322 2144
rect 9006 2208 9322 2209
rect 9006 2144 9012 2208
rect 9076 2144 9092 2208
rect 9156 2144 9172 2208
rect 9236 2144 9252 2208
rect 9316 2144 9322 2208
rect 9006 2143 9322 2144
rect 15006 2208 15322 2209
rect 15006 2144 15012 2208
rect 15076 2144 15092 2208
rect 15156 2144 15172 2208
rect 15236 2144 15252 2208
rect 15316 2144 15322 2208
rect 15006 2143 15322 2144
rect 21006 2208 21322 2209
rect 21006 2144 21012 2208
rect 21076 2144 21092 2208
rect 21156 2144 21172 2208
rect 21236 2144 21252 2208
rect 21316 2144 21322 2208
rect 21006 2143 21322 2144
rect 27006 2208 27322 2209
rect 27006 2144 27012 2208
rect 27076 2144 27092 2208
rect 27156 2144 27172 2208
rect 27236 2144 27252 2208
rect 27316 2144 27322 2208
rect 27006 2143 27322 2144
rect 33006 2208 33322 2209
rect 33006 2144 33012 2208
rect 33076 2144 33092 2208
rect 33156 2144 33172 2208
rect 33236 2144 33252 2208
rect 33316 2144 33322 2208
rect 33006 2143 33322 2144
rect 39006 2208 39322 2209
rect 39006 2144 39012 2208
rect 39076 2144 39092 2208
rect 39156 2144 39172 2208
rect 39236 2144 39252 2208
rect 39316 2144 39322 2208
rect 40880 2184 41000 2214
rect 39006 2143 39322 2144
rect 10501 2138 10567 2141
rect 14641 2138 14707 2141
rect 10501 2136 14707 2138
rect 10501 2080 10506 2136
rect 10562 2080 14646 2136
rect 14702 2080 14707 2136
rect 10501 2078 14707 2080
rect 10501 2075 10567 2078
rect 14641 2075 14707 2078
rect 0 2002 120 2032
rect 2313 2002 2379 2005
rect 0 2000 2379 2002
rect 0 1944 2318 2000
rect 2374 1944 2379 2000
rect 0 1942 2379 1944
rect 0 1912 120 1942
rect 2313 1939 2379 1942
rect 7097 2002 7163 2005
rect 19333 2002 19399 2005
rect 7097 2000 19399 2002
rect 7097 1944 7102 2000
rect 7158 1944 19338 2000
rect 19394 1944 19399 2000
rect 7097 1942 19399 1944
rect 7097 1939 7163 1942
rect 19333 1939 19399 1942
rect 26509 2002 26575 2005
rect 37089 2002 37155 2005
rect 26509 2000 37155 2002
rect 26509 1944 26514 2000
rect 26570 1944 37094 2000
rect 37150 1944 37155 2000
rect 26509 1942 37155 1944
rect 26509 1939 26575 1942
rect 37089 1939 37155 1942
rect 38929 2002 38995 2005
rect 40880 2002 41000 2032
rect 38929 2000 41000 2002
rect 38929 1944 38934 2000
rect 38990 1944 41000 2000
rect 38929 1942 41000 1944
rect 38929 1939 38995 1942
rect 40880 1912 41000 1942
rect 4061 1866 4127 1869
rect 19793 1866 19859 1869
rect 38745 1866 38811 1869
rect 4061 1864 19859 1866
rect 4061 1808 4066 1864
rect 4122 1808 19798 1864
rect 19854 1808 19859 1864
rect 4061 1806 19859 1808
rect 4061 1803 4127 1806
rect 19793 1803 19859 1806
rect 22050 1864 38811 1866
rect 22050 1808 38750 1864
rect 38806 1808 38811 1864
rect 22050 1806 38811 1808
rect 0 1730 120 1760
rect 381 1730 447 1733
rect 0 1728 447 1730
rect 0 1672 386 1728
rect 442 1672 447 1728
rect 0 1670 447 1672
rect 0 1640 120 1670
rect 381 1667 447 1670
rect 7046 1668 7052 1732
rect 7116 1730 7122 1732
rect 17861 1730 17927 1733
rect 22050 1730 22110 1806
rect 38745 1803 38811 1806
rect 7116 1670 16590 1730
rect 7116 1668 7122 1670
rect 9581 1594 9647 1597
rect 11145 1594 11211 1597
rect 9581 1592 11211 1594
rect 9581 1536 9586 1592
rect 9642 1536 11150 1592
rect 11206 1536 11211 1592
rect 9581 1534 11211 1536
rect 16530 1594 16590 1670
rect 17861 1728 22110 1730
rect 17861 1672 17866 1728
rect 17922 1672 22110 1728
rect 17861 1670 22110 1672
rect 37917 1730 37983 1733
rect 40880 1730 41000 1760
rect 37917 1728 41000 1730
rect 37917 1672 37922 1728
rect 37978 1672 41000 1728
rect 37917 1670 41000 1672
rect 17861 1667 17927 1670
rect 37917 1667 37983 1670
rect 40880 1640 41000 1670
rect 27337 1594 27403 1597
rect 16530 1592 27403 1594
rect 16530 1536 27342 1592
rect 27398 1536 27403 1592
rect 16530 1534 27403 1536
rect 9581 1531 9647 1534
rect 11145 1531 11211 1534
rect 27337 1531 27403 1534
rect 0 1458 120 1488
rect 933 1458 999 1461
rect 0 1456 999 1458
rect 0 1400 938 1456
rect 994 1400 999 1456
rect 0 1398 999 1400
rect 0 1368 120 1398
rect 933 1395 999 1398
rect 3918 1396 3924 1460
rect 3988 1458 3994 1460
rect 17493 1458 17559 1461
rect 3988 1456 17559 1458
rect 3988 1400 17498 1456
rect 17554 1400 17559 1456
rect 3988 1398 17559 1400
rect 3988 1396 3994 1398
rect 17493 1395 17559 1398
rect 38285 1458 38351 1461
rect 40880 1458 41000 1488
rect 38285 1456 41000 1458
rect 38285 1400 38290 1456
rect 38346 1400 41000 1456
rect 38285 1398 41000 1400
rect 38285 1395 38351 1398
rect 40880 1368 41000 1398
rect 4613 1322 4679 1325
rect 39849 1322 39915 1325
rect 4613 1320 39915 1322
rect 4613 1264 4618 1320
rect 4674 1264 39854 1320
rect 39910 1264 39915 1320
rect 4613 1262 39915 1264
rect 4613 1259 4679 1262
rect 39849 1259 39915 1262
rect 5574 1124 5580 1188
rect 5644 1186 5650 1188
rect 39665 1186 39731 1189
rect 5644 1184 39731 1186
rect 5644 1128 39670 1184
rect 39726 1128 39731 1184
rect 5644 1126 39731 1128
rect 5644 1124 5650 1126
rect 39665 1123 39731 1126
rect 2446 988 2452 1052
rect 2516 1050 2522 1052
rect 33501 1050 33567 1053
rect 2516 1048 33567 1050
rect 2516 992 33506 1048
rect 33562 992 33567 1048
rect 2516 990 33567 992
rect 2516 988 2522 990
rect 33501 987 33567 990
rect 6678 852 6684 916
rect 6748 914 6754 916
rect 35801 914 35867 917
rect 6748 912 35867 914
rect 6748 856 35806 912
rect 35862 856 35867 912
rect 6748 854 35867 856
rect 6748 852 6754 854
rect 35801 851 35867 854
rect 3969 778 4035 781
rect 27705 778 27771 781
rect 3969 776 27771 778
rect 3969 720 3974 776
rect 4030 720 27710 776
rect 27766 720 27771 776
rect 3969 718 27771 720
rect 3969 715 4035 718
rect 27705 715 27771 718
rect 29821 778 29887 781
rect 35709 778 35775 781
rect 29821 776 35775 778
rect 29821 720 29826 776
rect 29882 720 35714 776
rect 35770 720 35775 776
rect 29821 718 35775 720
rect 29821 715 29887 718
rect 35709 715 35775 718
rect 2589 642 2655 645
rect 25262 642 25268 644
rect 2589 640 25268 642
rect 2589 584 2594 640
rect 2650 584 25268 640
rect 2589 582 25268 584
rect 2589 579 2655 582
rect 25262 580 25268 582
rect 25332 580 25338 644
rect 5625 506 5691 509
rect 22134 506 22140 508
rect 5625 504 22140 506
rect 5625 448 5630 504
rect 5686 448 22140 504
rect 5625 446 22140 448
rect 5625 443 5691 446
rect 22134 444 22140 446
rect 22204 444 22210 508
<< via3 >>
rect 2636 10100 2700 10164
rect 26740 10372 26804 10436
rect 24900 10236 24964 10300
rect 7788 9964 7852 10028
rect 23428 9964 23492 10028
rect 33732 9888 33796 9892
rect 33732 9832 33782 9888
rect 33782 9832 33796 9888
rect 33732 9828 33796 9832
rect 15516 9420 15580 9484
rect 32444 9420 32508 9484
rect 7604 9284 7668 9348
rect 24164 9148 24228 9212
rect 32812 9012 32876 9076
rect 3012 8732 3076 8736
rect 3012 8676 3016 8732
rect 3016 8676 3072 8732
rect 3072 8676 3076 8732
rect 3012 8672 3076 8676
rect 3092 8732 3156 8736
rect 3092 8676 3096 8732
rect 3096 8676 3152 8732
rect 3152 8676 3156 8732
rect 3092 8672 3156 8676
rect 3172 8732 3236 8736
rect 3172 8676 3176 8732
rect 3176 8676 3232 8732
rect 3232 8676 3236 8732
rect 3172 8672 3236 8676
rect 3252 8732 3316 8736
rect 3252 8676 3256 8732
rect 3256 8676 3312 8732
rect 3312 8676 3316 8732
rect 3252 8672 3316 8676
rect 9628 8740 9692 8804
rect 9012 8732 9076 8736
rect 9012 8676 9016 8732
rect 9016 8676 9072 8732
rect 9072 8676 9076 8732
rect 9012 8672 9076 8676
rect 9092 8732 9156 8736
rect 9092 8676 9096 8732
rect 9096 8676 9152 8732
rect 9152 8676 9156 8732
rect 9092 8672 9156 8676
rect 9172 8732 9236 8736
rect 9172 8676 9176 8732
rect 9176 8676 9232 8732
rect 9232 8676 9236 8732
rect 9172 8672 9236 8676
rect 9252 8732 9316 8736
rect 9252 8676 9256 8732
rect 9256 8676 9312 8732
rect 9312 8676 9316 8732
rect 9252 8672 9316 8676
rect 7052 8468 7116 8532
rect 15012 8732 15076 8736
rect 15012 8676 15016 8732
rect 15016 8676 15072 8732
rect 15072 8676 15076 8732
rect 15012 8672 15076 8676
rect 15092 8732 15156 8736
rect 15092 8676 15096 8732
rect 15096 8676 15152 8732
rect 15152 8676 15156 8732
rect 15092 8672 15156 8676
rect 15172 8732 15236 8736
rect 15172 8676 15176 8732
rect 15176 8676 15232 8732
rect 15232 8676 15236 8732
rect 15172 8672 15236 8676
rect 15252 8732 15316 8736
rect 15252 8676 15256 8732
rect 15256 8676 15312 8732
rect 15312 8676 15316 8732
rect 15252 8672 15316 8676
rect 21012 8732 21076 8736
rect 21012 8676 21016 8732
rect 21016 8676 21072 8732
rect 21072 8676 21076 8732
rect 21012 8672 21076 8676
rect 21092 8732 21156 8736
rect 21092 8676 21096 8732
rect 21096 8676 21152 8732
rect 21152 8676 21156 8732
rect 21092 8672 21156 8676
rect 21172 8732 21236 8736
rect 21172 8676 21176 8732
rect 21176 8676 21232 8732
rect 21232 8676 21236 8732
rect 21172 8672 21236 8676
rect 21252 8732 21316 8736
rect 21252 8676 21256 8732
rect 21256 8676 21312 8732
rect 21312 8676 21316 8732
rect 21252 8672 21316 8676
rect 27012 8732 27076 8736
rect 27012 8676 27016 8732
rect 27016 8676 27072 8732
rect 27072 8676 27076 8732
rect 27012 8672 27076 8676
rect 27092 8732 27156 8736
rect 27092 8676 27096 8732
rect 27096 8676 27152 8732
rect 27152 8676 27156 8732
rect 27092 8672 27156 8676
rect 27172 8732 27236 8736
rect 27172 8676 27176 8732
rect 27176 8676 27232 8732
rect 27232 8676 27236 8732
rect 27172 8672 27236 8676
rect 27252 8732 27316 8736
rect 27252 8676 27256 8732
rect 27256 8676 27312 8732
rect 27312 8676 27316 8732
rect 27252 8672 27316 8676
rect 33012 8732 33076 8736
rect 33012 8676 33016 8732
rect 33016 8676 33072 8732
rect 33072 8676 33076 8732
rect 33012 8672 33076 8676
rect 33092 8732 33156 8736
rect 33092 8676 33096 8732
rect 33096 8676 33152 8732
rect 33152 8676 33156 8732
rect 33092 8672 33156 8676
rect 33172 8732 33236 8736
rect 33172 8676 33176 8732
rect 33176 8676 33232 8732
rect 33232 8676 33236 8732
rect 33172 8672 33236 8676
rect 33252 8732 33316 8736
rect 33252 8676 33256 8732
rect 33256 8676 33312 8732
rect 33312 8676 33316 8732
rect 33252 8672 33316 8676
rect 39012 8732 39076 8736
rect 39012 8676 39016 8732
rect 39016 8676 39072 8732
rect 39072 8676 39076 8732
rect 39012 8672 39076 8676
rect 39092 8732 39156 8736
rect 39092 8676 39096 8732
rect 39096 8676 39152 8732
rect 39152 8676 39156 8732
rect 39092 8672 39156 8676
rect 39172 8732 39236 8736
rect 39172 8676 39176 8732
rect 39176 8676 39232 8732
rect 39232 8676 39236 8732
rect 39172 8672 39236 8676
rect 39252 8732 39316 8736
rect 39252 8676 39256 8732
rect 39256 8676 39312 8732
rect 39312 8676 39316 8732
rect 39252 8672 39316 8676
rect 18644 8664 18708 8668
rect 18644 8608 18694 8664
rect 18694 8608 18708 8664
rect 18644 8604 18708 8608
rect 28028 8664 28092 8668
rect 28028 8608 28078 8664
rect 28078 8608 28092 8664
rect 16804 8468 16868 8532
rect 28028 8604 28092 8608
rect 25268 8528 25332 8532
rect 25268 8472 25282 8528
rect 25282 8472 25332 8528
rect 25268 8468 25332 8472
rect 26556 8468 26620 8532
rect 17908 8332 17972 8396
rect 7788 8256 7852 8260
rect 7788 8200 7802 8256
rect 7802 8200 7852 8256
rect 7788 8196 7852 8200
rect 8524 8196 8588 8260
rect 25452 8196 25516 8260
rect 1952 8188 2016 8192
rect 1952 8132 1956 8188
rect 1956 8132 2012 8188
rect 2012 8132 2016 8188
rect 1952 8128 2016 8132
rect 2032 8188 2096 8192
rect 2032 8132 2036 8188
rect 2036 8132 2092 8188
rect 2092 8132 2096 8188
rect 2032 8128 2096 8132
rect 2112 8188 2176 8192
rect 2112 8132 2116 8188
rect 2116 8132 2172 8188
rect 2172 8132 2176 8188
rect 2112 8128 2176 8132
rect 2192 8188 2256 8192
rect 2192 8132 2196 8188
rect 2196 8132 2252 8188
rect 2252 8132 2256 8188
rect 2192 8128 2256 8132
rect 7952 8188 8016 8192
rect 7952 8132 7956 8188
rect 7956 8132 8012 8188
rect 8012 8132 8016 8188
rect 7952 8128 8016 8132
rect 8032 8188 8096 8192
rect 8032 8132 8036 8188
rect 8036 8132 8092 8188
rect 8092 8132 8096 8188
rect 8032 8128 8096 8132
rect 8112 8188 8176 8192
rect 8112 8132 8116 8188
rect 8116 8132 8172 8188
rect 8172 8132 8176 8188
rect 8112 8128 8176 8132
rect 8192 8188 8256 8192
rect 8192 8132 8196 8188
rect 8196 8132 8252 8188
rect 8252 8132 8256 8188
rect 8192 8128 8256 8132
rect 13952 8188 14016 8192
rect 13952 8132 13956 8188
rect 13956 8132 14012 8188
rect 14012 8132 14016 8188
rect 13952 8128 14016 8132
rect 14032 8188 14096 8192
rect 14032 8132 14036 8188
rect 14036 8132 14092 8188
rect 14092 8132 14096 8188
rect 14032 8128 14096 8132
rect 14112 8188 14176 8192
rect 14112 8132 14116 8188
rect 14116 8132 14172 8188
rect 14172 8132 14176 8188
rect 14112 8128 14176 8132
rect 14192 8188 14256 8192
rect 14192 8132 14196 8188
rect 14196 8132 14252 8188
rect 14252 8132 14256 8188
rect 14192 8128 14256 8132
rect 19952 8188 20016 8192
rect 19952 8132 19956 8188
rect 19956 8132 20012 8188
rect 20012 8132 20016 8188
rect 19952 8128 20016 8132
rect 20032 8188 20096 8192
rect 20032 8132 20036 8188
rect 20036 8132 20092 8188
rect 20092 8132 20096 8188
rect 20032 8128 20096 8132
rect 20112 8188 20176 8192
rect 20112 8132 20116 8188
rect 20116 8132 20172 8188
rect 20172 8132 20176 8188
rect 20112 8128 20176 8132
rect 20192 8188 20256 8192
rect 20192 8132 20196 8188
rect 20196 8132 20252 8188
rect 20252 8132 20256 8188
rect 20192 8128 20256 8132
rect 25952 8188 26016 8192
rect 25952 8132 25956 8188
rect 25956 8132 26012 8188
rect 26012 8132 26016 8188
rect 25952 8128 26016 8132
rect 26032 8188 26096 8192
rect 26032 8132 26036 8188
rect 26036 8132 26092 8188
rect 26092 8132 26096 8188
rect 26032 8128 26096 8132
rect 26112 8188 26176 8192
rect 26112 8132 26116 8188
rect 26116 8132 26172 8188
rect 26172 8132 26176 8188
rect 26112 8128 26176 8132
rect 26192 8188 26256 8192
rect 26192 8132 26196 8188
rect 26196 8132 26252 8188
rect 26252 8132 26256 8188
rect 26192 8128 26256 8132
rect 18460 8060 18524 8124
rect 19012 8120 19076 8124
rect 19012 8064 19062 8120
rect 19062 8064 19076 8120
rect 19012 8060 19076 8064
rect 25636 8060 25700 8124
rect 26372 8060 26436 8124
rect 31952 8188 32016 8192
rect 31952 8132 31956 8188
rect 31956 8132 32012 8188
rect 32012 8132 32016 8188
rect 31952 8128 32016 8132
rect 32032 8188 32096 8192
rect 32032 8132 32036 8188
rect 32036 8132 32092 8188
rect 32092 8132 32096 8188
rect 32032 8128 32096 8132
rect 32112 8188 32176 8192
rect 32112 8132 32116 8188
rect 32116 8132 32172 8188
rect 32172 8132 32176 8188
rect 32112 8128 32176 8132
rect 32192 8188 32256 8192
rect 32192 8132 32196 8188
rect 32196 8132 32252 8188
rect 32252 8132 32256 8188
rect 32192 8128 32256 8132
rect 37952 8188 38016 8192
rect 37952 8132 37956 8188
rect 37956 8132 38012 8188
rect 38012 8132 38016 8188
rect 37952 8128 38016 8132
rect 38032 8188 38096 8192
rect 38032 8132 38036 8188
rect 38036 8132 38092 8188
rect 38092 8132 38096 8188
rect 38032 8128 38096 8132
rect 38112 8188 38176 8192
rect 38112 8132 38116 8188
rect 38116 8132 38172 8188
rect 38172 8132 38176 8188
rect 38112 8128 38176 8132
rect 38192 8188 38256 8192
rect 38192 8132 38196 8188
rect 38196 8132 38252 8188
rect 38252 8132 38256 8188
rect 38192 8128 38256 8132
rect 30604 8060 30668 8124
rect 32628 8060 32692 8124
rect 3012 7644 3076 7648
rect 3012 7588 3016 7644
rect 3016 7588 3072 7644
rect 3072 7588 3076 7644
rect 3012 7584 3076 7588
rect 3092 7644 3156 7648
rect 3092 7588 3096 7644
rect 3096 7588 3152 7644
rect 3152 7588 3156 7644
rect 3092 7584 3156 7588
rect 3172 7644 3236 7648
rect 3172 7588 3176 7644
rect 3176 7588 3232 7644
rect 3232 7588 3236 7644
rect 3172 7584 3236 7588
rect 3252 7644 3316 7648
rect 3252 7588 3256 7644
rect 3256 7588 3312 7644
rect 3312 7588 3316 7644
rect 3252 7584 3316 7588
rect 10916 7788 10980 7852
rect 9012 7644 9076 7648
rect 9012 7588 9016 7644
rect 9016 7588 9072 7644
rect 9072 7588 9076 7644
rect 9012 7584 9076 7588
rect 9092 7644 9156 7648
rect 9092 7588 9096 7644
rect 9096 7588 9152 7644
rect 9152 7588 9156 7644
rect 9092 7584 9156 7588
rect 9172 7644 9236 7648
rect 9172 7588 9176 7644
rect 9176 7588 9232 7644
rect 9232 7588 9236 7644
rect 9172 7584 9236 7588
rect 9252 7644 9316 7648
rect 9252 7588 9256 7644
rect 9256 7588 9312 7644
rect 9312 7588 9316 7644
rect 9252 7584 9316 7588
rect 10364 7576 10428 7580
rect 10364 7520 10378 7576
rect 10378 7520 10428 7576
rect 10364 7516 10428 7520
rect 15012 7644 15076 7648
rect 15012 7588 15016 7644
rect 15016 7588 15072 7644
rect 15072 7588 15076 7644
rect 15012 7584 15076 7588
rect 15092 7644 15156 7648
rect 15092 7588 15096 7644
rect 15096 7588 15152 7644
rect 15152 7588 15156 7644
rect 15092 7584 15156 7588
rect 15172 7644 15236 7648
rect 15172 7588 15176 7644
rect 15176 7588 15232 7644
rect 15232 7588 15236 7644
rect 15172 7584 15236 7588
rect 15252 7644 15316 7648
rect 15252 7588 15256 7644
rect 15256 7588 15312 7644
rect 15312 7588 15316 7644
rect 15252 7584 15316 7588
rect 21012 7644 21076 7648
rect 21012 7588 21016 7644
rect 21016 7588 21072 7644
rect 21072 7588 21076 7644
rect 21012 7584 21076 7588
rect 21092 7644 21156 7648
rect 21092 7588 21096 7644
rect 21096 7588 21152 7644
rect 21152 7588 21156 7644
rect 21092 7584 21156 7588
rect 21172 7644 21236 7648
rect 21172 7588 21176 7644
rect 21176 7588 21232 7644
rect 21232 7588 21236 7644
rect 21172 7584 21236 7588
rect 21252 7644 21316 7648
rect 21252 7588 21256 7644
rect 21256 7588 21312 7644
rect 21312 7588 21316 7644
rect 21252 7584 21316 7588
rect 27012 7644 27076 7648
rect 27012 7588 27016 7644
rect 27016 7588 27072 7644
rect 27072 7588 27076 7644
rect 27012 7584 27076 7588
rect 27092 7644 27156 7648
rect 27092 7588 27096 7644
rect 27096 7588 27152 7644
rect 27152 7588 27156 7644
rect 27092 7584 27156 7588
rect 27172 7644 27236 7648
rect 27172 7588 27176 7644
rect 27176 7588 27232 7644
rect 27232 7588 27236 7644
rect 27172 7584 27236 7588
rect 27252 7644 27316 7648
rect 27252 7588 27256 7644
rect 27256 7588 27312 7644
rect 27312 7588 27316 7644
rect 27252 7584 27316 7588
rect 33012 7644 33076 7648
rect 33012 7588 33016 7644
rect 33016 7588 33072 7644
rect 33072 7588 33076 7644
rect 33012 7584 33076 7588
rect 33092 7644 33156 7648
rect 33092 7588 33096 7644
rect 33096 7588 33152 7644
rect 33152 7588 33156 7644
rect 33092 7584 33156 7588
rect 33172 7644 33236 7648
rect 33172 7588 33176 7644
rect 33176 7588 33232 7644
rect 33232 7588 33236 7644
rect 33172 7584 33236 7588
rect 33252 7644 33316 7648
rect 33252 7588 33256 7644
rect 33256 7588 33312 7644
rect 33312 7588 33316 7644
rect 33252 7584 33316 7588
rect 39012 7644 39076 7648
rect 39012 7588 39016 7644
rect 39016 7588 39072 7644
rect 39072 7588 39076 7644
rect 39012 7584 39076 7588
rect 39092 7644 39156 7648
rect 39092 7588 39096 7644
rect 39096 7588 39152 7644
rect 39152 7588 39156 7644
rect 39092 7584 39156 7588
rect 39172 7644 39236 7648
rect 39172 7588 39176 7644
rect 39176 7588 39232 7644
rect 39232 7588 39236 7644
rect 39172 7584 39236 7588
rect 39252 7644 39316 7648
rect 39252 7588 39256 7644
rect 39256 7588 39312 7644
rect 39312 7588 39316 7644
rect 39252 7584 39316 7588
rect 31340 7516 31404 7580
rect 32628 7516 32692 7580
rect 8708 7244 8772 7308
rect 1952 7100 2016 7104
rect 1952 7044 1956 7100
rect 1956 7044 2012 7100
rect 2012 7044 2016 7100
rect 1952 7040 2016 7044
rect 2032 7100 2096 7104
rect 2032 7044 2036 7100
rect 2036 7044 2092 7100
rect 2092 7044 2096 7100
rect 2032 7040 2096 7044
rect 2112 7100 2176 7104
rect 2112 7044 2116 7100
rect 2116 7044 2172 7100
rect 2172 7044 2176 7100
rect 2112 7040 2176 7044
rect 2192 7100 2256 7104
rect 2192 7044 2196 7100
rect 2196 7044 2252 7100
rect 2252 7044 2256 7100
rect 2192 7040 2256 7044
rect 3924 6972 3988 7036
rect 6684 6972 6748 7036
rect 8524 7108 8588 7172
rect 14780 7108 14844 7172
rect 16252 7108 16316 7172
rect 7952 7100 8016 7104
rect 7952 7044 7956 7100
rect 7956 7044 8012 7100
rect 8012 7044 8016 7100
rect 7952 7040 8016 7044
rect 8032 7100 8096 7104
rect 8032 7044 8036 7100
rect 8036 7044 8092 7100
rect 8092 7044 8096 7100
rect 8032 7040 8096 7044
rect 8112 7100 8176 7104
rect 8112 7044 8116 7100
rect 8116 7044 8172 7100
rect 8172 7044 8176 7100
rect 8112 7040 8176 7044
rect 8192 7100 8256 7104
rect 8192 7044 8196 7100
rect 8196 7044 8252 7100
rect 8252 7044 8256 7100
rect 8192 7040 8256 7044
rect 13952 7100 14016 7104
rect 13952 7044 13956 7100
rect 13956 7044 14012 7100
rect 14012 7044 14016 7100
rect 13952 7040 14016 7044
rect 14032 7100 14096 7104
rect 14032 7044 14036 7100
rect 14036 7044 14092 7100
rect 14092 7044 14096 7100
rect 14032 7040 14096 7044
rect 14112 7100 14176 7104
rect 14112 7044 14116 7100
rect 14116 7044 14172 7100
rect 14172 7044 14176 7100
rect 14112 7040 14176 7044
rect 14192 7100 14256 7104
rect 14192 7044 14196 7100
rect 14196 7044 14252 7100
rect 14252 7044 14256 7100
rect 14192 7040 14256 7044
rect 19952 7100 20016 7104
rect 19952 7044 19956 7100
rect 19956 7044 20012 7100
rect 20012 7044 20016 7100
rect 19952 7040 20016 7044
rect 20032 7100 20096 7104
rect 20032 7044 20036 7100
rect 20036 7044 20092 7100
rect 20092 7044 20096 7100
rect 20032 7040 20096 7044
rect 20112 7100 20176 7104
rect 20112 7044 20116 7100
rect 20116 7044 20172 7100
rect 20172 7044 20176 7100
rect 20112 7040 20176 7044
rect 20192 7100 20256 7104
rect 20192 7044 20196 7100
rect 20196 7044 20252 7100
rect 20252 7044 20256 7100
rect 20192 7040 20256 7044
rect 15884 7032 15948 7036
rect 15884 6976 15934 7032
rect 15934 6976 15948 7032
rect 15884 6972 15948 6976
rect 18644 6972 18708 7036
rect 25952 7100 26016 7104
rect 25952 7044 25956 7100
rect 25956 7044 26012 7100
rect 26012 7044 26016 7100
rect 25952 7040 26016 7044
rect 26032 7100 26096 7104
rect 26032 7044 26036 7100
rect 26036 7044 26092 7100
rect 26092 7044 26096 7100
rect 26032 7040 26096 7044
rect 26112 7100 26176 7104
rect 26112 7044 26116 7100
rect 26116 7044 26172 7100
rect 26172 7044 26176 7100
rect 26112 7040 26176 7044
rect 26192 7100 26256 7104
rect 26192 7044 26196 7100
rect 26196 7044 26252 7100
rect 26252 7044 26256 7100
rect 26192 7040 26256 7044
rect 31952 7100 32016 7104
rect 31952 7044 31956 7100
rect 31956 7044 32012 7100
rect 32012 7044 32016 7100
rect 31952 7040 32016 7044
rect 32032 7100 32096 7104
rect 32032 7044 32036 7100
rect 32036 7044 32092 7100
rect 32092 7044 32096 7100
rect 32032 7040 32096 7044
rect 32112 7100 32176 7104
rect 32112 7044 32116 7100
rect 32116 7044 32172 7100
rect 32172 7044 32176 7100
rect 32112 7040 32176 7044
rect 32192 7100 32256 7104
rect 32192 7044 32196 7100
rect 32196 7044 32252 7100
rect 32252 7044 32256 7100
rect 32192 7040 32256 7044
rect 37952 7100 38016 7104
rect 37952 7044 37956 7100
rect 37956 7044 38012 7100
rect 38012 7044 38016 7100
rect 37952 7040 38016 7044
rect 38032 7100 38096 7104
rect 38032 7044 38036 7100
rect 38036 7044 38092 7100
rect 38092 7044 38096 7100
rect 38032 7040 38096 7044
rect 38112 7100 38176 7104
rect 38112 7044 38116 7100
rect 38116 7044 38172 7100
rect 38172 7044 38176 7100
rect 38112 7040 38176 7044
rect 38192 7100 38256 7104
rect 38192 7044 38196 7100
rect 38196 7044 38252 7100
rect 38252 7044 38256 7100
rect 38192 7040 38256 7044
rect 26740 6972 26804 7036
rect 23428 6896 23492 6900
rect 23428 6840 23478 6896
rect 23478 6840 23492 6896
rect 23428 6836 23492 6840
rect 25636 6836 25700 6900
rect 5396 6624 5460 6628
rect 5396 6568 5446 6624
rect 5446 6568 5460 6624
rect 5396 6564 5460 6568
rect 3012 6556 3076 6560
rect 3012 6500 3016 6556
rect 3016 6500 3072 6556
rect 3072 6500 3076 6556
rect 3012 6496 3076 6500
rect 3092 6556 3156 6560
rect 3092 6500 3096 6556
rect 3096 6500 3152 6556
rect 3152 6500 3156 6556
rect 3092 6496 3156 6500
rect 3172 6556 3236 6560
rect 3172 6500 3176 6556
rect 3176 6500 3232 6556
rect 3232 6500 3236 6556
rect 3172 6496 3236 6500
rect 3252 6556 3316 6560
rect 3252 6500 3256 6556
rect 3256 6500 3312 6556
rect 3312 6500 3316 6556
rect 3252 6496 3316 6500
rect 2452 6292 2516 6356
rect 9012 6556 9076 6560
rect 9012 6500 9016 6556
rect 9016 6500 9072 6556
rect 9072 6500 9076 6556
rect 9012 6496 9076 6500
rect 9092 6556 9156 6560
rect 9092 6500 9096 6556
rect 9096 6500 9152 6556
rect 9152 6500 9156 6556
rect 9092 6496 9156 6500
rect 9172 6556 9236 6560
rect 9172 6500 9176 6556
rect 9176 6500 9232 6556
rect 9232 6500 9236 6556
rect 9172 6496 9236 6500
rect 9252 6556 9316 6560
rect 9252 6500 9256 6556
rect 9256 6500 9312 6556
rect 9312 6500 9316 6556
rect 9252 6496 9316 6500
rect 15012 6556 15076 6560
rect 15012 6500 15016 6556
rect 15016 6500 15072 6556
rect 15072 6500 15076 6556
rect 15012 6496 15076 6500
rect 15092 6556 15156 6560
rect 15092 6500 15096 6556
rect 15096 6500 15152 6556
rect 15152 6500 15156 6556
rect 15092 6496 15156 6500
rect 15172 6556 15236 6560
rect 15172 6500 15176 6556
rect 15176 6500 15232 6556
rect 15232 6500 15236 6556
rect 15172 6496 15236 6500
rect 15252 6556 15316 6560
rect 15252 6500 15256 6556
rect 15256 6500 15312 6556
rect 15312 6500 15316 6556
rect 15252 6496 15316 6500
rect 16068 6488 16132 6492
rect 21012 6556 21076 6560
rect 21012 6500 21016 6556
rect 21016 6500 21072 6556
rect 21072 6500 21076 6556
rect 21012 6496 21076 6500
rect 21092 6556 21156 6560
rect 21092 6500 21096 6556
rect 21096 6500 21152 6556
rect 21152 6500 21156 6556
rect 21092 6496 21156 6500
rect 21172 6556 21236 6560
rect 21172 6500 21176 6556
rect 21176 6500 21232 6556
rect 21232 6500 21236 6556
rect 21172 6496 21236 6500
rect 21252 6556 21316 6560
rect 21252 6500 21256 6556
rect 21256 6500 21312 6556
rect 21312 6500 21316 6556
rect 21252 6496 21316 6500
rect 16068 6432 16082 6488
rect 16082 6432 16132 6488
rect 16068 6428 16132 6432
rect 19012 6488 19076 6492
rect 19012 6432 19062 6488
rect 19062 6432 19076 6488
rect 19012 6428 19076 6432
rect 24900 6428 24964 6492
rect 27012 6556 27076 6560
rect 27012 6500 27016 6556
rect 27016 6500 27072 6556
rect 27072 6500 27076 6556
rect 27012 6496 27076 6500
rect 27092 6556 27156 6560
rect 27092 6500 27096 6556
rect 27096 6500 27152 6556
rect 27152 6500 27156 6556
rect 27092 6496 27156 6500
rect 27172 6556 27236 6560
rect 27172 6500 27176 6556
rect 27176 6500 27232 6556
rect 27232 6500 27236 6556
rect 27172 6496 27236 6500
rect 27252 6556 27316 6560
rect 27252 6500 27256 6556
rect 27256 6500 27312 6556
rect 27312 6500 27316 6556
rect 27252 6496 27316 6500
rect 33012 6556 33076 6560
rect 33012 6500 33016 6556
rect 33016 6500 33072 6556
rect 33072 6500 33076 6556
rect 33012 6496 33076 6500
rect 33092 6556 33156 6560
rect 33092 6500 33096 6556
rect 33096 6500 33152 6556
rect 33152 6500 33156 6556
rect 33092 6496 33156 6500
rect 33172 6556 33236 6560
rect 33172 6500 33176 6556
rect 33176 6500 33232 6556
rect 33232 6500 33236 6556
rect 33172 6496 33236 6500
rect 33252 6556 33316 6560
rect 33252 6500 33256 6556
rect 33256 6500 33312 6556
rect 33312 6500 33316 6556
rect 33252 6496 33316 6500
rect 39012 6556 39076 6560
rect 39012 6500 39016 6556
rect 39016 6500 39072 6556
rect 39072 6500 39076 6556
rect 39012 6496 39076 6500
rect 39092 6556 39156 6560
rect 39092 6500 39096 6556
rect 39096 6500 39152 6556
rect 39152 6500 39156 6556
rect 39092 6496 39156 6500
rect 39172 6556 39236 6560
rect 39172 6500 39176 6556
rect 39176 6500 39232 6556
rect 39232 6500 39236 6556
rect 39172 6496 39236 6500
rect 39252 6556 39316 6560
rect 39252 6500 39256 6556
rect 39256 6500 39312 6556
rect 39312 6500 39316 6556
rect 39252 6496 39316 6500
rect 31340 6428 31404 6492
rect 18276 6292 18340 6356
rect 28028 6292 28092 6356
rect 32444 6156 32508 6220
rect 16252 6020 16316 6084
rect 18276 6020 18340 6084
rect 1952 6012 2016 6016
rect 1952 5956 1956 6012
rect 1956 5956 2012 6012
rect 2012 5956 2016 6012
rect 1952 5952 2016 5956
rect 2032 6012 2096 6016
rect 2032 5956 2036 6012
rect 2036 5956 2092 6012
rect 2092 5956 2096 6012
rect 2032 5952 2096 5956
rect 2112 6012 2176 6016
rect 2112 5956 2116 6012
rect 2116 5956 2172 6012
rect 2172 5956 2176 6012
rect 2112 5952 2176 5956
rect 2192 6012 2256 6016
rect 2192 5956 2196 6012
rect 2196 5956 2252 6012
rect 2252 5956 2256 6012
rect 2192 5952 2256 5956
rect 7952 6012 8016 6016
rect 7952 5956 7956 6012
rect 7956 5956 8012 6012
rect 8012 5956 8016 6012
rect 7952 5952 8016 5956
rect 8032 6012 8096 6016
rect 8032 5956 8036 6012
rect 8036 5956 8092 6012
rect 8092 5956 8096 6012
rect 8032 5952 8096 5956
rect 8112 6012 8176 6016
rect 8112 5956 8116 6012
rect 8116 5956 8172 6012
rect 8172 5956 8176 6012
rect 8112 5952 8176 5956
rect 8192 6012 8256 6016
rect 8192 5956 8196 6012
rect 8196 5956 8252 6012
rect 8252 5956 8256 6012
rect 8192 5952 8256 5956
rect 13952 6012 14016 6016
rect 13952 5956 13956 6012
rect 13956 5956 14012 6012
rect 14012 5956 14016 6012
rect 13952 5952 14016 5956
rect 14032 6012 14096 6016
rect 14032 5956 14036 6012
rect 14036 5956 14092 6012
rect 14092 5956 14096 6012
rect 14032 5952 14096 5956
rect 14112 6012 14176 6016
rect 14112 5956 14116 6012
rect 14116 5956 14172 6012
rect 14172 5956 14176 6012
rect 14112 5952 14176 5956
rect 14192 6012 14256 6016
rect 14192 5956 14196 6012
rect 14196 5956 14252 6012
rect 14252 5956 14256 6012
rect 14192 5952 14256 5956
rect 19952 6012 20016 6016
rect 19952 5956 19956 6012
rect 19956 5956 20012 6012
rect 20012 5956 20016 6012
rect 19952 5952 20016 5956
rect 20032 6012 20096 6016
rect 20032 5956 20036 6012
rect 20036 5956 20092 6012
rect 20092 5956 20096 6012
rect 20032 5952 20096 5956
rect 20112 6012 20176 6016
rect 20112 5956 20116 6012
rect 20116 5956 20172 6012
rect 20172 5956 20176 6012
rect 20112 5952 20176 5956
rect 20192 6012 20256 6016
rect 20192 5956 20196 6012
rect 20196 5956 20252 6012
rect 20252 5956 20256 6012
rect 20192 5952 20256 5956
rect 25952 6012 26016 6016
rect 25952 5956 25956 6012
rect 25956 5956 26012 6012
rect 26012 5956 26016 6012
rect 25952 5952 26016 5956
rect 26032 6012 26096 6016
rect 26032 5956 26036 6012
rect 26036 5956 26092 6012
rect 26092 5956 26096 6012
rect 26032 5952 26096 5956
rect 26112 6012 26176 6016
rect 26112 5956 26116 6012
rect 26116 5956 26172 6012
rect 26172 5956 26176 6012
rect 26112 5952 26176 5956
rect 26192 6012 26256 6016
rect 26192 5956 26196 6012
rect 26196 5956 26252 6012
rect 26252 5956 26256 6012
rect 26192 5952 26256 5956
rect 31952 6012 32016 6016
rect 31952 5956 31956 6012
rect 31956 5956 32012 6012
rect 32012 5956 32016 6012
rect 31952 5952 32016 5956
rect 32032 6012 32096 6016
rect 32032 5956 32036 6012
rect 32036 5956 32092 6012
rect 32092 5956 32096 6012
rect 32032 5952 32096 5956
rect 32112 6012 32176 6016
rect 32112 5956 32116 6012
rect 32116 5956 32172 6012
rect 32172 5956 32176 6012
rect 32112 5952 32176 5956
rect 32192 6012 32256 6016
rect 32192 5956 32196 6012
rect 32196 5956 32252 6012
rect 32252 5956 32256 6012
rect 32192 5952 32256 5956
rect 37952 6012 38016 6016
rect 37952 5956 37956 6012
rect 37956 5956 38012 6012
rect 38012 5956 38016 6012
rect 37952 5952 38016 5956
rect 38032 6012 38096 6016
rect 38032 5956 38036 6012
rect 38036 5956 38092 6012
rect 38092 5956 38096 6012
rect 38032 5952 38096 5956
rect 38112 6012 38176 6016
rect 38112 5956 38116 6012
rect 38116 5956 38172 6012
rect 38172 5956 38176 6012
rect 38112 5952 38176 5956
rect 38192 6012 38256 6016
rect 38192 5956 38196 6012
rect 38196 5956 38252 6012
rect 38252 5956 38256 6012
rect 38192 5952 38256 5956
rect 2636 5884 2700 5948
rect 5580 5884 5644 5948
rect 14596 5884 14660 5948
rect 33732 5884 33796 5948
rect 8524 5476 8588 5540
rect 22140 5612 22204 5676
rect 37780 5612 37844 5676
rect 3012 5468 3076 5472
rect 3012 5412 3016 5468
rect 3016 5412 3072 5468
rect 3072 5412 3076 5468
rect 3012 5408 3076 5412
rect 3092 5468 3156 5472
rect 3092 5412 3096 5468
rect 3096 5412 3152 5468
rect 3152 5412 3156 5468
rect 3092 5408 3156 5412
rect 3172 5468 3236 5472
rect 3172 5412 3176 5468
rect 3176 5412 3232 5468
rect 3232 5412 3236 5468
rect 3172 5408 3236 5412
rect 3252 5468 3316 5472
rect 3252 5412 3256 5468
rect 3256 5412 3312 5468
rect 3312 5412 3316 5468
rect 3252 5408 3316 5412
rect 9012 5468 9076 5472
rect 9012 5412 9016 5468
rect 9016 5412 9072 5468
rect 9072 5412 9076 5468
rect 9012 5408 9076 5412
rect 9092 5468 9156 5472
rect 9092 5412 9096 5468
rect 9096 5412 9152 5468
rect 9152 5412 9156 5468
rect 9092 5408 9156 5412
rect 9172 5468 9236 5472
rect 9172 5412 9176 5468
rect 9176 5412 9232 5468
rect 9232 5412 9236 5468
rect 9172 5408 9236 5412
rect 9252 5468 9316 5472
rect 9252 5412 9256 5468
rect 9256 5412 9312 5468
rect 9312 5412 9316 5468
rect 9252 5408 9316 5412
rect 15012 5468 15076 5472
rect 15012 5412 15016 5468
rect 15016 5412 15072 5468
rect 15072 5412 15076 5468
rect 15012 5408 15076 5412
rect 15092 5468 15156 5472
rect 15092 5412 15096 5468
rect 15096 5412 15152 5468
rect 15152 5412 15156 5468
rect 15092 5408 15156 5412
rect 15172 5468 15236 5472
rect 15172 5412 15176 5468
rect 15176 5412 15232 5468
rect 15232 5412 15236 5468
rect 15172 5408 15236 5412
rect 15252 5468 15316 5472
rect 15252 5412 15256 5468
rect 15256 5412 15312 5468
rect 15312 5412 15316 5468
rect 15252 5408 15316 5412
rect 21012 5468 21076 5472
rect 21012 5412 21016 5468
rect 21016 5412 21072 5468
rect 21072 5412 21076 5468
rect 21012 5408 21076 5412
rect 21092 5468 21156 5472
rect 21092 5412 21096 5468
rect 21096 5412 21152 5468
rect 21152 5412 21156 5468
rect 21092 5408 21156 5412
rect 21172 5468 21236 5472
rect 21172 5412 21176 5468
rect 21176 5412 21232 5468
rect 21232 5412 21236 5468
rect 21172 5408 21236 5412
rect 21252 5468 21316 5472
rect 21252 5412 21256 5468
rect 21256 5412 21312 5468
rect 21312 5412 21316 5468
rect 21252 5408 21316 5412
rect 27012 5468 27076 5472
rect 27012 5412 27016 5468
rect 27016 5412 27072 5468
rect 27072 5412 27076 5468
rect 27012 5408 27076 5412
rect 27092 5468 27156 5472
rect 27092 5412 27096 5468
rect 27096 5412 27152 5468
rect 27152 5412 27156 5468
rect 27092 5408 27156 5412
rect 27172 5468 27236 5472
rect 27172 5412 27176 5468
rect 27176 5412 27232 5468
rect 27232 5412 27236 5468
rect 27172 5408 27236 5412
rect 27252 5468 27316 5472
rect 27252 5412 27256 5468
rect 27256 5412 27312 5468
rect 27312 5412 27316 5468
rect 27252 5408 27316 5412
rect 33012 5468 33076 5472
rect 33012 5412 33016 5468
rect 33016 5412 33072 5468
rect 33072 5412 33076 5468
rect 33012 5408 33076 5412
rect 33092 5468 33156 5472
rect 33092 5412 33096 5468
rect 33096 5412 33152 5468
rect 33152 5412 33156 5468
rect 33092 5408 33156 5412
rect 33172 5468 33236 5472
rect 33172 5412 33176 5468
rect 33176 5412 33232 5468
rect 33232 5412 33236 5468
rect 33172 5408 33236 5412
rect 33252 5468 33316 5472
rect 33252 5412 33256 5468
rect 33256 5412 33312 5468
rect 33312 5412 33316 5468
rect 33252 5408 33316 5412
rect 39012 5468 39076 5472
rect 39012 5412 39016 5468
rect 39016 5412 39072 5468
rect 39072 5412 39076 5468
rect 39012 5408 39076 5412
rect 39092 5468 39156 5472
rect 39092 5412 39096 5468
rect 39096 5412 39152 5468
rect 39152 5412 39156 5468
rect 39092 5408 39156 5412
rect 39172 5468 39236 5472
rect 39172 5412 39176 5468
rect 39176 5412 39232 5468
rect 39232 5412 39236 5468
rect 39172 5408 39236 5412
rect 39252 5468 39316 5472
rect 39252 5412 39256 5468
rect 39256 5412 39312 5468
rect 39312 5412 39316 5468
rect 39252 5408 39316 5412
rect 7052 5400 7116 5404
rect 7052 5344 7066 5400
rect 7066 5344 7116 5400
rect 7052 5340 7116 5344
rect 8708 5340 8772 5404
rect 9812 5204 9876 5268
rect 18460 5204 18524 5268
rect 8524 4932 8588 4996
rect 1952 4924 2016 4928
rect 1952 4868 1956 4924
rect 1956 4868 2012 4924
rect 2012 4868 2016 4924
rect 1952 4864 2016 4868
rect 2032 4924 2096 4928
rect 2032 4868 2036 4924
rect 2036 4868 2092 4924
rect 2092 4868 2096 4924
rect 2032 4864 2096 4868
rect 2112 4924 2176 4928
rect 2112 4868 2116 4924
rect 2116 4868 2172 4924
rect 2172 4868 2176 4924
rect 2112 4864 2176 4868
rect 2192 4924 2256 4928
rect 2192 4868 2196 4924
rect 2196 4868 2252 4924
rect 2252 4868 2256 4924
rect 2192 4864 2256 4868
rect 7952 4924 8016 4928
rect 7952 4868 7956 4924
rect 7956 4868 8012 4924
rect 8012 4868 8016 4924
rect 7952 4864 8016 4868
rect 8032 4924 8096 4928
rect 8032 4868 8036 4924
rect 8036 4868 8092 4924
rect 8092 4868 8096 4924
rect 8032 4864 8096 4868
rect 8112 4924 8176 4928
rect 8112 4868 8116 4924
rect 8116 4868 8172 4924
rect 8172 4868 8176 4924
rect 8112 4864 8176 4868
rect 8192 4924 8256 4928
rect 8192 4868 8196 4924
rect 8196 4868 8252 4924
rect 8252 4868 8256 4924
rect 8192 4864 8256 4868
rect 13952 4924 14016 4928
rect 13952 4868 13956 4924
rect 13956 4868 14012 4924
rect 14012 4868 14016 4924
rect 13952 4864 14016 4868
rect 14032 4924 14096 4928
rect 14032 4868 14036 4924
rect 14036 4868 14092 4924
rect 14092 4868 14096 4924
rect 14032 4864 14096 4868
rect 14112 4924 14176 4928
rect 14112 4868 14116 4924
rect 14116 4868 14172 4924
rect 14172 4868 14176 4924
rect 14112 4864 14176 4868
rect 14192 4924 14256 4928
rect 14192 4868 14196 4924
rect 14196 4868 14252 4924
rect 14252 4868 14256 4924
rect 14192 4864 14256 4868
rect 19952 4924 20016 4928
rect 19952 4868 19956 4924
rect 19956 4868 20012 4924
rect 20012 4868 20016 4924
rect 19952 4864 20016 4868
rect 20032 4924 20096 4928
rect 20032 4868 20036 4924
rect 20036 4868 20092 4924
rect 20092 4868 20096 4924
rect 20032 4864 20096 4868
rect 20112 4924 20176 4928
rect 20112 4868 20116 4924
rect 20116 4868 20172 4924
rect 20172 4868 20176 4924
rect 20112 4864 20176 4868
rect 20192 4924 20256 4928
rect 20192 4868 20196 4924
rect 20196 4868 20252 4924
rect 20252 4868 20256 4924
rect 20192 4864 20256 4868
rect 25952 4924 26016 4928
rect 25952 4868 25956 4924
rect 25956 4868 26012 4924
rect 26012 4868 26016 4924
rect 25952 4864 26016 4868
rect 26032 4924 26096 4928
rect 26032 4868 26036 4924
rect 26036 4868 26092 4924
rect 26092 4868 26096 4924
rect 26032 4864 26096 4868
rect 26112 4924 26176 4928
rect 26112 4868 26116 4924
rect 26116 4868 26172 4924
rect 26172 4868 26176 4924
rect 26112 4864 26176 4868
rect 26192 4924 26256 4928
rect 26192 4868 26196 4924
rect 26196 4868 26252 4924
rect 26252 4868 26256 4924
rect 26192 4864 26256 4868
rect 31952 4924 32016 4928
rect 31952 4868 31956 4924
rect 31956 4868 32012 4924
rect 32012 4868 32016 4924
rect 31952 4864 32016 4868
rect 32032 4924 32096 4928
rect 32032 4868 32036 4924
rect 32036 4868 32092 4924
rect 32092 4868 32096 4924
rect 32032 4864 32096 4868
rect 32112 4924 32176 4928
rect 32112 4868 32116 4924
rect 32116 4868 32172 4924
rect 32172 4868 32176 4924
rect 32112 4864 32176 4868
rect 32192 4924 32256 4928
rect 32192 4868 32196 4924
rect 32196 4868 32252 4924
rect 32252 4868 32256 4924
rect 32192 4864 32256 4868
rect 37952 4924 38016 4928
rect 37952 4868 37956 4924
rect 37956 4868 38012 4924
rect 38012 4868 38016 4924
rect 37952 4864 38016 4868
rect 38032 4924 38096 4928
rect 38032 4868 38036 4924
rect 38036 4868 38092 4924
rect 38092 4868 38096 4924
rect 38032 4864 38096 4868
rect 38112 4924 38176 4928
rect 38112 4868 38116 4924
rect 38116 4868 38172 4924
rect 38172 4868 38176 4924
rect 38112 4864 38176 4868
rect 38192 4924 38256 4928
rect 38192 4868 38196 4924
rect 38196 4868 38252 4924
rect 38252 4868 38256 4924
rect 38192 4864 38256 4868
rect 30604 4856 30668 4860
rect 30604 4800 30618 4856
rect 30618 4800 30668 4856
rect 30604 4796 30668 4800
rect 14780 4448 14844 4452
rect 14780 4392 14794 4448
rect 14794 4392 14844 4448
rect 14780 4388 14844 4392
rect 3012 4380 3076 4384
rect 3012 4324 3016 4380
rect 3016 4324 3072 4380
rect 3072 4324 3076 4380
rect 3012 4320 3076 4324
rect 3092 4380 3156 4384
rect 3092 4324 3096 4380
rect 3096 4324 3152 4380
rect 3152 4324 3156 4380
rect 3092 4320 3156 4324
rect 3172 4380 3236 4384
rect 3172 4324 3176 4380
rect 3176 4324 3232 4380
rect 3232 4324 3236 4380
rect 3172 4320 3236 4324
rect 3252 4380 3316 4384
rect 3252 4324 3256 4380
rect 3256 4324 3312 4380
rect 3312 4324 3316 4380
rect 3252 4320 3316 4324
rect 9012 4380 9076 4384
rect 9012 4324 9016 4380
rect 9016 4324 9072 4380
rect 9072 4324 9076 4380
rect 9012 4320 9076 4324
rect 9092 4380 9156 4384
rect 9092 4324 9096 4380
rect 9096 4324 9152 4380
rect 9152 4324 9156 4380
rect 9092 4320 9156 4324
rect 9172 4380 9236 4384
rect 9172 4324 9176 4380
rect 9176 4324 9232 4380
rect 9232 4324 9236 4380
rect 9172 4320 9236 4324
rect 9252 4380 9316 4384
rect 9252 4324 9256 4380
rect 9256 4324 9312 4380
rect 9312 4324 9316 4380
rect 9252 4320 9316 4324
rect 15012 4380 15076 4384
rect 15012 4324 15016 4380
rect 15016 4324 15072 4380
rect 15072 4324 15076 4380
rect 15012 4320 15076 4324
rect 15092 4380 15156 4384
rect 15092 4324 15096 4380
rect 15096 4324 15152 4380
rect 15152 4324 15156 4380
rect 15092 4320 15156 4324
rect 15172 4380 15236 4384
rect 15172 4324 15176 4380
rect 15176 4324 15232 4380
rect 15232 4324 15236 4380
rect 15172 4320 15236 4324
rect 15252 4380 15316 4384
rect 15252 4324 15256 4380
rect 15256 4324 15312 4380
rect 15312 4324 15316 4380
rect 15252 4320 15316 4324
rect 21012 4380 21076 4384
rect 21012 4324 21016 4380
rect 21016 4324 21072 4380
rect 21072 4324 21076 4380
rect 21012 4320 21076 4324
rect 21092 4380 21156 4384
rect 21092 4324 21096 4380
rect 21096 4324 21152 4380
rect 21152 4324 21156 4380
rect 21092 4320 21156 4324
rect 21172 4380 21236 4384
rect 21172 4324 21176 4380
rect 21176 4324 21232 4380
rect 21232 4324 21236 4380
rect 21172 4320 21236 4324
rect 21252 4380 21316 4384
rect 21252 4324 21256 4380
rect 21256 4324 21312 4380
rect 21312 4324 21316 4380
rect 21252 4320 21316 4324
rect 27012 4380 27076 4384
rect 27012 4324 27016 4380
rect 27016 4324 27072 4380
rect 27072 4324 27076 4380
rect 27012 4320 27076 4324
rect 27092 4380 27156 4384
rect 27092 4324 27096 4380
rect 27096 4324 27152 4380
rect 27152 4324 27156 4380
rect 27092 4320 27156 4324
rect 27172 4380 27236 4384
rect 27172 4324 27176 4380
rect 27176 4324 27232 4380
rect 27232 4324 27236 4380
rect 27172 4320 27236 4324
rect 27252 4380 27316 4384
rect 27252 4324 27256 4380
rect 27256 4324 27312 4380
rect 27312 4324 27316 4380
rect 27252 4320 27316 4324
rect 33012 4380 33076 4384
rect 33012 4324 33016 4380
rect 33016 4324 33072 4380
rect 33072 4324 33076 4380
rect 33012 4320 33076 4324
rect 33092 4380 33156 4384
rect 33092 4324 33096 4380
rect 33096 4324 33152 4380
rect 33152 4324 33156 4380
rect 33092 4320 33156 4324
rect 33172 4380 33236 4384
rect 33172 4324 33176 4380
rect 33176 4324 33232 4380
rect 33232 4324 33236 4380
rect 33172 4320 33236 4324
rect 33252 4380 33316 4384
rect 33252 4324 33256 4380
rect 33256 4324 33312 4380
rect 33312 4324 33316 4380
rect 33252 4320 33316 4324
rect 39012 4380 39076 4384
rect 39012 4324 39016 4380
rect 39016 4324 39072 4380
rect 39072 4324 39076 4380
rect 39012 4320 39076 4324
rect 39092 4380 39156 4384
rect 39092 4324 39096 4380
rect 39096 4324 39152 4380
rect 39152 4324 39156 4380
rect 39092 4320 39156 4324
rect 39172 4380 39236 4384
rect 39172 4324 39176 4380
rect 39176 4324 39232 4380
rect 39232 4324 39236 4380
rect 39172 4320 39236 4324
rect 39252 4380 39316 4384
rect 39252 4324 39256 4380
rect 39256 4324 39312 4380
rect 39312 4324 39316 4380
rect 39252 4320 39316 4324
rect 7052 4116 7116 4180
rect 10916 4252 10980 4316
rect 16068 4176 16132 4180
rect 16068 4120 16082 4176
rect 16082 4120 16132 4176
rect 16068 4116 16132 4120
rect 32812 4116 32876 4180
rect 5396 3904 5460 3908
rect 5396 3848 5410 3904
rect 5410 3848 5460 3904
rect 5396 3844 5460 3848
rect 9812 3844 9876 3908
rect 15884 3844 15948 3908
rect 1952 3836 2016 3840
rect 1952 3780 1956 3836
rect 1956 3780 2012 3836
rect 2012 3780 2016 3836
rect 1952 3776 2016 3780
rect 2032 3836 2096 3840
rect 2032 3780 2036 3836
rect 2036 3780 2092 3836
rect 2092 3780 2096 3836
rect 2032 3776 2096 3780
rect 2112 3836 2176 3840
rect 2112 3780 2116 3836
rect 2116 3780 2172 3836
rect 2172 3780 2176 3836
rect 2112 3776 2176 3780
rect 2192 3836 2256 3840
rect 2192 3780 2196 3836
rect 2196 3780 2252 3836
rect 2252 3780 2256 3836
rect 2192 3776 2256 3780
rect 7952 3836 8016 3840
rect 7952 3780 7956 3836
rect 7956 3780 8012 3836
rect 8012 3780 8016 3836
rect 7952 3776 8016 3780
rect 8032 3836 8096 3840
rect 8032 3780 8036 3836
rect 8036 3780 8092 3836
rect 8092 3780 8096 3836
rect 8032 3776 8096 3780
rect 8112 3836 8176 3840
rect 8112 3780 8116 3836
rect 8116 3780 8172 3836
rect 8172 3780 8176 3836
rect 8112 3776 8176 3780
rect 8192 3836 8256 3840
rect 8192 3780 8196 3836
rect 8196 3780 8252 3836
rect 8252 3780 8256 3836
rect 8192 3776 8256 3780
rect 13952 3836 14016 3840
rect 13952 3780 13956 3836
rect 13956 3780 14012 3836
rect 14012 3780 14016 3836
rect 13952 3776 14016 3780
rect 14032 3836 14096 3840
rect 14032 3780 14036 3836
rect 14036 3780 14092 3836
rect 14092 3780 14096 3836
rect 14032 3776 14096 3780
rect 14112 3836 14176 3840
rect 14112 3780 14116 3836
rect 14116 3780 14172 3836
rect 14172 3780 14176 3836
rect 14112 3776 14176 3780
rect 14192 3836 14256 3840
rect 14192 3780 14196 3836
rect 14196 3780 14252 3836
rect 14252 3780 14256 3836
rect 14192 3776 14256 3780
rect 19952 3836 20016 3840
rect 19952 3780 19956 3836
rect 19956 3780 20012 3836
rect 20012 3780 20016 3836
rect 19952 3776 20016 3780
rect 20032 3836 20096 3840
rect 20032 3780 20036 3836
rect 20036 3780 20092 3836
rect 20092 3780 20096 3836
rect 20032 3776 20096 3780
rect 20112 3836 20176 3840
rect 20112 3780 20116 3836
rect 20116 3780 20172 3836
rect 20172 3780 20176 3836
rect 20112 3776 20176 3780
rect 20192 3836 20256 3840
rect 20192 3780 20196 3836
rect 20196 3780 20252 3836
rect 20252 3780 20256 3836
rect 20192 3776 20256 3780
rect 25952 3836 26016 3840
rect 25952 3780 25956 3836
rect 25956 3780 26012 3836
rect 26012 3780 26016 3836
rect 25952 3776 26016 3780
rect 26032 3836 26096 3840
rect 26032 3780 26036 3836
rect 26036 3780 26092 3836
rect 26092 3780 26096 3836
rect 26032 3776 26096 3780
rect 26112 3836 26176 3840
rect 26112 3780 26116 3836
rect 26116 3780 26172 3836
rect 26172 3780 26176 3836
rect 26112 3776 26176 3780
rect 26192 3836 26256 3840
rect 26192 3780 26196 3836
rect 26196 3780 26252 3836
rect 26252 3780 26256 3836
rect 26192 3776 26256 3780
rect 31952 3836 32016 3840
rect 31952 3780 31956 3836
rect 31956 3780 32012 3836
rect 32012 3780 32016 3836
rect 31952 3776 32016 3780
rect 32032 3836 32096 3840
rect 32032 3780 32036 3836
rect 32036 3780 32092 3836
rect 32092 3780 32096 3836
rect 32032 3776 32096 3780
rect 32112 3836 32176 3840
rect 32112 3780 32116 3836
rect 32116 3780 32172 3836
rect 32172 3780 32176 3836
rect 32112 3776 32176 3780
rect 32192 3836 32256 3840
rect 32192 3780 32196 3836
rect 32196 3780 32252 3836
rect 32252 3780 32256 3836
rect 32192 3776 32256 3780
rect 37952 3836 38016 3840
rect 37952 3780 37956 3836
rect 37956 3780 38012 3836
rect 38012 3780 38016 3836
rect 37952 3776 38016 3780
rect 38032 3836 38096 3840
rect 38032 3780 38036 3836
rect 38036 3780 38092 3836
rect 38092 3780 38096 3836
rect 38032 3776 38096 3780
rect 38112 3836 38176 3840
rect 38112 3780 38116 3836
rect 38116 3780 38172 3836
rect 38172 3780 38176 3836
rect 38112 3776 38176 3780
rect 38192 3836 38256 3840
rect 38192 3780 38196 3836
rect 38196 3780 38252 3836
rect 38252 3780 38256 3836
rect 38192 3776 38256 3780
rect 7604 3708 7668 3772
rect 15516 3708 15580 3772
rect 16804 3708 16868 3772
rect 9628 3572 9692 3636
rect 17908 3436 17972 3500
rect 3012 3292 3076 3296
rect 3012 3236 3016 3292
rect 3016 3236 3072 3292
rect 3072 3236 3076 3292
rect 3012 3232 3076 3236
rect 3092 3292 3156 3296
rect 3092 3236 3096 3292
rect 3096 3236 3152 3292
rect 3152 3236 3156 3292
rect 3092 3232 3156 3236
rect 3172 3292 3236 3296
rect 3172 3236 3176 3292
rect 3176 3236 3232 3292
rect 3232 3236 3236 3292
rect 3172 3232 3236 3236
rect 3252 3292 3316 3296
rect 3252 3236 3256 3292
rect 3256 3236 3312 3292
rect 3312 3236 3316 3292
rect 3252 3232 3316 3236
rect 9012 3292 9076 3296
rect 9012 3236 9016 3292
rect 9016 3236 9072 3292
rect 9072 3236 9076 3292
rect 9012 3232 9076 3236
rect 9092 3292 9156 3296
rect 9092 3236 9096 3292
rect 9096 3236 9152 3292
rect 9152 3236 9156 3292
rect 9092 3232 9156 3236
rect 9172 3292 9236 3296
rect 9172 3236 9176 3292
rect 9176 3236 9232 3292
rect 9232 3236 9236 3292
rect 9172 3232 9236 3236
rect 9252 3292 9316 3296
rect 9252 3236 9256 3292
rect 9256 3236 9312 3292
rect 9312 3236 9316 3292
rect 9252 3232 9316 3236
rect 15012 3292 15076 3296
rect 15012 3236 15016 3292
rect 15016 3236 15072 3292
rect 15072 3236 15076 3292
rect 15012 3232 15076 3236
rect 15092 3292 15156 3296
rect 15092 3236 15096 3292
rect 15096 3236 15152 3292
rect 15152 3236 15156 3292
rect 15092 3232 15156 3236
rect 15172 3292 15236 3296
rect 15172 3236 15176 3292
rect 15176 3236 15232 3292
rect 15232 3236 15236 3292
rect 15172 3232 15236 3236
rect 15252 3292 15316 3296
rect 15252 3236 15256 3292
rect 15256 3236 15312 3292
rect 15312 3236 15316 3292
rect 15252 3232 15316 3236
rect 21012 3292 21076 3296
rect 21012 3236 21016 3292
rect 21016 3236 21072 3292
rect 21072 3236 21076 3292
rect 21012 3232 21076 3236
rect 21092 3292 21156 3296
rect 21092 3236 21096 3292
rect 21096 3236 21152 3292
rect 21152 3236 21156 3292
rect 21092 3232 21156 3236
rect 21172 3292 21236 3296
rect 21172 3236 21176 3292
rect 21176 3236 21232 3292
rect 21232 3236 21236 3292
rect 21172 3232 21236 3236
rect 21252 3292 21316 3296
rect 21252 3236 21256 3292
rect 21256 3236 21312 3292
rect 21312 3236 21316 3292
rect 21252 3232 21316 3236
rect 27012 3292 27076 3296
rect 27012 3236 27016 3292
rect 27016 3236 27072 3292
rect 27072 3236 27076 3292
rect 27012 3232 27076 3236
rect 27092 3292 27156 3296
rect 27092 3236 27096 3292
rect 27096 3236 27152 3292
rect 27152 3236 27156 3292
rect 27092 3232 27156 3236
rect 27172 3292 27236 3296
rect 27172 3236 27176 3292
rect 27176 3236 27232 3292
rect 27232 3236 27236 3292
rect 27172 3232 27236 3236
rect 27252 3292 27316 3296
rect 27252 3236 27256 3292
rect 27256 3236 27312 3292
rect 27312 3236 27316 3292
rect 27252 3232 27316 3236
rect 33012 3292 33076 3296
rect 33012 3236 33016 3292
rect 33016 3236 33072 3292
rect 33072 3236 33076 3292
rect 33012 3232 33076 3236
rect 33092 3292 33156 3296
rect 33092 3236 33096 3292
rect 33096 3236 33152 3292
rect 33152 3236 33156 3292
rect 33092 3232 33156 3236
rect 33172 3292 33236 3296
rect 33172 3236 33176 3292
rect 33176 3236 33232 3292
rect 33232 3236 33236 3292
rect 33172 3232 33236 3236
rect 33252 3292 33316 3296
rect 33252 3236 33256 3292
rect 33256 3236 33312 3292
rect 33312 3236 33316 3292
rect 33252 3232 33316 3236
rect 39012 3292 39076 3296
rect 39012 3236 39016 3292
rect 39016 3236 39072 3292
rect 39072 3236 39076 3292
rect 39012 3232 39076 3236
rect 39092 3292 39156 3296
rect 39092 3236 39096 3292
rect 39096 3236 39152 3292
rect 39152 3236 39156 3292
rect 39092 3232 39156 3236
rect 39172 3292 39236 3296
rect 39172 3236 39176 3292
rect 39176 3236 39232 3292
rect 39232 3236 39236 3292
rect 39172 3232 39236 3236
rect 39252 3292 39316 3296
rect 39252 3236 39256 3292
rect 39256 3236 39312 3292
rect 39312 3236 39316 3292
rect 39252 3232 39316 3236
rect 24164 3224 24228 3228
rect 24164 3168 24178 3224
rect 24178 3168 24228 3224
rect 24164 3164 24228 3168
rect 25452 3028 25516 3092
rect 26372 2892 26436 2956
rect 26556 2952 26620 2956
rect 26556 2896 26606 2952
rect 26606 2896 26620 2952
rect 26556 2892 26620 2896
rect 1952 2748 2016 2752
rect 1952 2692 1956 2748
rect 1956 2692 2012 2748
rect 2012 2692 2016 2748
rect 1952 2688 2016 2692
rect 2032 2748 2096 2752
rect 2032 2692 2036 2748
rect 2036 2692 2092 2748
rect 2092 2692 2096 2748
rect 2032 2688 2096 2692
rect 2112 2748 2176 2752
rect 2112 2692 2116 2748
rect 2116 2692 2172 2748
rect 2172 2692 2176 2748
rect 2112 2688 2176 2692
rect 2192 2748 2256 2752
rect 2192 2692 2196 2748
rect 2196 2692 2252 2748
rect 2252 2692 2256 2748
rect 2192 2688 2256 2692
rect 7952 2748 8016 2752
rect 7952 2692 7956 2748
rect 7956 2692 8012 2748
rect 8012 2692 8016 2748
rect 7952 2688 8016 2692
rect 8032 2748 8096 2752
rect 8032 2692 8036 2748
rect 8036 2692 8092 2748
rect 8092 2692 8096 2748
rect 8032 2688 8096 2692
rect 8112 2748 8176 2752
rect 8112 2692 8116 2748
rect 8116 2692 8172 2748
rect 8172 2692 8176 2748
rect 8112 2688 8176 2692
rect 8192 2748 8256 2752
rect 8192 2692 8196 2748
rect 8196 2692 8252 2748
rect 8252 2692 8256 2748
rect 8192 2688 8256 2692
rect 13952 2748 14016 2752
rect 13952 2692 13956 2748
rect 13956 2692 14012 2748
rect 14012 2692 14016 2748
rect 13952 2688 14016 2692
rect 14032 2748 14096 2752
rect 14032 2692 14036 2748
rect 14036 2692 14092 2748
rect 14092 2692 14096 2748
rect 14032 2688 14096 2692
rect 14112 2748 14176 2752
rect 14112 2692 14116 2748
rect 14116 2692 14172 2748
rect 14172 2692 14176 2748
rect 14112 2688 14176 2692
rect 14192 2748 14256 2752
rect 14192 2692 14196 2748
rect 14196 2692 14252 2748
rect 14252 2692 14256 2748
rect 14192 2688 14256 2692
rect 19952 2748 20016 2752
rect 19952 2692 19956 2748
rect 19956 2692 20012 2748
rect 20012 2692 20016 2748
rect 19952 2688 20016 2692
rect 20032 2748 20096 2752
rect 20032 2692 20036 2748
rect 20036 2692 20092 2748
rect 20092 2692 20096 2748
rect 20032 2688 20096 2692
rect 20112 2748 20176 2752
rect 20112 2692 20116 2748
rect 20116 2692 20172 2748
rect 20172 2692 20176 2748
rect 20112 2688 20176 2692
rect 20192 2748 20256 2752
rect 20192 2692 20196 2748
rect 20196 2692 20252 2748
rect 20252 2692 20256 2748
rect 20192 2688 20256 2692
rect 25952 2748 26016 2752
rect 25952 2692 25956 2748
rect 25956 2692 26012 2748
rect 26012 2692 26016 2748
rect 25952 2688 26016 2692
rect 26032 2748 26096 2752
rect 26032 2692 26036 2748
rect 26036 2692 26092 2748
rect 26092 2692 26096 2748
rect 26032 2688 26096 2692
rect 26112 2748 26176 2752
rect 26112 2692 26116 2748
rect 26116 2692 26172 2748
rect 26172 2692 26176 2748
rect 26112 2688 26176 2692
rect 26192 2748 26256 2752
rect 26192 2692 26196 2748
rect 26196 2692 26252 2748
rect 26252 2692 26256 2748
rect 26192 2688 26256 2692
rect 31952 2748 32016 2752
rect 31952 2692 31956 2748
rect 31956 2692 32012 2748
rect 32012 2692 32016 2748
rect 31952 2688 32016 2692
rect 32032 2748 32096 2752
rect 32032 2692 32036 2748
rect 32036 2692 32092 2748
rect 32092 2692 32096 2748
rect 32032 2688 32096 2692
rect 32112 2748 32176 2752
rect 32112 2692 32116 2748
rect 32116 2692 32172 2748
rect 32172 2692 32176 2748
rect 32112 2688 32176 2692
rect 32192 2748 32256 2752
rect 32192 2692 32196 2748
rect 32196 2692 32252 2748
rect 32252 2692 32256 2748
rect 32192 2688 32256 2692
rect 37952 2748 38016 2752
rect 37952 2692 37956 2748
rect 37956 2692 38012 2748
rect 38012 2692 38016 2748
rect 37952 2688 38016 2692
rect 38032 2748 38096 2752
rect 38032 2692 38036 2748
rect 38036 2692 38092 2748
rect 38092 2692 38096 2748
rect 38032 2688 38096 2692
rect 38112 2748 38176 2752
rect 38112 2692 38116 2748
rect 38116 2692 38172 2748
rect 38172 2692 38176 2748
rect 38112 2688 38176 2692
rect 38192 2748 38256 2752
rect 38192 2692 38196 2748
rect 38196 2692 38252 2748
rect 38252 2692 38256 2748
rect 38192 2688 38256 2692
rect 14596 2544 14660 2548
rect 14596 2488 14610 2544
rect 14610 2488 14660 2544
rect 14596 2484 14660 2488
rect 37780 2484 37844 2548
rect 10364 2272 10428 2276
rect 10364 2216 10378 2272
rect 10378 2216 10428 2272
rect 10364 2212 10428 2216
rect 3012 2204 3076 2208
rect 3012 2148 3016 2204
rect 3016 2148 3072 2204
rect 3072 2148 3076 2204
rect 3012 2144 3076 2148
rect 3092 2204 3156 2208
rect 3092 2148 3096 2204
rect 3096 2148 3152 2204
rect 3152 2148 3156 2204
rect 3092 2144 3156 2148
rect 3172 2204 3236 2208
rect 3172 2148 3176 2204
rect 3176 2148 3232 2204
rect 3232 2148 3236 2204
rect 3172 2144 3236 2148
rect 3252 2204 3316 2208
rect 3252 2148 3256 2204
rect 3256 2148 3312 2204
rect 3312 2148 3316 2204
rect 3252 2144 3316 2148
rect 9012 2204 9076 2208
rect 9012 2148 9016 2204
rect 9016 2148 9072 2204
rect 9072 2148 9076 2204
rect 9012 2144 9076 2148
rect 9092 2204 9156 2208
rect 9092 2148 9096 2204
rect 9096 2148 9152 2204
rect 9152 2148 9156 2204
rect 9092 2144 9156 2148
rect 9172 2204 9236 2208
rect 9172 2148 9176 2204
rect 9176 2148 9232 2204
rect 9232 2148 9236 2204
rect 9172 2144 9236 2148
rect 9252 2204 9316 2208
rect 9252 2148 9256 2204
rect 9256 2148 9312 2204
rect 9312 2148 9316 2204
rect 9252 2144 9316 2148
rect 15012 2204 15076 2208
rect 15012 2148 15016 2204
rect 15016 2148 15072 2204
rect 15072 2148 15076 2204
rect 15012 2144 15076 2148
rect 15092 2204 15156 2208
rect 15092 2148 15096 2204
rect 15096 2148 15152 2204
rect 15152 2148 15156 2204
rect 15092 2144 15156 2148
rect 15172 2204 15236 2208
rect 15172 2148 15176 2204
rect 15176 2148 15232 2204
rect 15232 2148 15236 2204
rect 15172 2144 15236 2148
rect 15252 2204 15316 2208
rect 15252 2148 15256 2204
rect 15256 2148 15312 2204
rect 15312 2148 15316 2204
rect 15252 2144 15316 2148
rect 21012 2204 21076 2208
rect 21012 2148 21016 2204
rect 21016 2148 21072 2204
rect 21072 2148 21076 2204
rect 21012 2144 21076 2148
rect 21092 2204 21156 2208
rect 21092 2148 21096 2204
rect 21096 2148 21152 2204
rect 21152 2148 21156 2204
rect 21092 2144 21156 2148
rect 21172 2204 21236 2208
rect 21172 2148 21176 2204
rect 21176 2148 21232 2204
rect 21232 2148 21236 2204
rect 21172 2144 21236 2148
rect 21252 2204 21316 2208
rect 21252 2148 21256 2204
rect 21256 2148 21312 2204
rect 21312 2148 21316 2204
rect 21252 2144 21316 2148
rect 27012 2204 27076 2208
rect 27012 2148 27016 2204
rect 27016 2148 27072 2204
rect 27072 2148 27076 2204
rect 27012 2144 27076 2148
rect 27092 2204 27156 2208
rect 27092 2148 27096 2204
rect 27096 2148 27152 2204
rect 27152 2148 27156 2204
rect 27092 2144 27156 2148
rect 27172 2204 27236 2208
rect 27172 2148 27176 2204
rect 27176 2148 27232 2204
rect 27232 2148 27236 2204
rect 27172 2144 27236 2148
rect 27252 2204 27316 2208
rect 27252 2148 27256 2204
rect 27256 2148 27312 2204
rect 27312 2148 27316 2204
rect 27252 2144 27316 2148
rect 33012 2204 33076 2208
rect 33012 2148 33016 2204
rect 33016 2148 33072 2204
rect 33072 2148 33076 2204
rect 33012 2144 33076 2148
rect 33092 2204 33156 2208
rect 33092 2148 33096 2204
rect 33096 2148 33152 2204
rect 33152 2148 33156 2204
rect 33092 2144 33156 2148
rect 33172 2204 33236 2208
rect 33172 2148 33176 2204
rect 33176 2148 33232 2204
rect 33232 2148 33236 2204
rect 33172 2144 33236 2148
rect 33252 2204 33316 2208
rect 33252 2148 33256 2204
rect 33256 2148 33312 2204
rect 33312 2148 33316 2204
rect 33252 2144 33316 2148
rect 39012 2204 39076 2208
rect 39012 2148 39016 2204
rect 39016 2148 39072 2204
rect 39072 2148 39076 2204
rect 39012 2144 39076 2148
rect 39092 2204 39156 2208
rect 39092 2148 39096 2204
rect 39096 2148 39152 2204
rect 39152 2148 39156 2204
rect 39092 2144 39156 2148
rect 39172 2204 39236 2208
rect 39172 2148 39176 2204
rect 39176 2148 39232 2204
rect 39232 2148 39236 2204
rect 39172 2144 39236 2148
rect 39252 2204 39316 2208
rect 39252 2148 39256 2204
rect 39256 2148 39312 2204
rect 39312 2148 39316 2204
rect 39252 2144 39316 2148
rect 7052 1668 7116 1732
rect 3924 1396 3988 1460
rect 5580 1124 5644 1188
rect 2452 988 2516 1052
rect 6684 852 6748 916
rect 25268 580 25332 644
rect 22140 444 22204 508
<< metal4 >>
rect 1944 8192 2264 11250
rect 2635 10164 2701 10165
rect 2635 10100 2636 10164
rect 2700 10100 2701 10164
rect 2635 10099 2701 10100
rect 1944 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2264 8192
rect 1944 7104 2264 8128
rect 1944 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2264 7104
rect 1944 6016 2264 7040
rect 2451 6356 2517 6357
rect 2451 6292 2452 6356
rect 2516 6292 2517 6356
rect 2451 6291 2517 6292
rect 1944 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2264 6016
rect 1944 4928 2264 5952
rect 1944 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2264 4928
rect 1944 3840 2264 4864
rect 1944 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2264 3840
rect 1944 2752 2264 3776
rect 1944 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2264 2752
rect 1944 0 2264 2688
rect 2454 1053 2514 6291
rect 2638 5949 2698 10099
rect 3004 8736 3324 11250
rect 7787 10028 7853 10029
rect 7787 9964 7788 10028
rect 7852 9964 7853 10028
rect 7787 9963 7853 9964
rect 7603 9348 7669 9349
rect 7603 9284 7604 9348
rect 7668 9284 7669 9348
rect 7603 9283 7669 9284
rect 3004 8672 3012 8736
rect 3076 8672 3092 8736
rect 3156 8672 3172 8736
rect 3236 8672 3252 8736
rect 3316 8672 3324 8736
rect 3004 7648 3324 8672
rect 7051 8532 7117 8533
rect 7051 8468 7052 8532
rect 7116 8468 7117 8532
rect 7051 8467 7117 8468
rect 3004 7584 3012 7648
rect 3076 7584 3092 7648
rect 3156 7584 3172 7648
rect 3236 7584 3252 7648
rect 3316 7584 3324 7648
rect 3004 6560 3324 7584
rect 3923 7036 3989 7037
rect 3923 6972 3924 7036
rect 3988 6972 3989 7036
rect 3923 6971 3989 6972
rect 6683 7036 6749 7037
rect 6683 6972 6684 7036
rect 6748 6972 6749 7036
rect 6683 6971 6749 6972
rect 3004 6496 3012 6560
rect 3076 6496 3092 6560
rect 3156 6496 3172 6560
rect 3236 6496 3252 6560
rect 3316 6496 3324 6560
rect 2635 5948 2701 5949
rect 2635 5884 2636 5948
rect 2700 5884 2701 5948
rect 2635 5883 2701 5884
rect 3004 5472 3324 6496
rect 3004 5408 3012 5472
rect 3076 5408 3092 5472
rect 3156 5408 3172 5472
rect 3236 5408 3252 5472
rect 3316 5408 3324 5472
rect 3004 4384 3324 5408
rect 3004 4320 3012 4384
rect 3076 4320 3092 4384
rect 3156 4320 3172 4384
rect 3236 4320 3252 4384
rect 3316 4320 3324 4384
rect 3004 3296 3324 4320
rect 3004 3232 3012 3296
rect 3076 3232 3092 3296
rect 3156 3232 3172 3296
rect 3236 3232 3252 3296
rect 3316 3232 3324 3296
rect 3004 2208 3324 3232
rect 3004 2144 3012 2208
rect 3076 2144 3092 2208
rect 3156 2144 3172 2208
rect 3236 2144 3252 2208
rect 3316 2144 3324 2208
rect 2451 1052 2517 1053
rect 2451 988 2452 1052
rect 2516 988 2517 1052
rect 2451 987 2517 988
rect 3004 0 3324 2144
rect 3926 1461 3986 6971
rect 5395 6628 5461 6629
rect 5395 6564 5396 6628
rect 5460 6564 5461 6628
rect 5395 6563 5461 6564
rect 5398 3909 5458 6563
rect 5579 5948 5645 5949
rect 5579 5884 5580 5948
rect 5644 5884 5645 5948
rect 5579 5883 5645 5884
rect 5395 3908 5461 3909
rect 5395 3844 5396 3908
rect 5460 3844 5461 3908
rect 5395 3843 5461 3844
rect 3923 1460 3989 1461
rect 3923 1396 3924 1460
rect 3988 1396 3989 1460
rect 3923 1395 3989 1396
rect 5582 1189 5642 5883
rect 5579 1188 5645 1189
rect 5579 1124 5580 1188
rect 5644 1124 5645 1188
rect 5579 1123 5645 1124
rect 6686 917 6746 6971
rect 7054 5405 7114 8467
rect 7051 5404 7117 5405
rect 7051 5340 7052 5404
rect 7116 5340 7117 5404
rect 7051 5339 7117 5340
rect 7051 4180 7117 4181
rect 7051 4116 7052 4180
rect 7116 4116 7117 4180
rect 7051 4115 7117 4116
rect 7054 1733 7114 4115
rect 7606 3773 7666 9283
rect 7790 8261 7850 9963
rect 7787 8260 7853 8261
rect 7787 8196 7788 8260
rect 7852 8196 7853 8260
rect 7787 8195 7853 8196
rect 7944 8192 8264 11250
rect 9004 8736 9324 11250
rect 9627 8804 9693 8805
rect 9627 8740 9628 8804
rect 9692 8740 9693 8804
rect 9627 8739 9693 8740
rect 9004 8672 9012 8736
rect 9076 8672 9092 8736
rect 9156 8672 9172 8736
rect 9236 8672 9252 8736
rect 9316 8672 9324 8736
rect 8523 8260 8589 8261
rect 8523 8196 8524 8260
rect 8588 8196 8589 8260
rect 8523 8195 8589 8196
rect 7944 8128 7952 8192
rect 8016 8128 8032 8192
rect 8096 8128 8112 8192
rect 8176 8128 8192 8192
rect 8256 8128 8264 8192
rect 7944 7104 8264 8128
rect 8526 7173 8586 8195
rect 9004 7648 9324 8672
rect 9004 7584 9012 7648
rect 9076 7584 9092 7648
rect 9156 7584 9172 7648
rect 9236 7584 9252 7648
rect 9316 7584 9324 7648
rect 8707 7308 8773 7309
rect 8707 7244 8708 7308
rect 8772 7244 8773 7308
rect 8707 7243 8773 7244
rect 8523 7172 8589 7173
rect 8523 7108 8524 7172
rect 8588 7108 8589 7172
rect 8523 7107 8589 7108
rect 7944 7040 7952 7104
rect 8016 7040 8032 7104
rect 8096 7040 8112 7104
rect 8176 7040 8192 7104
rect 8256 7040 8264 7104
rect 7944 6016 8264 7040
rect 7944 5952 7952 6016
rect 8016 5952 8032 6016
rect 8096 5952 8112 6016
rect 8176 5952 8192 6016
rect 8256 5952 8264 6016
rect 7944 4928 8264 5952
rect 8523 5540 8589 5541
rect 8523 5476 8524 5540
rect 8588 5476 8589 5540
rect 8523 5475 8589 5476
rect 8526 4997 8586 5475
rect 8710 5405 8770 7243
rect 9004 6560 9324 7584
rect 9004 6496 9012 6560
rect 9076 6496 9092 6560
rect 9156 6496 9172 6560
rect 9236 6496 9252 6560
rect 9316 6496 9324 6560
rect 9004 5472 9324 6496
rect 9004 5408 9012 5472
rect 9076 5408 9092 5472
rect 9156 5408 9172 5472
rect 9236 5408 9252 5472
rect 9316 5408 9324 5472
rect 8707 5404 8773 5405
rect 8707 5340 8708 5404
rect 8772 5340 8773 5404
rect 8707 5339 8773 5340
rect 8523 4996 8589 4997
rect 8523 4932 8524 4996
rect 8588 4932 8589 4996
rect 8523 4931 8589 4932
rect 7944 4864 7952 4928
rect 8016 4864 8032 4928
rect 8096 4864 8112 4928
rect 8176 4864 8192 4928
rect 8256 4864 8264 4928
rect 7944 3840 8264 4864
rect 7944 3776 7952 3840
rect 8016 3776 8032 3840
rect 8096 3776 8112 3840
rect 8176 3776 8192 3840
rect 8256 3776 8264 3840
rect 7603 3772 7669 3773
rect 7603 3708 7604 3772
rect 7668 3708 7669 3772
rect 7603 3707 7669 3708
rect 7944 2752 8264 3776
rect 7944 2688 7952 2752
rect 8016 2688 8032 2752
rect 8096 2688 8112 2752
rect 8176 2688 8192 2752
rect 8256 2688 8264 2752
rect 7051 1732 7117 1733
rect 7051 1668 7052 1732
rect 7116 1668 7117 1732
rect 7051 1667 7117 1668
rect 6683 916 6749 917
rect 6683 852 6684 916
rect 6748 852 6749 916
rect 6683 851 6749 852
rect 7944 0 8264 2688
rect 9004 4384 9324 5408
rect 9004 4320 9012 4384
rect 9076 4320 9092 4384
rect 9156 4320 9172 4384
rect 9236 4320 9252 4384
rect 9316 4320 9324 4384
rect 9004 3296 9324 4320
rect 9630 3637 9690 8739
rect 13944 8192 14264 11250
rect 13944 8128 13952 8192
rect 14016 8128 14032 8192
rect 14096 8128 14112 8192
rect 14176 8128 14192 8192
rect 14256 8128 14264 8192
rect 10915 7852 10981 7853
rect 10915 7788 10916 7852
rect 10980 7788 10981 7852
rect 10915 7787 10981 7788
rect 10363 7580 10429 7581
rect 10363 7516 10364 7580
rect 10428 7516 10429 7580
rect 10363 7515 10429 7516
rect 9811 5268 9877 5269
rect 9811 5204 9812 5268
rect 9876 5204 9877 5268
rect 9811 5203 9877 5204
rect 9814 3909 9874 5203
rect 9811 3908 9877 3909
rect 9811 3844 9812 3908
rect 9876 3844 9877 3908
rect 9811 3843 9877 3844
rect 9627 3636 9693 3637
rect 9627 3572 9628 3636
rect 9692 3572 9693 3636
rect 9627 3571 9693 3572
rect 9004 3232 9012 3296
rect 9076 3232 9092 3296
rect 9156 3232 9172 3296
rect 9236 3232 9252 3296
rect 9316 3232 9324 3296
rect 9004 2208 9324 3232
rect 10366 2277 10426 7515
rect 10918 4317 10978 7787
rect 13944 7104 14264 8128
rect 15004 8736 15324 11250
rect 15515 9484 15581 9485
rect 15515 9420 15516 9484
rect 15580 9420 15581 9484
rect 15515 9419 15581 9420
rect 15004 8672 15012 8736
rect 15076 8672 15092 8736
rect 15156 8672 15172 8736
rect 15236 8672 15252 8736
rect 15316 8672 15324 8736
rect 15004 7648 15324 8672
rect 15004 7584 15012 7648
rect 15076 7584 15092 7648
rect 15156 7584 15172 7648
rect 15236 7584 15252 7648
rect 15316 7584 15324 7648
rect 14779 7172 14845 7173
rect 14779 7108 14780 7172
rect 14844 7108 14845 7172
rect 14779 7107 14845 7108
rect 13944 7040 13952 7104
rect 14016 7040 14032 7104
rect 14096 7040 14112 7104
rect 14176 7040 14192 7104
rect 14256 7040 14264 7104
rect 13944 6016 14264 7040
rect 13944 5952 13952 6016
rect 14016 5952 14032 6016
rect 14096 5952 14112 6016
rect 14176 5952 14192 6016
rect 14256 5952 14264 6016
rect 13944 4928 14264 5952
rect 14595 5948 14661 5949
rect 14595 5884 14596 5948
rect 14660 5884 14661 5948
rect 14595 5883 14661 5884
rect 13944 4864 13952 4928
rect 14016 4864 14032 4928
rect 14096 4864 14112 4928
rect 14176 4864 14192 4928
rect 14256 4864 14264 4928
rect 10915 4316 10981 4317
rect 10915 4252 10916 4316
rect 10980 4252 10981 4316
rect 10915 4251 10981 4252
rect 13944 3840 14264 4864
rect 13944 3776 13952 3840
rect 14016 3776 14032 3840
rect 14096 3776 14112 3840
rect 14176 3776 14192 3840
rect 14256 3776 14264 3840
rect 13944 2752 14264 3776
rect 13944 2688 13952 2752
rect 14016 2688 14032 2752
rect 14096 2688 14112 2752
rect 14176 2688 14192 2752
rect 14256 2688 14264 2752
rect 10363 2276 10429 2277
rect 10363 2212 10364 2276
rect 10428 2212 10429 2276
rect 10363 2211 10429 2212
rect 9004 2144 9012 2208
rect 9076 2144 9092 2208
rect 9156 2144 9172 2208
rect 9236 2144 9252 2208
rect 9316 2144 9324 2208
rect 9004 0 9324 2144
rect 13944 0 14264 2688
rect 14598 2549 14658 5883
rect 14782 4453 14842 7107
rect 15004 6560 15324 7584
rect 15004 6496 15012 6560
rect 15076 6496 15092 6560
rect 15156 6496 15172 6560
rect 15236 6496 15252 6560
rect 15316 6496 15324 6560
rect 15004 5472 15324 6496
rect 15004 5408 15012 5472
rect 15076 5408 15092 5472
rect 15156 5408 15172 5472
rect 15236 5408 15252 5472
rect 15316 5408 15324 5472
rect 14779 4452 14845 4453
rect 14779 4388 14780 4452
rect 14844 4388 14845 4452
rect 14779 4387 14845 4388
rect 15004 4384 15324 5408
rect 15004 4320 15012 4384
rect 15076 4320 15092 4384
rect 15156 4320 15172 4384
rect 15236 4320 15252 4384
rect 15316 4320 15324 4384
rect 15004 3296 15324 4320
rect 15518 3773 15578 9419
rect 18643 8668 18709 8669
rect 18643 8604 18644 8668
rect 18708 8604 18709 8668
rect 18643 8603 18709 8604
rect 16803 8532 16869 8533
rect 16803 8468 16804 8532
rect 16868 8468 16869 8532
rect 16803 8467 16869 8468
rect 16251 7172 16317 7173
rect 16251 7108 16252 7172
rect 16316 7108 16317 7172
rect 16251 7107 16317 7108
rect 15883 7036 15949 7037
rect 15883 6972 15884 7036
rect 15948 6972 15949 7036
rect 15883 6971 15949 6972
rect 15886 3909 15946 6971
rect 16067 6492 16133 6493
rect 16067 6428 16068 6492
rect 16132 6428 16133 6492
rect 16067 6427 16133 6428
rect 16070 4181 16130 6427
rect 16254 6085 16314 7107
rect 16251 6084 16317 6085
rect 16251 6020 16252 6084
rect 16316 6020 16317 6084
rect 16251 6019 16317 6020
rect 16067 4180 16133 4181
rect 16067 4116 16068 4180
rect 16132 4116 16133 4180
rect 16067 4115 16133 4116
rect 15883 3908 15949 3909
rect 15883 3844 15884 3908
rect 15948 3844 15949 3908
rect 15883 3843 15949 3844
rect 16806 3773 16866 8467
rect 17907 8396 17973 8397
rect 17907 8332 17908 8396
rect 17972 8332 17973 8396
rect 17907 8331 17973 8332
rect 15515 3772 15581 3773
rect 15515 3708 15516 3772
rect 15580 3708 15581 3772
rect 15515 3707 15581 3708
rect 16803 3772 16869 3773
rect 16803 3708 16804 3772
rect 16868 3708 16869 3772
rect 16803 3707 16869 3708
rect 17910 3501 17970 8331
rect 18459 8124 18525 8125
rect 18459 8060 18460 8124
rect 18524 8060 18525 8124
rect 18459 8059 18525 8060
rect 18275 6356 18341 6357
rect 18275 6292 18276 6356
rect 18340 6292 18341 6356
rect 18275 6291 18341 6292
rect 18278 6085 18338 6291
rect 18275 6084 18341 6085
rect 18275 6020 18276 6084
rect 18340 6020 18341 6084
rect 18275 6019 18341 6020
rect 18462 5269 18522 8059
rect 18646 7037 18706 8603
rect 19944 8192 20264 11250
rect 19944 8128 19952 8192
rect 20016 8128 20032 8192
rect 20096 8128 20112 8192
rect 20176 8128 20192 8192
rect 20256 8128 20264 8192
rect 19011 8124 19077 8125
rect 19011 8060 19012 8124
rect 19076 8060 19077 8124
rect 19011 8059 19077 8060
rect 18643 7036 18709 7037
rect 18643 6972 18644 7036
rect 18708 6972 18709 7036
rect 18643 6971 18709 6972
rect 19014 6493 19074 8059
rect 19944 7104 20264 8128
rect 19944 7040 19952 7104
rect 20016 7040 20032 7104
rect 20096 7040 20112 7104
rect 20176 7040 20192 7104
rect 20256 7040 20264 7104
rect 19011 6492 19077 6493
rect 19011 6428 19012 6492
rect 19076 6428 19077 6492
rect 19011 6427 19077 6428
rect 19944 6016 20264 7040
rect 19944 5952 19952 6016
rect 20016 5952 20032 6016
rect 20096 5952 20112 6016
rect 20176 5952 20192 6016
rect 20256 5952 20264 6016
rect 18459 5268 18525 5269
rect 18459 5204 18460 5268
rect 18524 5204 18525 5268
rect 18459 5203 18525 5204
rect 19944 4928 20264 5952
rect 19944 4864 19952 4928
rect 20016 4864 20032 4928
rect 20096 4864 20112 4928
rect 20176 4864 20192 4928
rect 20256 4864 20264 4928
rect 19944 3840 20264 4864
rect 19944 3776 19952 3840
rect 20016 3776 20032 3840
rect 20096 3776 20112 3840
rect 20176 3776 20192 3840
rect 20256 3776 20264 3840
rect 17907 3500 17973 3501
rect 17907 3436 17908 3500
rect 17972 3436 17973 3500
rect 17907 3435 17973 3436
rect 15004 3232 15012 3296
rect 15076 3232 15092 3296
rect 15156 3232 15172 3296
rect 15236 3232 15252 3296
rect 15316 3232 15324 3296
rect 14595 2548 14661 2549
rect 14595 2484 14596 2548
rect 14660 2484 14661 2548
rect 14595 2483 14661 2484
rect 15004 2208 15324 3232
rect 15004 2144 15012 2208
rect 15076 2144 15092 2208
rect 15156 2144 15172 2208
rect 15236 2144 15252 2208
rect 15316 2144 15324 2208
rect 15004 0 15324 2144
rect 19944 2752 20264 3776
rect 19944 2688 19952 2752
rect 20016 2688 20032 2752
rect 20096 2688 20112 2752
rect 20176 2688 20192 2752
rect 20256 2688 20264 2752
rect 19944 0 20264 2688
rect 21004 8736 21324 11250
rect 24899 10300 24965 10301
rect 24899 10236 24900 10300
rect 24964 10236 24965 10300
rect 24899 10235 24965 10236
rect 23427 10028 23493 10029
rect 23427 9964 23428 10028
rect 23492 9964 23493 10028
rect 23427 9963 23493 9964
rect 21004 8672 21012 8736
rect 21076 8672 21092 8736
rect 21156 8672 21172 8736
rect 21236 8672 21252 8736
rect 21316 8672 21324 8736
rect 21004 7648 21324 8672
rect 21004 7584 21012 7648
rect 21076 7584 21092 7648
rect 21156 7584 21172 7648
rect 21236 7584 21252 7648
rect 21316 7584 21324 7648
rect 21004 6560 21324 7584
rect 23430 6901 23490 9963
rect 24163 9212 24229 9213
rect 24163 9148 24164 9212
rect 24228 9148 24229 9212
rect 24163 9147 24229 9148
rect 23427 6900 23493 6901
rect 23427 6836 23428 6900
rect 23492 6836 23493 6900
rect 23427 6835 23493 6836
rect 21004 6496 21012 6560
rect 21076 6496 21092 6560
rect 21156 6496 21172 6560
rect 21236 6496 21252 6560
rect 21316 6496 21324 6560
rect 21004 5472 21324 6496
rect 22139 5676 22205 5677
rect 22139 5612 22140 5676
rect 22204 5612 22205 5676
rect 22139 5611 22205 5612
rect 21004 5408 21012 5472
rect 21076 5408 21092 5472
rect 21156 5408 21172 5472
rect 21236 5408 21252 5472
rect 21316 5408 21324 5472
rect 21004 4384 21324 5408
rect 21004 4320 21012 4384
rect 21076 4320 21092 4384
rect 21156 4320 21172 4384
rect 21236 4320 21252 4384
rect 21316 4320 21324 4384
rect 21004 3296 21324 4320
rect 21004 3232 21012 3296
rect 21076 3232 21092 3296
rect 21156 3232 21172 3296
rect 21236 3232 21252 3296
rect 21316 3232 21324 3296
rect 21004 2208 21324 3232
rect 21004 2144 21012 2208
rect 21076 2144 21092 2208
rect 21156 2144 21172 2208
rect 21236 2144 21252 2208
rect 21316 2144 21324 2208
rect 21004 0 21324 2144
rect 22142 509 22202 5611
rect 24166 3229 24226 9147
rect 24902 6493 24962 10235
rect 25267 8532 25333 8533
rect 25267 8468 25268 8532
rect 25332 8468 25333 8532
rect 25267 8467 25333 8468
rect 24899 6492 24965 6493
rect 24899 6428 24900 6492
rect 24964 6428 24965 6492
rect 24899 6427 24965 6428
rect 24163 3228 24229 3229
rect 24163 3164 24164 3228
rect 24228 3164 24229 3228
rect 24163 3163 24229 3164
rect 25270 645 25330 8467
rect 25451 8260 25517 8261
rect 25451 8196 25452 8260
rect 25516 8196 25517 8260
rect 25451 8195 25517 8196
rect 25454 3093 25514 8195
rect 25944 8192 26264 11250
rect 26739 10436 26805 10437
rect 26739 10372 26740 10436
rect 26804 10372 26805 10436
rect 26739 10371 26805 10372
rect 26555 8532 26621 8533
rect 26555 8468 26556 8532
rect 26620 8468 26621 8532
rect 26555 8467 26621 8468
rect 25944 8128 25952 8192
rect 26016 8128 26032 8192
rect 26096 8128 26112 8192
rect 26176 8128 26192 8192
rect 26256 8128 26264 8192
rect 25635 8124 25701 8125
rect 25635 8060 25636 8124
rect 25700 8060 25701 8124
rect 25635 8059 25701 8060
rect 25638 6901 25698 8059
rect 25944 7104 26264 8128
rect 26371 8124 26437 8125
rect 26371 8060 26372 8124
rect 26436 8060 26437 8124
rect 26371 8059 26437 8060
rect 25944 7040 25952 7104
rect 26016 7040 26032 7104
rect 26096 7040 26112 7104
rect 26176 7040 26192 7104
rect 26256 7040 26264 7104
rect 25635 6900 25701 6901
rect 25635 6836 25636 6900
rect 25700 6836 25701 6900
rect 25635 6835 25701 6836
rect 25944 6016 26264 7040
rect 25944 5952 25952 6016
rect 26016 5952 26032 6016
rect 26096 5952 26112 6016
rect 26176 5952 26192 6016
rect 26256 5952 26264 6016
rect 25944 4928 26264 5952
rect 25944 4864 25952 4928
rect 26016 4864 26032 4928
rect 26096 4864 26112 4928
rect 26176 4864 26192 4928
rect 26256 4864 26264 4928
rect 25944 3840 26264 4864
rect 25944 3776 25952 3840
rect 26016 3776 26032 3840
rect 26096 3776 26112 3840
rect 26176 3776 26192 3840
rect 26256 3776 26264 3840
rect 25451 3092 25517 3093
rect 25451 3028 25452 3092
rect 25516 3028 25517 3092
rect 25451 3027 25517 3028
rect 25944 2752 26264 3776
rect 26374 2957 26434 8059
rect 26558 2957 26618 8467
rect 26742 7037 26802 10371
rect 27004 8736 27324 11250
rect 27004 8672 27012 8736
rect 27076 8672 27092 8736
rect 27156 8672 27172 8736
rect 27236 8672 27252 8736
rect 27316 8672 27324 8736
rect 27004 7648 27324 8672
rect 28027 8668 28093 8669
rect 28027 8604 28028 8668
rect 28092 8604 28093 8668
rect 28027 8603 28093 8604
rect 27004 7584 27012 7648
rect 27076 7584 27092 7648
rect 27156 7584 27172 7648
rect 27236 7584 27252 7648
rect 27316 7584 27324 7648
rect 26739 7036 26805 7037
rect 26739 6972 26740 7036
rect 26804 6972 26805 7036
rect 26739 6971 26805 6972
rect 27004 6560 27324 7584
rect 27004 6496 27012 6560
rect 27076 6496 27092 6560
rect 27156 6496 27172 6560
rect 27236 6496 27252 6560
rect 27316 6496 27324 6560
rect 27004 5472 27324 6496
rect 28030 6357 28090 8603
rect 31944 8192 32264 11250
rect 32443 9484 32509 9485
rect 32443 9420 32444 9484
rect 32508 9420 32509 9484
rect 32443 9419 32509 9420
rect 31944 8128 31952 8192
rect 32016 8128 32032 8192
rect 32096 8128 32112 8192
rect 32176 8128 32192 8192
rect 32256 8128 32264 8192
rect 30603 8124 30669 8125
rect 30603 8060 30604 8124
rect 30668 8060 30669 8124
rect 30603 8059 30669 8060
rect 28027 6356 28093 6357
rect 28027 6292 28028 6356
rect 28092 6292 28093 6356
rect 28027 6291 28093 6292
rect 27004 5408 27012 5472
rect 27076 5408 27092 5472
rect 27156 5408 27172 5472
rect 27236 5408 27252 5472
rect 27316 5408 27324 5472
rect 27004 4384 27324 5408
rect 30606 4861 30666 8059
rect 31339 7580 31405 7581
rect 31339 7516 31340 7580
rect 31404 7516 31405 7580
rect 31339 7515 31405 7516
rect 31342 6493 31402 7515
rect 31944 7104 32264 8128
rect 31944 7040 31952 7104
rect 32016 7040 32032 7104
rect 32096 7040 32112 7104
rect 32176 7040 32192 7104
rect 32256 7040 32264 7104
rect 31339 6492 31405 6493
rect 31339 6428 31340 6492
rect 31404 6428 31405 6492
rect 31339 6427 31405 6428
rect 31944 6016 32264 7040
rect 32446 6221 32506 9419
rect 32811 9076 32877 9077
rect 32811 9012 32812 9076
rect 32876 9012 32877 9076
rect 32811 9011 32877 9012
rect 32627 8124 32693 8125
rect 32627 8060 32628 8124
rect 32692 8060 32693 8124
rect 32627 8059 32693 8060
rect 32630 7581 32690 8059
rect 32627 7580 32693 7581
rect 32627 7516 32628 7580
rect 32692 7516 32693 7580
rect 32627 7515 32693 7516
rect 32443 6220 32509 6221
rect 32443 6156 32444 6220
rect 32508 6156 32509 6220
rect 32443 6155 32509 6156
rect 31944 5952 31952 6016
rect 32016 5952 32032 6016
rect 32096 5952 32112 6016
rect 32176 5952 32192 6016
rect 32256 5952 32264 6016
rect 31944 4928 32264 5952
rect 31944 4864 31952 4928
rect 32016 4864 32032 4928
rect 32096 4864 32112 4928
rect 32176 4864 32192 4928
rect 32256 4864 32264 4928
rect 30603 4860 30669 4861
rect 30603 4796 30604 4860
rect 30668 4796 30669 4860
rect 30603 4795 30669 4796
rect 27004 4320 27012 4384
rect 27076 4320 27092 4384
rect 27156 4320 27172 4384
rect 27236 4320 27252 4384
rect 27316 4320 27324 4384
rect 27004 3296 27324 4320
rect 27004 3232 27012 3296
rect 27076 3232 27092 3296
rect 27156 3232 27172 3296
rect 27236 3232 27252 3296
rect 27316 3232 27324 3296
rect 26371 2956 26437 2957
rect 26371 2892 26372 2956
rect 26436 2892 26437 2956
rect 26371 2891 26437 2892
rect 26555 2956 26621 2957
rect 26555 2892 26556 2956
rect 26620 2892 26621 2956
rect 26555 2891 26621 2892
rect 25944 2688 25952 2752
rect 26016 2688 26032 2752
rect 26096 2688 26112 2752
rect 26176 2688 26192 2752
rect 26256 2688 26264 2752
rect 25267 644 25333 645
rect 25267 580 25268 644
rect 25332 580 25333 644
rect 25267 579 25333 580
rect 22139 508 22205 509
rect 22139 444 22140 508
rect 22204 444 22205 508
rect 22139 443 22205 444
rect 25944 0 26264 2688
rect 27004 2208 27324 3232
rect 27004 2144 27012 2208
rect 27076 2144 27092 2208
rect 27156 2144 27172 2208
rect 27236 2144 27252 2208
rect 27316 2144 27324 2208
rect 27004 0 27324 2144
rect 31944 3840 32264 4864
rect 32814 4181 32874 9011
rect 33004 8736 33324 11250
rect 33731 9892 33797 9893
rect 33731 9828 33732 9892
rect 33796 9828 33797 9892
rect 33731 9827 33797 9828
rect 33004 8672 33012 8736
rect 33076 8672 33092 8736
rect 33156 8672 33172 8736
rect 33236 8672 33252 8736
rect 33316 8672 33324 8736
rect 33004 7648 33324 8672
rect 33004 7584 33012 7648
rect 33076 7584 33092 7648
rect 33156 7584 33172 7648
rect 33236 7584 33252 7648
rect 33316 7584 33324 7648
rect 33004 6560 33324 7584
rect 33004 6496 33012 6560
rect 33076 6496 33092 6560
rect 33156 6496 33172 6560
rect 33236 6496 33252 6560
rect 33316 6496 33324 6560
rect 33004 5472 33324 6496
rect 33734 5949 33794 9827
rect 37944 8192 38264 11250
rect 37944 8128 37952 8192
rect 38016 8128 38032 8192
rect 38096 8128 38112 8192
rect 38176 8128 38192 8192
rect 38256 8128 38264 8192
rect 37944 7104 38264 8128
rect 37944 7040 37952 7104
rect 38016 7040 38032 7104
rect 38096 7040 38112 7104
rect 38176 7040 38192 7104
rect 38256 7040 38264 7104
rect 37944 6016 38264 7040
rect 37944 5952 37952 6016
rect 38016 5952 38032 6016
rect 38096 5952 38112 6016
rect 38176 5952 38192 6016
rect 38256 5952 38264 6016
rect 33731 5948 33797 5949
rect 33731 5884 33732 5948
rect 33796 5884 33797 5948
rect 33731 5883 33797 5884
rect 37779 5676 37845 5677
rect 37779 5612 37780 5676
rect 37844 5612 37845 5676
rect 37779 5611 37845 5612
rect 33004 5408 33012 5472
rect 33076 5408 33092 5472
rect 33156 5408 33172 5472
rect 33236 5408 33252 5472
rect 33316 5408 33324 5472
rect 33004 4384 33324 5408
rect 33004 4320 33012 4384
rect 33076 4320 33092 4384
rect 33156 4320 33172 4384
rect 33236 4320 33252 4384
rect 33316 4320 33324 4384
rect 32811 4180 32877 4181
rect 32811 4116 32812 4180
rect 32876 4116 32877 4180
rect 32811 4115 32877 4116
rect 31944 3776 31952 3840
rect 32016 3776 32032 3840
rect 32096 3776 32112 3840
rect 32176 3776 32192 3840
rect 32256 3776 32264 3840
rect 31944 2752 32264 3776
rect 31944 2688 31952 2752
rect 32016 2688 32032 2752
rect 32096 2688 32112 2752
rect 32176 2688 32192 2752
rect 32256 2688 32264 2752
rect 31944 0 32264 2688
rect 33004 3296 33324 4320
rect 33004 3232 33012 3296
rect 33076 3232 33092 3296
rect 33156 3232 33172 3296
rect 33236 3232 33252 3296
rect 33316 3232 33324 3296
rect 33004 2208 33324 3232
rect 37782 2549 37842 5611
rect 37944 4928 38264 5952
rect 37944 4864 37952 4928
rect 38016 4864 38032 4928
rect 38096 4864 38112 4928
rect 38176 4864 38192 4928
rect 38256 4864 38264 4928
rect 37944 3840 38264 4864
rect 37944 3776 37952 3840
rect 38016 3776 38032 3840
rect 38096 3776 38112 3840
rect 38176 3776 38192 3840
rect 38256 3776 38264 3840
rect 37944 2752 38264 3776
rect 37944 2688 37952 2752
rect 38016 2688 38032 2752
rect 38096 2688 38112 2752
rect 38176 2688 38192 2752
rect 38256 2688 38264 2752
rect 37779 2548 37845 2549
rect 37779 2484 37780 2548
rect 37844 2484 37845 2548
rect 37779 2483 37845 2484
rect 33004 2144 33012 2208
rect 33076 2144 33092 2208
rect 33156 2144 33172 2208
rect 33236 2144 33252 2208
rect 33316 2144 33324 2208
rect 33004 0 33324 2144
rect 37944 0 38264 2688
rect 39004 8736 39324 11250
rect 39004 8672 39012 8736
rect 39076 8672 39092 8736
rect 39156 8672 39172 8736
rect 39236 8672 39252 8736
rect 39316 8672 39324 8736
rect 39004 7648 39324 8672
rect 39004 7584 39012 7648
rect 39076 7584 39092 7648
rect 39156 7584 39172 7648
rect 39236 7584 39252 7648
rect 39316 7584 39324 7648
rect 39004 6560 39324 7584
rect 39004 6496 39012 6560
rect 39076 6496 39092 6560
rect 39156 6496 39172 6560
rect 39236 6496 39252 6560
rect 39316 6496 39324 6560
rect 39004 5472 39324 6496
rect 39004 5408 39012 5472
rect 39076 5408 39092 5472
rect 39156 5408 39172 5472
rect 39236 5408 39252 5472
rect 39316 5408 39324 5472
rect 39004 4384 39324 5408
rect 39004 4320 39012 4384
rect 39076 4320 39092 4384
rect 39156 4320 39172 4384
rect 39236 4320 39252 4384
rect 39316 4320 39324 4384
rect 39004 3296 39324 4320
rect 39004 3232 39012 3296
rect 39076 3232 39092 3296
rect 39156 3232 39172 3296
rect 39236 3232 39252 3296
rect 39316 3232 39324 3296
rect 39004 2208 39324 3232
rect 39004 2144 39012 2208
rect 39076 2144 39092 2208
rect 39156 2144 39172 2208
rect 39236 2144 39252 2208
rect 39316 2144 39324 2208
rect 39004 0 39324 2144
use sky130_fd_sc_hd__inv_2  _081_
timestamp -3599
transform 1 0 17020 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  _082_
timestamp -3599
transform -1 0 18952 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _083_
timestamp -3599
transform -1 0 22080 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _084_
timestamp -3599
transform -1 0 13616 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _085_
timestamp -3599
transform 1 0 30084 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _086_
timestamp -3599
transform 1 0 6348 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _087_
timestamp -3599
transform 1 0 3772 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _088_
timestamp -3599
transform -1 0 14444 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _089_
timestamp -3599
transform 1 0 23092 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _090_
timestamp -3599
transform -1 0 18584 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _091_
timestamp -3599
transform 1 0 4876 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _092_
timestamp -3599
transform 1 0 33396 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _093_
timestamp -3599
transform 1 0 32936 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _094_
timestamp -3599
transform 1 0 34500 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _095_
timestamp -3599
transform 1 0 36064 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _096_
timestamp -3599
transform 1 0 35972 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _097_
timestamp -3599
transform 1 0 32476 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _098_
timestamp -3599
transform -1 0 21620 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _099_
timestamp -3599
transform -1 0 25208 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _100_
timestamp -3599
transform 1 0 8924 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _101_
timestamp -3599
transform -1 0 17572 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _102_
timestamp -3599
transform 1 0 27140 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _103_
timestamp -3599
transform -1 0 23092 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _104_
timestamp -3599
transform 1 0 24380 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _105_
timestamp -3599
transform 1 0 18492 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _106_
timestamp -3599
transform 1 0 27600 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _107_
timestamp -3599
transform -1 0 18124 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _108_
timestamp -3599
transform -1 0 5704 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _109_
timestamp -3599
transform 1 0 14444 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _110_
timestamp -3599
transform 1 0 11500 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _111_
timestamp -3599
transform 1 0 4876 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _112_
timestamp -3599
transform 1 0 3864 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _113_
timestamp -3599
transform 1 0 13156 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _114_
timestamp -3599
transform 1 0 27232 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _115_
timestamp -3599
transform 1 0 20884 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _116_
timestamp -3599
transform -1 0 6716 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _117_
timestamp -3599
transform 1 0 17572 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _118_
timestamp -3599
transform 1 0 21804 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__nand2b_1  _119_
timestamp -3599
transform -1 0 21252 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _120_
timestamp -3599
transform 1 0 23276 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _121_
timestamp -3599
transform 1 0 23552 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _122_
timestamp -3599
transform 1 0 21252 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__nor2_1  _123_
timestamp -3599
transform -1 0 23000 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _124_
timestamp -3599
transform -1 0 23552 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _125_
timestamp -3599
transform -1 0 25576 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _126_
timestamp -3599
transform -1 0 28980 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _127_
timestamp -3599
transform -1 0 26404 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__a21bo_1  _128_
timestamp -3599
transform -1 0 29900 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__mux4_1  _129_
timestamp -3599
transform 1 0 27324 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__o22a_1  _130_
timestamp -3599
transform 1 0 28152 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _131_
timestamp -3599
transform -1 0 24288 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _132_
timestamp -3599
transform -1 0 11408 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _133_
timestamp -3599
transform 1 0 10304 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _134_
timestamp -3599
transform 1 0 14444 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_1  _135_
timestamp -3599
transform 1 0 18124 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _136_
timestamp -3599
transform 1 0 16652 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _137_
timestamp -3599
transform 1 0 30452 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _138_
timestamp -3599
transform 1 0 29440 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _139_
timestamp -3599
transform 1 0 28796 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _140_
timestamp -3599
transform -1 0 31740 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _141_
timestamp -3599
transform -1 0 31096 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _142_
timestamp -3599
transform 1 0 22172 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _143_
timestamp -3599
transform -1 0 23828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _144_
timestamp -3599
transform -1 0 23276 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o211ai_1  _145_
timestamp -3599
transform -1 0 19136 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _146_
timestamp -3599
transform -1 0 16560 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _147_
timestamp -3599
transform 1 0 17388 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _148_
timestamp -3599
transform -1 0 20424 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _149_
timestamp -3599
transform -1 0 25668 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _150_
timestamp -3599
transform -1 0 25852 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _151_
timestamp -3599
transform 1 0 24380 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _152_
timestamp -3599
transform 1 0 24748 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _153_
timestamp -3599
transform -1 0 23736 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _154_
timestamp -3599
transform 1 0 32108 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _155_
timestamp -3599
transform -1 0 34592 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _156_
timestamp -3599
transform -1 0 7176 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _157_
timestamp -3599
transform -1 0 18584 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _158_
timestamp -3599
transform -1 0 30360 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _159_
timestamp -3599
transform 1 0 6532 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _160_
timestamp -3599
transform 1 0 2760 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _161_
timestamp -3599
transform -1 0 9752 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _162_
timestamp -3599
transform -1 0 11408 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _163_
timestamp -3599
transform 1 0 6900 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _164_
timestamp -3599
transform 1 0 4048 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _165_
timestamp -3599
transform -1 0 15824 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _166_
timestamp -3599
transform 1 0 26956 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _167_
timestamp -3599
transform 1 0 26956 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _168_
timestamp -3599
transform 1 0 21804 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _169_
timestamp -3599
transform 1 0 20424 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _170_
timestamp -3599
transform -1 0 14352 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _171_
timestamp -3599
transform -1 0 15916 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _172_
timestamp -3599
transform -1 0 19136 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _173_
timestamp -3599
transform 1 0 13708 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _174_
timestamp -3599
transform 1 0 13064 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _175_
timestamp -3599
transform 1 0 18584 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _176_
timestamp -3599
transform 1 0 15180 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _177_
timestamp -3599
transform -1 0 17020 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _178_
timestamp -3599
transform -1 0 16284 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _179_
timestamp -3599
transform -1 0 17112 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _180_
timestamp -3599
transform 1 0 15548 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _181_
timestamp -3599
transform 1 0 8740 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _182_
timestamp -3599
transform -1 0 9476 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _183_
timestamp -3599
transform 1 0 8096 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _184_
timestamp -3599
transform -1 0 11776 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _185_
timestamp -3599
transform 1 0 10948 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _186_
timestamp -3599
transform -1 0 12144 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _187_
timestamp -3599
transform 1 0 1932 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _188_
timestamp -3599
transform 1 0 9016 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _189_
timestamp -3599
transform -1 0 11132 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _190_
timestamp -3599
transform 1 0 1656 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _191_
timestamp -3599
transform 1 0 7820 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _192_
timestamp -3599
transform -1 0 8832 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _193_
timestamp -3599
transform 1 0 8464 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _194_
timestamp -3599
transform 1 0 7820 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _195_
timestamp -3599
transform 1 0 8280 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _196_
timestamp -3599
transform 1 0 9016 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _197_
timestamp -3599
transform 1 0 8372 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _198_
timestamp -3599
transform 1 0 9936 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _199_
timestamp -3599
transform 1 0 9292 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _200_
timestamp -3599
transform 1 0 11500 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _201_
timestamp -3599
transform -1 0 12236 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _202_
timestamp -3599
transform 1 0 10304 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _203_
timestamp -3599
transform -1 0 14536 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _204_
timestamp -3599
transform -1 0 12696 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _205_
timestamp -3599
transform 1 0 10488 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _206_
timestamp -3599
transform -1 0 15088 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _207_
timestamp -3599
transform -1 0 32660 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a21boi_1  _208_
timestamp -3599
transform 1 0 31096 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _209_
timestamp -3599
transform -1 0 33580 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _210_
timestamp -3599
transform 1 0 29532 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _211_
timestamp -3599
transform 1 0 30084 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _212_
timestamp -3599
transform -1 0 29992 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _213_
timestamp -3599
transform -1 0 29164 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _214_
timestamp -3599
transform -1 0 30084 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _215_
timestamp -3599
transform -1 0 28704 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  _216_
timestamp -3599
transform 1 0 19228 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _217_
timestamp -3599
transform 1 0 18768 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _218_
timestamp -3599
transform -1 0 18124 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _219_
timestamp -3599
transform -1 0 24196 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _220_
timestamp -3599
transform 1 0 20240 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _221_
timestamp -3599
transform 1 0 17112 0 -1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _222_
timestamp -3599
transform -1 0 24104 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dlxtp_1  _223_
timestamp -3599
transform 1 0 30176 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _224_
timestamp -3599
transform 1 0 30360 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _225_
timestamp -3599
transform 1 0 28796 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _226_
timestamp -3599
transform 1 0 27692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _227_
timestamp -3599
transform -1 0 19044 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _228_
timestamp -3599
transform 1 0 15088 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _229_
timestamp -3599
transform 1 0 3864 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _230_
timestamp -3599
transform 1 0 4416 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _231_
timestamp -3599
transform 1 0 20516 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _232_
timestamp -3599
transform 1 0 19320 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _233_
timestamp -3599
transform 1 0 25760 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _234_
timestamp -3599
transform 1 0 26772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _235_
timestamp -3599
transform 1 0 11776 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _236_
timestamp -3599
transform 1 0 3312 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _237_
timestamp -3599
transform -1 0 6256 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _238_
timestamp -3599
transform 1 0 10304 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _239_
timestamp -3599
transform 1 0 8648 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _240_
timestamp -3599
transform 1 0 3312 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _241_
timestamp -3599
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _242_
timestamp -3599
transform 1 0 27876 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _243_
timestamp -3599
transform 1 0 17296 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _244_
timestamp -3599
transform 1 0 6716 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _245_
timestamp -3599
transform -1 0 26864 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _246_
timestamp -3599
transform 1 0 26220 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _247_
timestamp -3599
transform -1 0 18308 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _248_
timestamp -3599
transform 1 0 7636 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _249_
timestamp -3599
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _250_
timestamp -3599
transform 1 0 20424 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _251_
timestamp -3599
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _252_
timestamp -3599
transform 1 0 34868 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _253_
timestamp -3599
transform 1 0 34960 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _254_
timestamp -3599
transform 1 0 33396 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _255_
timestamp -3599
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _256_
timestamp -3599
transform 1 0 32292 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _257_
timestamp -3599
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _258_
timestamp -3599
transform 1 0 17388 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _259_
timestamp -3599
transform 1 0 21988 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _260_
timestamp -3599
transform 1 0 12880 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _261_
timestamp -3599
transform 1 0 2760 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _262_
timestamp -3599
transform 1 0 4968 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _263_
timestamp -3599
transform 1 0 19504 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _264_
timestamp -3599
transform 1 0 19412 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _265_
timestamp -3599
transform 1 0 25760 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _266_
timestamp -3599
transform -1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _267_
timestamp -3599
transform 1 0 13984 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _268_
timestamp -3599
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _269_
timestamp -3599
transform 1 0 5704 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _270_
timestamp -3599
transform 1 0 10396 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _271_
timestamp -3599
transform 1 0 7544 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _272_
timestamp -3599
transform -1 0 3680 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _273_
timestamp -3599
transform 1 0 5428 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _274_
timestamp -3599
transform -1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _275_
timestamp -3599
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _276_
timestamp -3599
transform 1 0 5704 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _277_
timestamp -3599
transform 1 0 32660 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _278_
timestamp -3599
transform 1 0 30912 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _279_
timestamp -3599
transform 1 0 22080 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _280_
timestamp -3599
transform 1 0 23184 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _281_
timestamp -3599
transform 1 0 23828 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _282_
timestamp -3599
transform 1 0 24196 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _283_
timestamp -3599
transform -1 0 32016 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _284_
timestamp -3599
transform -1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _285_
timestamp -3599
transform 1 0 34776 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _286_
timestamp -3599
transform -1 0 31924 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _287_
timestamp -3599
transform -1 0 30820 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _288_
timestamp -3599
transform -1 0 31280 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _289_
timestamp -3599
transform -1 0 15640 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _290_
timestamp -3599
transform 1 0 14720 0 1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _291_
timestamp -3599
transform -1 0 16284 0 -1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _292_
timestamp -3599
transform -1 0 8464 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _293_
timestamp -3599
transform 1 0 11868 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _294_
timestamp -3599
transform 1 0 10764 0 1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _295_
timestamp -3599
transform 1 0 8924 0 1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _296_
timestamp -3599
transform -1 0 8832 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _297_
timestamp -3599
transform 1 0 9476 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _298_
timestamp -3599
transform 1 0 11592 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _299_
timestamp -3599
transform 1 0 12328 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _300_
timestamp -3599
transform 1 0 15088 0 1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _301_
timestamp -3599
transform 1 0 30452 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _302_
timestamp -3599
transform 1 0 30544 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _303_
timestamp -3599
transform 1 0 27968 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _304_
timestamp -3599
transform 1 0 27692 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _305_
timestamp -3599
transform -1 0 16008 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _306_
timestamp -3599
transform -1 0 15548 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _307_
timestamp -3599
transform 1 0 8464 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _308_
timestamp -3599
transform 1 0 11500 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _309_
timestamp -3599
transform 1 0 9936 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _310_
timestamp -3599
transform 1 0 8280 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _311_
timestamp -3599
transform 1 0 8924 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _312_
timestamp -3599
transform 1 0 9016 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _313_
timestamp -3599
transform 1 0 11592 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _314_
timestamp -3599
transform -1 0 13432 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _315_
timestamp -3599
transform -1 0 15272 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_1  _317_
timestamp -3599
transform 1 0 26864 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _318_
timestamp -3599
transform 1 0 26588 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _319_
timestamp -3599
transform 1 0 21436 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _320_
timestamp -3599
transform 1 0 12880 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _321_
timestamp -3599
transform 1 0 3772 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _322_
timestamp -3599
transform 1 0 4600 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _323_
timestamp -3599
transform 1 0 19228 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _324_
timestamp -3599
transform 1 0 19136 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _325_
timestamp -3599
transform 1 0 26956 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _326_
timestamp -3599
transform 1 0 28060 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _327_
timestamp -3599
transform 1 0 10764 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _328_
timestamp -3599
transform 1 0 2024 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _329_
timestamp -3599
transform 1 0 3588 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _330_
timestamp -3599
transform 1 0 10028 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _331_
timestamp -3599
transform 1 0 8464 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _332_
timestamp -3599
transform 1 0 4416 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _333_
timestamp -3599
transform -1 0 16560 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _334_
timestamp -3599
transform 1 0 28980 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _335_
timestamp -3599
transform 1 0 16928 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _336_
timestamp -3599
transform 1 0 6348 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _337_
timestamp -3599
transform 1 0 26312 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _338_
timestamp -3599
transform -1 0 30912 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _339_
timestamp -3599
transform 1 0 20792 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _340_
timestamp -3599
transform 1 0 7268 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _341_
timestamp -3599
transform 1 0 23460 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _342_
timestamp -3599
transform 1 0 23920 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _343_
timestamp -3599
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _344_
timestamp -3599
transform -1 0 36064 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _345_
timestamp -3599
transform -1 0 35604 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _346_
timestamp -3599
transform -1 0 33764 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _347_
timestamp -3599
transform -1 0 32292 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _348_
timestamp -3599
transform -1 0 32016 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _349_
timestamp -3599
transform -1 0 30912 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _350_
timestamp -3599
transform -1 0 26036 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _351_
timestamp -3599
transform -1 0 31740 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _352_
timestamp -3599
transform 1 0 38548 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _353_
timestamp -3599
transform 1 0 37260 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _354_
timestamp -3599
transform 1 0 38272 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _355_
timestamp -3599
transform 1 0 38272 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _356_
timestamp -3599
transform 1 0 38364 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _357_
timestamp -3599
transform 1 0 37352 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _358_
timestamp -3599
transform 1 0 38180 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _359_
timestamp -3599
transform 1 0 37720 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _360_
timestamp -3599
transform 1 0 38548 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _361_
timestamp -3599
transform 1 0 37444 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _362_
timestamp -3599
transform 1 0 37444 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _363_
timestamp -3599
transform -1 0 35604 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _364_
timestamp -3599
transform 1 0 37352 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _365_
timestamp -3599
transform 1 0 38364 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _366_
timestamp -3599
transform -1 0 37996 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _367_
timestamp -3599
transform 1 0 38548 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _368_
timestamp -3599
transform -1 0 36892 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _369_
timestamp -3599
transform -1 0 19504 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _370_
timestamp -3599
transform 1 0 5520 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _371_
timestamp -3599
transform -1 0 23460 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _372_
timestamp -3599
transform -1 0 29808 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _373_
timestamp -3599
transform -1 0 13616 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _374_
timestamp -3599
transform 1 0 3036 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _375_
timestamp -3599
transform -1 0 2576 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _376_
timestamp -3599
transform 1 0 10488 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _377_
timestamp -3599
transform -1 0 13984 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _378_
timestamp -3599
transform -1 0 5796 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _379_
timestamp -3599
transform -1 0 18676 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _380_
timestamp -3599
transform -1 0 27600 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _381_
timestamp -3599
transform -1 0 18860 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _382_
timestamp -3599
transform -1 0 24472 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _383_
timestamp -3599
transform -1 0 23368 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _384_
timestamp -3599
transform -1 0 27232 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _385_
timestamp -3599
transform -1 0 17756 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _386_
timestamp -3599
transform 1 0 8004 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _387_
timestamp -3599
transform -1 0 25300 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _388_
timestamp -3599
transform -1 0 21344 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _389_
timestamp -3599
transform -1 0 32752 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _390_
timestamp -3599
transform -1 0 36064 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _391_
timestamp -3599
transform -1 0 36064 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _392_
timestamp -3599
transform -1 0 34500 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _393_
timestamp -3599
transform -1 0 33028 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _394_
timestamp -3599
transform -1 0 33488 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _395_
timestamp -3599
transform 1 0 4968 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _396_
timestamp -3599
transform 1 0 18308 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _397_
timestamp -3599
transform -1 0 23184 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _398_
timestamp -3599
transform 1 0 15640 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _399_
timestamp -3599
transform 1 0 3220 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _400_
timestamp -3599
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _401_
timestamp -3599
transform -1 0 20884 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _402_
timestamp -3599
transform 1 0 21344 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _403_
timestamp -3599
transform -1 0 27140 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _404_
timestamp -3599
transform -1 0 26864 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _405_
timestamp -3599
transform 1 0 15640 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _406_
timestamp -3599
transform -1 0 2760 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _407_
timestamp -3599
transform -1 0 1656 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _408_
timestamp -3599
transform 1 0 11500 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _409_
timestamp -3599
transform -1 0 10028 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _410_
timestamp -3599
transform 1 0 2852 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _411_
timestamp -3599
transform -1 0 5520 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _412_
timestamp -3599
transform -1 0 30636 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _413_
timestamp -3599
transform 1 0 18860 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _414_
timestamp -3599
transform 1 0 6716 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _415_
timestamp -3599
transform -1 0 34592 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _416_
timestamp -3599
transform -1 0 32476 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _417_
timestamp -3599
transform 1 0 23736 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _418_
timestamp -3599
transform -1 0 24748 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _419_
timestamp -3599
transform 1 0 24012 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _420_
timestamp -3599
transform -1 0 25576 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _421_
timestamp -3599
transform 1 0 27600 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp -3599
transform 1 0 39008 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp -3599
transform -1 0 38180 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp -3599
transform -1 0 2300 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp -3599
transform 1 0 7360 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp -3599
transform -1 0 3312 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp -3599
transform -1 0 5520 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp -3599
transform -1 0 7084 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp -3599
transform -1 0 7728 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp -3599
transform -1 0 12880 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp -3599
transform 1 0 4600 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp -3599
transform -1 0 4048 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp -3599
transform 1 0 38180 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp -3599
transform -1 0 2576 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp -3599
transform 1 0 6808 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp -3599
transform -1 0 4784 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp -3599
transform -1 0 4876 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp -3599
transform 1 0 39008 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_UserCLK
timestamp -3599
transform 1 0 24472 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_UserCLK_regs
timestamp -3599
transform 1 0 19504 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_UserCLK
timestamp -3599
transform -1 0 26312 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_UserCLK_regs
timestamp -3599
transform -1 0 13984 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_UserCLK_regs
timestamp -3599
transform -1 0 13708 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_UserCLK_regs
timestamp -3599
transform 1 0 26312 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_UserCLK_regs
timestamp -3599
transform -1 0 22264 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_regs_0_UserCLK
timestamp -3599
transform -1 0 18492 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__bufinv_16  clkload0
timestamp -3599
transform 1 0 12328 0 -1 5440
box -38 -48 2246 592
use sky130_fd_sc_hd__clkinv_4  clkload1
timestamp -3599
transform -1 0 27600 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__bufinv_16  clkload2
timestamp -3599
transform 1 0 20424 0 1 7616
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_2  fanout33
timestamp -3599
transform 1 0 16652 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout34
timestamp -3599
transform -1 0 7820 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout35
timestamp -3599
transform -1 0 16284 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout36
timestamp -3599
transform 1 0 15272 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout37
timestamp -3599
transform -1 0 14812 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout38
timestamp -3599
transform 1 0 19504 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  fanout39
timestamp -3599
transform -1 0 32016 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout40
timestamp -3599
transform -1 0 3680 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout41
timestamp -3599
transform -1 0 29992 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout42
timestamp -3599
transform -1 0 30360 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout43
timestamp -3599
transform 1 0 30360 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23
timestamp -3599
transform 1 0 3220 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27
timestamp -3599
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33
timestamp -3599
transform 1 0 4140 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41
timestamp -3599
transform 1 0 4876 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57
timestamp -3599
transform 1 0 6348 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65
timestamp -3599
transform 1 0 7084 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71
timestamp -3599
transform 1 0 7636 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_94
timestamp -3599
transform 1 0 9752 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101
timestamp -3599
transform 1 0 10396 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_126
timestamp -3599
transform 1 0 12696 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_149
timestamp -3599
transform 1 0 14812 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_164
timestamp -3599
transform 1 0 16192 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_173
timestamp -3599
transform 1 0 17020 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_177
timestamp -3599
transform 1 0 17388 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_181
timestamp -3599
transform 1 0 17756 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_195
timestamp -3599
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_200
timestamp -3599
transform 1 0 19504 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_204
timestamp -3599
transform 1 0 19872 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_208
timestamp -3599
transform 1 0 20240 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_223
timestamp -3599
transform 1 0 21620 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_228
timestamp -3599
transform 1 0 22080 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_236
timestamp -3599
transform 1 0 22816 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_240
timestamp 1636964856
transform 1 0 23184 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_253
timestamp 1636964856
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_265
timestamp 1636964856
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp -3599
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_290
timestamp 1636964856
transform 1 0 27784 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_302
timestamp -3599
transform 1 0 28888 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_309
timestamp 1636964856
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_324
timestamp -3599
transform 1 0 30912 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_332
timestamp -3599
transform 1 0 31648 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_337
timestamp -3599
transform 1 0 32108 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_350
timestamp -3599
transform 1 0 33304 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_355
timestamp -3599
transform 1 0 33764 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_363
timestamp -3599
transform 1 0 34500 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_365
timestamp 1636964856
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_377
timestamp 1636964856
transform 1 0 35788 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_389
timestamp -3599
transform 1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_393
timestamp -3599
transform 1 0 37260 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_397
timestamp -3599
transform 1 0 37628 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3
timestamp -3599
transform 1 0 1380 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_22
timestamp 1636964856
transform 1 0 3128 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_34
timestamp -3599
transform 1 0 4232 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp -3599
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_66
timestamp -3599
transform 1 0 7176 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_97
timestamp -3599
transform 1 0 10028 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_164
timestamp -3599
transform 1 0 16192 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_169
timestamp -3599
transform 1 0 16652 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_222
timestamp -3599
transform 1 0 21528 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_225
timestamp -3599
transform 1 0 21804 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_266
timestamp -3599
transform 1 0 25576 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_271
timestamp -3599
transform 1 0 26036 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_296
timestamp 1636964856
transform 1 0 28336 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_308
timestamp -3599
transform 1 0 29440 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_321
timestamp -3599
transform 1 0 30636 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp -3599
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_349
timestamp -3599
transform 1 0 33212 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_375
timestamp -3599
transform 1 0 35604 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_383
timestamp -3599
transform 1 0 36340 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_389
timestamp -3599
transform 1 0 36892 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_393
timestamp 1636964856
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_405
timestamp -3599
transform 1 0 38364 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_22
timestamp -3599
transform 1 0 3128 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_33
timestamp -3599
transform 1 0 4140 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_51
timestamp 1636964856
transform 1 0 5796 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_63
timestamp -3599
transform 1 0 6900 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp -3599
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_94
timestamp -3599
transform 1 0 9752 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_116
timestamp -3599
transform 1 0 11776 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_136
timestamp -3599
transform 1 0 13616 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_161
timestamp -3599
transform 1 0 15916 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_169
timestamp -3599
transform 1 0 16652 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1636964856
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_209
timestamp -3599
transform 1 0 20332 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_213
timestamp -3599
transform 1 0 20700 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_220
timestamp -3599
transform 1 0 21344 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_224
timestamp -3599
transform 1 0 21712 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_253
timestamp -3599
transform 1 0 24380 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_275
timestamp -3599
transform 1 0 26404 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_306
timestamp -3599
transform 1 0 29256 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_321
timestamp -3599
transform 1 0 30636 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_336
timestamp -3599
transform 1 0 32016 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_340
timestamp -3599
transform 1 0 32384 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_344
timestamp 1636964856
transform 1 0 32752 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_356
timestamp -3599
transform 1 0 33856 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_365
timestamp -3599
transform 1 0 34684 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_373
timestamp -3599
transform 1 0 35420 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_380
timestamp 1636964856
transform 1 0 36064 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_392
timestamp 1636964856
transform 1 0 37168 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_404
timestamp -3599
transform 1 0 38272 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_3_13
timestamp -3599
transform 1 0 2300 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp -3599
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_66
timestamp -3599
transform 1 0 7176 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_74
timestamp -3599
transform 1 0 7912 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_78
timestamp -3599
transform 1 0 8280 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_129
timestamp -3599
transform 1 0 12972 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_161
timestamp -3599
transform 1 0 15916 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_198
timestamp 1636964856
transform 1 0 19320 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_219
timestamp -3599
transform 1 0 21252 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp -3599
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_234
timestamp -3599
transform 1 0 22632 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_249
timestamp -3599
transform 1 0 24012 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_254
timestamp -3599
transform 1 0 24472 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_3_269
timestamp -3599
transform 1 0 25852 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_277
timestamp -3599
transform 1 0 26588 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_281
timestamp -3599
transform 1 0 26956 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_303
timestamp -3599
transform 1 0 28980 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_309
timestamp -3599
transform 1 0 29532 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_324
timestamp 1636964856
transform 1 0 30912 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_337
timestamp -3599
transform 1 0 32108 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_341
timestamp -3599
transform 1 0 32476 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_347
timestamp 1636964856
transform 1 0 33028 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_359
timestamp -3599
transform 1 0 34132 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_388
timestamp -3599
transform 1 0 36800 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_393
timestamp -3599
transform 1 0 37260 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_397
timestamp 1636964856
transform 1 0 37628 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_409
timestamp -3599
transform 1 0 38732 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_11
timestamp -3599
transform 1 0 2116 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_18
timestamp -3599
transform 1 0 2760 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_22
timestamp -3599
transform 1 0 3128 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_26
timestamp -3599
transform 1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_73
timestamp -3599
transform 1 0 7820 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_85
timestamp -3599
transform 1 0 8924 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_112
timestamp -3599
transform 1 0 11408 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_130
timestamp -3599
transform 1 0 13064 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_146
timestamp -3599
transform 1 0 14536 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_191
timestamp -3599
transform 1 0 18676 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp -3599
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_236
timestamp -3599
transform 1 0 22816 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_240
timestamp -3599
transform 1 0 23184 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_250
timestamp -3599
transform 1 0 24104 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_262
timestamp -3599
transform 1 0 25208 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_270
timestamp -3599
transform 1 0 25944 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_306
timestamp -3599
transform 1 0 29256 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_309
timestamp -3599
transform 1 0 29532 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_323
timestamp -3599
transform 1 0 30820 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_336
timestamp -3599
transform 1 0 32016 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_355
timestamp -3599
transform 1 0 33764 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp -3599
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_380
timestamp 1636964856
transform 1 0 36064 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_392
timestamp -3599
transform 1 0 37168 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_397
timestamp -3599
transform 1 0 37628 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3
timestamp -3599
transform 1 0 1380 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_19
timestamp -3599
transform 1 0 2852 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_40
timestamp -3599
transform 1 0 4784 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_50
timestamp -3599
transform 1 0 5704 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_121
timestamp -3599
transform 1 0 12236 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_166
timestamp -3599
transform 1 0 16376 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_190
timestamp -3599
transform 1 0 18584 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_194
timestamp -3599
transform 1 0 18952 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp -3599
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_234
timestamp -3599
transform 1 0 22632 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_247
timestamp -3599
transform 1 0 23828 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_255
timestamp -3599
transform 1 0 24564 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_266
timestamp -3599
transform 1 0 25576 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_313
timestamp -3599
transform 1 0 29900 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_328
timestamp -3599
transform 1 0 31280 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1636964856
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1636964856
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1636964856
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp -3599
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp -3599
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_396
timestamp -3599
transform 1 0 37536 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3
timestamp -3599
transform 1 0 1380 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_37
timestamp -3599
transform 1 0 4508 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_62
timestamp -3599
transform 1 0 6808 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_67
timestamp -3599
transform 1 0 7268 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_73
timestamp -3599
transform 1 0 7820 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_85
timestamp -3599
transform 1 0 8924 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_110
timestamp -3599
transform 1 0 11224 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_177
timestamp -3599
transform 1 0 17388 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_213
timestamp -3599
transform 1 0 20700 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_243
timestamp -3599
transform 1 0 23460 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_6_262
timestamp 1636964856
transform 1 0 25208 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_274
timestamp -3599
transform 1 0 26312 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_6_292
timestamp -3599
transform 1 0 27968 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_315
timestamp -3599
transform 1 0 30084 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_328
timestamp -3599
transform 1 0 31280 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_332
timestamp -3599
transform 1 0 31648 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_339
timestamp -3599
transform 1 0 32292 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_347
timestamp -3599
transform 1 0 33028 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_352
timestamp 1636964856
transform 1 0 33488 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_365
timestamp -3599
transform 1 0 34684 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_378
timestamp 1636964856
transform 1 0 35880 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_390
timestamp -3599
transform 1 0 36984 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_394
timestamp -3599
transform 1 0 37352 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_401
timestamp -3599
transform 1 0 37996 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3
timestamp -3599
transform 1 0 1380 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_16
timestamp -3599
transform 1 0 2576 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_51
timestamp -3599
transform 1 0 5796 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_99
timestamp -3599
transform 1 0 10212 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_113
timestamp -3599
transform 1 0 11500 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_138
timestamp -3599
transform 1 0 13800 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_189
timestamp -3599
transform 1 0 18492 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_196
timestamp -3599
transform 1 0 19136 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp -3599
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_228
timestamp -3599
transform 1 0 22080 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_234
timestamp -3599
transform 1 0 22632 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_238
timestamp -3599
transform 1 0 23000 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_246
timestamp -3599
transform 1 0 23736 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_259
timestamp -3599
transform 1 0 24932 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_263
timestamp -3599
transform 1 0 25300 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_271
timestamp -3599
transform 1 0 26036 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_284
timestamp -3599
transform 1 0 27232 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_313
timestamp -3599
transform 1 0 29900 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_337
timestamp -3599
transform 1 0 32108 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_360
timestamp -3599
transform 1 0 34224 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_389
timestamp -3599
transform 1 0 36892 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1636964856
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_3
timestamp -3599
transform 1 0 1380 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_29
timestamp -3599
transform 1 0 3772 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_141
timestamp -3599
transform 1 0 14076 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_189
timestamp -3599
transform 1 0 18492 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_197
timestamp -3599
transform 1 0 19228 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_242
timestamp -3599
transform 1 0 23368 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_318
timestamp -3599
transform 1 0 30360 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_342
timestamp -3599
transform 1 0 32568 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_365
timestamp -3599
transform 1 0 34684 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_371
timestamp -3599
transform 1 0 35236 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_375
timestamp -3599
transform 1 0 35604 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_380
timestamp 1636964856
transform 1 0 36064 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_392
timestamp -3599
transform 1 0 37168 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_9_36
timestamp -3599
transform 1 0 4416 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_57
timestamp -3599
transform 1 0 6348 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_94
timestamp -3599
transform 1 0 9752 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_191
timestamp -3599
transform 1 0 18676 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_233
timestamp -3599
transform 1 0 22540 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_290
timestamp -3599
transform 1 0 27784 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_318
timestamp -3599
transform 1 0 30360 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_364
timestamp 1636964856
transform 1 0 34592 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_376
timestamp 1636964856
transform 1 0 35696 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_388
timestamp -3599
transform 1 0 36800 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_393
timestamp -3599
transform 1 0 37260 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_23
timestamp -3599
transform 1 0 3220 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_62
timestamp -3599
transform 1 0 6808 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_138
timestamp -3599
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_189
timestamp -3599
transform 1 0 18492 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_250
timestamp -3599
transform 1 0 24104 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_253
timestamp -3599
transform 1 0 24380 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_306
timestamp -3599
transform 1 0 29256 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_335
timestamp -3599
transform 1 0 31924 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_359
timestamp -3599
transform 1 0 34132 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp -3599
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_369
timestamp -3599
transform 1 0 35052 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_10_379
timestamp -3599
transform 1 0 35972 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_385
timestamp -3599
transform 1 0 36524 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_391
timestamp -3599
transform 1 0 37076 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_403
timestamp -3599
transform 1 0 38180 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_29
timestamp -3599
transform 1 0 3772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_41
timestamp -3599
transform 1 0 4876 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_57
timestamp -3599
transform 1 0 6348 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_85
timestamp -3599
transform 1 0 8924 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_98
timestamp -3599
transform 1 0 10120 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_113
timestamp -3599
transform 1 0 11500 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_197
timestamp -3599
transform 1 0 19228 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_210
timestamp -3599
transform 1 0 20424 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_220
timestamp -3599
transform 1 0 21344 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_225
timestamp -3599
transform 1 0 21804 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_267
timestamp -3599
transform 1 0 25668 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_317
timestamp -3599
transform 1 0 30268 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp -3599
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_340
timestamp -3599
transform 1 0 32384 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_362
timestamp -3599
transform 1 0 34408 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_389
timestamp -3599
transform 1 0 36892 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_409
timestamp -3599
transform 1 0 38732 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1
timestamp -3599
transform 1 0 21988 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp -3599
transform -1 0 14720 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp -3599
transform -1 0 20424 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp -3599
transform 1 0 14076 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp -3599
transform -1 0 13984 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp -3599
transform -1 0 13800 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp -3599
transform -1 0 11224 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp -3599
transform -1 0 17388 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp -3599
transform 1 0 15640 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp -3599
transform -1 0 10120 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp -3599
transform -1 0 11408 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp -3599
transform 1 0 21804 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp -3599
transform -1 0 10212 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp -3599
transform -1 0 11868 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp -3599
transform -1 0 11408 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp -3599
transform -1 0 10304 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp -3599
transform -1 0 19964 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp -3599
transform -1 0 21344 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp -3599
transform 1 0 32292 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input1
timestamp -3599
transform 1 0 2944 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input2
timestamp -3599
transform 1 0 1748 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input3
timestamp -3599
transform 1 0 1748 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp -3599
transform 1 0 2024 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp -3599
transform 1 0 2208 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp -3599
transform 1 0 2576 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input7
timestamp -3599
transform 1 0 2300 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input8
timestamp -3599
transform 1 0 1748 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input9
timestamp -3599
transform 1 0 2024 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input10
timestamp -3599
transform 1 0 2116 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input11
timestamp -3599
transform 1 0 2484 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input12
timestamp -3599
transform 1 0 1840 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input13
timestamp -3599
transform 1 0 1380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input14
timestamp -3599
transform 1 0 1840 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input15
timestamp -3599
transform 1 0 1380 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input16
timestamp -3599
transform 1 0 1380 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input17
timestamp -3599
transform 1 0 1380 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input18
timestamp -3599
transform 1 0 2300 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input19
timestamp -3599
transform 1 0 2208 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input20
timestamp -3599
transform 1 0 1472 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input21
timestamp -3599
transform 1 0 1748 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input22
timestamp -3599
transform 1 0 1472 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input23
timestamp -3599
transform 1 0 2484 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input24
timestamp -3599
transform 1 0 2300 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input25
timestamp -3599
transform 1 0 1840 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input26
timestamp -3599
transform 1 0 2208 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp -3599
transform -1 0 2944 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input28
timestamp -3599
transform 1 0 2576 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input29
timestamp -3599
transform 1 0 1472 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input30
timestamp -3599
transform 1 0 2852 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input31
timestamp -3599
transform 1 0 2852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input32
timestamp -3599
transform 1 0 1380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input33
timestamp -3599
transform 1 0 1380 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input34
timestamp -3599
transform 1 0 19964 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input35
timestamp -3599
transform 1 0 21804 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input36
timestamp -3599
transform 1 0 17480 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp -3599
transform -1 0 19044 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input38
timestamp -3599
transform -1 0 17296 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp -3599
transform 1 0 18584 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp -3599
transform -1 0 19688 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp -3599
transform -1 0 21712 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input42
timestamp -3599
transform -1 0 18584 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp -3599
transform 1 0 24012 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input44
timestamp -3599
transform 1 0 23736 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp -3599
transform 1 0 25484 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp -3599
transform 1 0 27968 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp -3599
transform 1 0 24196 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input48
timestamp -3599
transform 1 0 17112 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp -3599
transform 1 0 18860 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input50
timestamp -3599
transform -1 0 15088 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input51
timestamp -3599
transform -1 0 16560 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input52
timestamp -3599
transform -1 0 19136 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input53
timestamp -3599
transform -1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input54
timestamp -3599
transform -1 0 19504 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input55
timestamp -3599
transform -1 0 19136 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp -3599
transform 1 0 28428 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp -3599
transform -1 0 29256 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp -3599
transform -1 0 31924 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input59
timestamp -3599
transform 1 0 29164 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp -3599
transform -1 0 29808 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input61
timestamp -3599
transform 1 0 29164 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input62
timestamp -3599
transform -1 0 32384 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp -3599
transform -1 0 26864 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp -3599
transform 1 0 25760 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input65
timestamp -3599
transform 1 0 25484 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input66
timestamp -3599
transform -1 0 28428 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input67
timestamp -3599
transform -1 0 26588 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input68
timestamp -3599
transform -1 0 28980 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input69
timestamp -3599
transform 1 0 29992 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input70
timestamp -3599
transform 1 0 27140 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input71
timestamp -3599
transform -1 0 27692 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input72
timestamp -3599
transform 1 0 32016 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input73
timestamp -3599
transform -1 0 33764 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input74
timestamp -3599
transform -1 0 32292 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input75
timestamp -3599
transform 1 0 33580 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input76
timestamp -3599
transform -1 0 32568 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input77
timestamp -3599
transform -1 0 34132 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input78
timestamp -3599
transform -1 0 34040 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input79
timestamp -3599
transform 1 0 27416 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input80
timestamp -3599
transform -1 0 30360 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input81
timestamp -3599
transform -1 0 30360 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input82
timestamp -3599
transform 1 0 32660 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input83
timestamp -3599
transform -1 0 30084 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input84
timestamp -3599
transform -1 0 33212 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input85
timestamp -3599
transform -1 0 32016 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input86
timestamp -3599
transform 1 0 31740 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input87
timestamp -3599
transform -1 0 33488 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output88
timestamp -3599
transform 1 0 38088 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp -3599
transform 1 0 39192 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp -3599
transform 1 0 38640 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp -3599
transform 1 0 39192 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp -3599
transform 1 0 38824 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp -3599
transform 1 0 39192 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp -3599
transform 1 0 38824 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp -3599
transform 1 0 39192 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp -3599
transform 1 0 38640 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp -3599
transform 1 0 38456 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp -3599
transform 1 0 39192 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp -3599
transform 1 0 37720 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output100
timestamp -3599
transform 1 0 37720 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output101
timestamp -3599
transform 1 0 39192 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp -3599
transform 1 0 38824 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output103
timestamp -3599
transform 1 0 39192 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output104
timestamp -3599
transform 1 0 39192 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output105
timestamp -3599
transform 1 0 38824 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output106
timestamp -3599
transform 1 0 38456 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output107
timestamp -3599
transform 1 0 38824 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output108
timestamp -3599
transform 1 0 39192 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output109
timestamp -3599
transform 1 0 38456 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output110
timestamp -3599
transform 1 0 38456 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output111
timestamp -3599
transform 1 0 38824 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output112
timestamp -3599
transform 1 0 38088 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output113
timestamp -3599
transform 1 0 38824 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output114
timestamp -3599
transform 1 0 39192 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output115
timestamp -3599
transform 1 0 38824 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output116
timestamp -3599
transform 1 0 39192 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output117
timestamp -3599
transform 1 0 38824 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output118
timestamp -3599
transform 1 0 39192 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output119
timestamp -3599
transform 1 0 38824 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output120
timestamp -3599
transform 1 0 32568 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output121
timestamp -3599
transform -1 0 36524 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output122
timestamp -3599
transform -1 0 35972 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output123
timestamp -3599
transform -1 0 36892 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output124
timestamp -3599
transform -1 0 36524 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output125
timestamp -3599
transform 1 0 37260 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output126
timestamp -3599
transform -1 0 37076 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output127
timestamp -3599
transform -1 0 37996 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output128
timestamp -3599
transform 1 0 37996 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output129
timestamp -3599
transform -1 0 38732 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output130
timestamp -3599
transform 1 0 37812 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output131
timestamp -3599
transform 1 0 32936 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output132
timestamp -3599
transform 1 0 33304 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output133
timestamp -3599
transform -1 0 34040 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output134
timestamp -3599
transform -1 0 34408 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output135
timestamp -3599
transform -1 0 35052 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output136
timestamp -3599
transform -1 0 35420 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output137
timestamp -3599
transform -1 0 35052 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output138
timestamp -3599
transform -1 0 35788 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output139
timestamp -3599
transform -1 0 36156 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output140
timestamp -3599
transform -1 0 2668 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output141
timestamp -3599
transform -1 0 2576 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output142
timestamp -3599
transform -1 0 1840 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output143
timestamp -3599
transform -1 0 3680 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output144
timestamp -3599
transform -1 0 4508 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output145
timestamp -3599
transform -1 0 2024 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output146
timestamp -3599
transform 1 0 2944 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output147
timestamp -3599
transform 1 0 3312 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output148
timestamp -3599
transform -1 0 4140 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output149
timestamp -3599
transform -1 0 3312 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output150
timestamp -3599
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output151
timestamp -3599
transform 1 0 2576 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output152
timestamp -3599
transform -1 0 6256 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output153
timestamp -3599
transform -1 0 4324 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output154
timestamp -3599
transform -1 0 7268 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output155
timestamp -3599
transform -1 0 7452 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output156
timestamp -3599
transform -1 0 7820 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output157
timestamp -3599
transform -1 0 2944 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output158
timestamp -3599
transform -1 0 6256 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output159
timestamp -3599
transform -1 0 4692 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output160
timestamp -3599
transform -1 0 7084 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output161
timestamp -3599
transform -1 0 6716 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output162
timestamp -3599
transform 1 0 4968 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output163
timestamp -3599
transform 1 0 5888 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output164
timestamp -3599
transform -1 0 7360 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output165
timestamp -3599
transform -1 0 8832 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output166
timestamp -3599
transform -1 0 8096 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output167
timestamp -3599
transform -1 0 6808 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output168
timestamp -3599
transform -1 0 6900 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output169
timestamp -3599
transform -1 0 5428 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output170
timestamp -3599
transform -1 0 8372 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output171
timestamp -3599
transform -1 0 7820 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output172
timestamp -3599
transform 1 0 3312 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output173
timestamp -3599
transform -1 0 5060 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output174
timestamp -3599
transform 1 0 4784 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output175
timestamp -3599
transform 1 0 5520 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output176
timestamp -3599
transform 1 0 7084 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output177
timestamp -3599
transform 1 0 7728 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output178
timestamp -3599
transform -1 0 15456 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output179
timestamp -3599
transform -1 0 15824 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output180
timestamp -3599
transform -1 0 16192 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output181
timestamp -3599
transform -1 0 16560 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output182
timestamp -3599
transform -1 0 18308 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output183
timestamp -3599
transform -1 0 18492 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output184
timestamp -3599
transform 1 0 16008 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output185
timestamp -3599
transform 1 0 8096 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output186
timestamp -3599
transform -1 0 9384 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output187
timestamp -3599
transform 1 0 13432 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output188
timestamp -3599
transform 1 0 10304 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output189
timestamp -3599
transform 1 0 11592 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output190
timestamp -3599
transform 1 0 12880 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output191
timestamp -3599
transform -1 0 13616 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output192
timestamp -3599
transform 1 0 13616 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output193
timestamp -3599
transform -1 0 4140 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  output194
timestamp -3599
transform -1 0 34316 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output195
timestamp -3599
transform -1 0 4876 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output196
timestamp -3599
transform -1 0 5980 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output197
timestamp -3599
transform -1 0 16192 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output198
timestamp -3599
transform -1 0 17020 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output199
timestamp -3599
transform -1 0 7084 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output200
timestamp -3599
transform -1 0 8096 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output201
timestamp -3599
transform -1 0 8464 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output202
timestamp -3599
transform -1 0 10396 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output203
timestamp -3599
transform 1 0 11040 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output204
timestamp -3599
transform -1 0 12696 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output205
timestamp -3599
transform -1 0 14444 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output206
timestamp -3599
transform 1 0 14076 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_12
timestamp -3599
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp -3599
transform -1 0 39836 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_13
timestamp -3599
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp -3599
transform -1 0 39836 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_14
timestamp -3599
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp -3599
transform -1 0 39836 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_15
timestamp -3599
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp -3599
transform -1 0 39836 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_16
timestamp -3599
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp -3599
transform -1 0 39836 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_17
timestamp -3599
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp -3599
transform -1 0 39836 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_18
timestamp -3599
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp -3599
transform -1 0 39836 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_19
timestamp -3599
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp -3599
transform -1 0 39836 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_20
timestamp -3599
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp -3599
transform -1 0 39836 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_21
timestamp -3599
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp -3599
transform -1 0 39836 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_22
timestamp -3599
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp -3599
transform -1 0 39836 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_23
timestamp -3599
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp -3599
transform -1 0 39836 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  S_EF_ADC12_207
timestamp -3599
transform 1 0 16376 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_24
timestamp -3599
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_25
timestamp -3599
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_26
timestamp -3599
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_27
timestamp -3599
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_28
timestamp -3599
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_29
timestamp -3599
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_30
timestamp -3599
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_31
timestamp -3599
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_32
timestamp -3599
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_33
timestamp -3599
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_34
timestamp -3599
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_35
timestamp -3599
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_36
timestamp -3599
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_37
timestamp -3599
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_38
timestamp -3599
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_39
timestamp -3599
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_40
timestamp -3599
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_41
timestamp -3599
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_42
timestamp -3599
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_43
timestamp -3599
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_44
timestamp -3599
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_45
timestamp -3599
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_46
timestamp -3599
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_47
timestamp -3599
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_48
timestamp -3599
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_49
timestamp -3599
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_50
timestamp -3599
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_51
timestamp -3599
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_52
timestamp -3599
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_53
timestamp -3599
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_54
timestamp -3599
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_55
timestamp -3599
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_56
timestamp -3599
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_57
timestamp -3599
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_58
timestamp -3599
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_59
timestamp -3599
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_60
timestamp -3599
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_61
timestamp -3599
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_62
timestamp -3599
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_63
timestamp -3599
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_64
timestamp -3599
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_65
timestamp -3599
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_66
timestamp -3599
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_67
timestamp -3599
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_68
timestamp -3599
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_69
timestamp -3599
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_70
timestamp -3599
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_71
timestamp -3599
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_72
timestamp -3599
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_73
timestamp -3599
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_74
timestamp -3599
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_75
timestamp -3599
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_76
timestamp -3599
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_77
timestamp -3599
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_78
timestamp -3599
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_79
timestamp -3599
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_80
timestamp -3599
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_81
timestamp -3599
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_82
timestamp -3599
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_83
timestamp -3599
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_84
timestamp -3599
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_85
timestamp -3599
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_86
timestamp -3599
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_87
timestamp -3599
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_88
timestamp -3599
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_89
timestamp -3599
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_90
timestamp -3599
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_91
timestamp -3599
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_92
timestamp -3599
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_93
timestamp -3599
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_94
timestamp -3599
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_95
timestamp -3599
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_96
timestamp -3599
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_97
timestamp -3599
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_98
timestamp -3599
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_99
timestamp -3599
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_100
timestamp -3599
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_101
timestamp -3599
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_102
timestamp -3599
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_103
timestamp -3599
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_104
timestamp -3599
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_105
timestamp -3599
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_106
timestamp -3599
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_107
timestamp -3599
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_108
timestamp -3599
transform 1 0 3680 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_109
timestamp -3599
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_110
timestamp -3599
transform 1 0 8832 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_111
timestamp -3599
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_112
timestamp -3599
transform 1 0 13984 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_113
timestamp -3599
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_114
timestamp -3599
transform 1 0 19136 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_115
timestamp -3599
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_116
timestamp -3599
transform 1 0 24288 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_117
timestamp -3599
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_118
timestamp -3599
transform 1 0 29440 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_119
timestamp -3599
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_120
timestamp -3599
transform 1 0 34592 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_121
timestamp -3599
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
<< labels >>
flabel metal2 s 1122 0 1178 56 0 FreeSans 224 0 0 0 CMP_top
port 0 nsew signal input
flabel metal2 s 17590 11194 17646 11250 0 FreeSans 224 0 0 0 Co
port 1 nsew signal output
flabel metal3 s 0 1368 120 1488 0 FreeSans 480 0 0 0 FrameData[0]
port 2 nsew signal input
flabel metal3 s 0 4088 120 4208 0 FreeSans 480 0 0 0 FrameData[10]
port 3 nsew signal input
flabel metal3 s 0 4360 120 4480 0 FreeSans 480 0 0 0 FrameData[11]
port 4 nsew signal input
flabel metal3 s 0 4632 120 4752 0 FreeSans 480 0 0 0 FrameData[12]
port 5 nsew signal input
flabel metal3 s 0 4904 120 5024 0 FreeSans 480 0 0 0 FrameData[13]
port 6 nsew signal input
flabel metal3 s 0 5176 120 5296 0 FreeSans 480 0 0 0 FrameData[14]
port 7 nsew signal input
flabel metal3 s 0 5448 120 5568 0 FreeSans 480 0 0 0 FrameData[15]
port 8 nsew signal input
flabel metal3 s 0 5720 120 5840 0 FreeSans 480 0 0 0 FrameData[16]
port 9 nsew signal input
flabel metal3 s 0 5992 120 6112 0 FreeSans 480 0 0 0 FrameData[17]
port 10 nsew signal input
flabel metal3 s 0 6264 120 6384 0 FreeSans 480 0 0 0 FrameData[18]
port 11 nsew signal input
flabel metal3 s 0 6536 120 6656 0 FreeSans 480 0 0 0 FrameData[19]
port 12 nsew signal input
flabel metal3 s 0 1640 120 1760 0 FreeSans 480 0 0 0 FrameData[1]
port 13 nsew signal input
flabel metal3 s 0 6808 120 6928 0 FreeSans 480 0 0 0 FrameData[20]
port 14 nsew signal input
flabel metal3 s 0 7080 120 7200 0 FreeSans 480 0 0 0 FrameData[21]
port 15 nsew signal input
flabel metal3 s 0 7352 120 7472 0 FreeSans 480 0 0 0 FrameData[22]
port 16 nsew signal input
flabel metal3 s 0 7624 120 7744 0 FreeSans 480 0 0 0 FrameData[23]
port 17 nsew signal input
flabel metal3 s 0 7896 120 8016 0 FreeSans 480 0 0 0 FrameData[24]
port 18 nsew signal input
flabel metal3 s 0 8168 120 8288 0 FreeSans 480 0 0 0 FrameData[25]
port 19 nsew signal input
flabel metal3 s 0 8440 120 8560 0 FreeSans 480 0 0 0 FrameData[26]
port 20 nsew signal input
flabel metal3 s 0 8712 120 8832 0 FreeSans 480 0 0 0 FrameData[27]
port 21 nsew signal input
flabel metal3 s 0 8984 120 9104 0 FreeSans 480 0 0 0 FrameData[28]
port 22 nsew signal input
flabel metal3 s 0 9256 120 9376 0 FreeSans 480 0 0 0 FrameData[29]
port 23 nsew signal input
flabel metal3 s 0 1912 120 2032 0 FreeSans 480 0 0 0 FrameData[2]
port 24 nsew signal input
flabel metal3 s 0 9528 120 9648 0 FreeSans 480 0 0 0 FrameData[30]
port 25 nsew signal input
flabel metal3 s 0 9800 120 9920 0 FreeSans 480 0 0 0 FrameData[31]
port 26 nsew signal input
flabel metal3 s 0 2184 120 2304 0 FreeSans 480 0 0 0 FrameData[3]
port 27 nsew signal input
flabel metal3 s 0 2456 120 2576 0 FreeSans 480 0 0 0 FrameData[4]
port 28 nsew signal input
flabel metal3 s 0 2728 120 2848 0 FreeSans 480 0 0 0 FrameData[5]
port 29 nsew signal input
flabel metal3 s 0 3000 120 3120 0 FreeSans 480 0 0 0 FrameData[6]
port 30 nsew signal input
flabel metal3 s 0 3272 120 3392 0 FreeSans 480 0 0 0 FrameData[7]
port 31 nsew signal input
flabel metal3 s 0 3544 120 3664 0 FreeSans 480 0 0 0 FrameData[8]
port 32 nsew signal input
flabel metal3 s 0 3816 120 3936 0 FreeSans 480 0 0 0 FrameData[9]
port 33 nsew signal input
flabel metal3 s 40880 1368 41000 1488 0 FreeSans 480 0 0 0 FrameData_O[0]
port 34 nsew signal output
flabel metal3 s 40880 4088 41000 4208 0 FreeSans 480 0 0 0 FrameData_O[10]
port 35 nsew signal output
flabel metal3 s 40880 4360 41000 4480 0 FreeSans 480 0 0 0 FrameData_O[11]
port 36 nsew signal output
flabel metal3 s 40880 4632 41000 4752 0 FreeSans 480 0 0 0 FrameData_O[12]
port 37 nsew signal output
flabel metal3 s 40880 4904 41000 5024 0 FreeSans 480 0 0 0 FrameData_O[13]
port 38 nsew signal output
flabel metal3 s 40880 5176 41000 5296 0 FreeSans 480 0 0 0 FrameData_O[14]
port 39 nsew signal output
flabel metal3 s 40880 5448 41000 5568 0 FreeSans 480 0 0 0 FrameData_O[15]
port 40 nsew signal output
flabel metal3 s 40880 5720 41000 5840 0 FreeSans 480 0 0 0 FrameData_O[16]
port 41 nsew signal output
flabel metal3 s 40880 5992 41000 6112 0 FreeSans 480 0 0 0 FrameData_O[17]
port 42 nsew signal output
flabel metal3 s 40880 6264 41000 6384 0 FreeSans 480 0 0 0 FrameData_O[18]
port 43 nsew signal output
flabel metal3 s 40880 6536 41000 6656 0 FreeSans 480 0 0 0 FrameData_O[19]
port 44 nsew signal output
flabel metal3 s 40880 1640 41000 1760 0 FreeSans 480 0 0 0 FrameData_O[1]
port 45 nsew signal output
flabel metal3 s 40880 6808 41000 6928 0 FreeSans 480 0 0 0 FrameData_O[20]
port 46 nsew signal output
flabel metal3 s 40880 7080 41000 7200 0 FreeSans 480 0 0 0 FrameData_O[21]
port 47 nsew signal output
flabel metal3 s 40880 7352 41000 7472 0 FreeSans 480 0 0 0 FrameData_O[22]
port 48 nsew signal output
flabel metal3 s 40880 7624 41000 7744 0 FreeSans 480 0 0 0 FrameData_O[23]
port 49 nsew signal output
flabel metal3 s 40880 7896 41000 8016 0 FreeSans 480 0 0 0 FrameData_O[24]
port 50 nsew signal output
flabel metal3 s 40880 8168 41000 8288 0 FreeSans 480 0 0 0 FrameData_O[25]
port 51 nsew signal output
flabel metal3 s 40880 8440 41000 8560 0 FreeSans 480 0 0 0 FrameData_O[26]
port 52 nsew signal output
flabel metal3 s 40880 8712 41000 8832 0 FreeSans 480 0 0 0 FrameData_O[27]
port 53 nsew signal output
flabel metal3 s 40880 8984 41000 9104 0 FreeSans 480 0 0 0 FrameData_O[28]
port 54 nsew signal output
flabel metal3 s 40880 9256 41000 9376 0 FreeSans 480 0 0 0 FrameData_O[29]
port 55 nsew signal output
flabel metal3 s 40880 1912 41000 2032 0 FreeSans 480 0 0 0 FrameData_O[2]
port 56 nsew signal output
flabel metal3 s 40880 9528 41000 9648 0 FreeSans 480 0 0 0 FrameData_O[30]
port 57 nsew signal output
flabel metal3 s 40880 9800 41000 9920 0 FreeSans 480 0 0 0 FrameData_O[31]
port 58 nsew signal output
flabel metal3 s 40880 2184 41000 2304 0 FreeSans 480 0 0 0 FrameData_O[3]
port 59 nsew signal output
flabel metal3 s 40880 2456 41000 2576 0 FreeSans 480 0 0 0 FrameData_O[4]
port 60 nsew signal output
flabel metal3 s 40880 2728 41000 2848 0 FreeSans 480 0 0 0 FrameData_O[5]
port 61 nsew signal output
flabel metal3 s 40880 3000 41000 3120 0 FreeSans 480 0 0 0 FrameData_O[6]
port 62 nsew signal output
flabel metal3 s 40880 3272 41000 3392 0 FreeSans 480 0 0 0 FrameData_O[7]
port 63 nsew signal output
flabel metal3 s 40880 3544 41000 3664 0 FreeSans 480 0 0 0 FrameData_O[8]
port 64 nsew signal output
flabel metal3 s 40880 3816 41000 3936 0 FreeSans 480 0 0 0 FrameData_O[9]
port 65 nsew signal output
flabel metal2 s 18786 0 18842 56 0 FreeSans 224 0 0 0 FrameStrobe[0]
port 66 nsew signal input
flabel metal2 s 29826 0 29882 56 0 FreeSans 224 0 0 0 FrameStrobe[10]
port 67 nsew signal input
flabel metal2 s 30930 0 30986 56 0 FreeSans 224 0 0 0 FrameStrobe[11]
port 68 nsew signal input
flabel metal2 s 32034 0 32090 56 0 FreeSans 224 0 0 0 FrameStrobe[12]
port 69 nsew signal input
flabel metal2 s 33138 0 33194 56 0 FreeSans 224 0 0 0 FrameStrobe[13]
port 70 nsew signal input
flabel metal2 s 34242 0 34298 56 0 FreeSans 224 0 0 0 FrameStrobe[14]
port 71 nsew signal input
flabel metal2 s 35346 0 35402 56 0 FreeSans 224 0 0 0 FrameStrobe[15]
port 72 nsew signal input
flabel metal2 s 36450 0 36506 56 0 FreeSans 224 0 0 0 FrameStrobe[16]
port 73 nsew signal input
flabel metal2 s 37554 0 37610 56 0 FreeSans 224 0 0 0 FrameStrobe[17]
port 74 nsew signal input
flabel metal2 s 38658 0 38714 56 0 FreeSans 224 0 0 0 FrameStrobe[18]
port 75 nsew signal input
flabel metal2 s 39762 0 39818 56 0 FreeSans 224 0 0 0 FrameStrobe[19]
port 76 nsew signal input
flabel metal2 s 19890 0 19946 56 0 FreeSans 224 0 0 0 FrameStrobe[1]
port 77 nsew signal input
flabel metal2 s 20994 0 21050 56 0 FreeSans 224 0 0 0 FrameStrobe[2]
port 78 nsew signal input
flabel metal2 s 22098 0 22154 56 0 FreeSans 224 0 0 0 FrameStrobe[3]
port 79 nsew signal input
flabel metal2 s 23202 0 23258 56 0 FreeSans 224 0 0 0 FrameStrobe[4]
port 80 nsew signal input
flabel metal2 s 24306 0 24362 56 0 FreeSans 224 0 0 0 FrameStrobe[5]
port 81 nsew signal input
flabel metal2 s 25410 0 25466 56 0 FreeSans 224 0 0 0 FrameStrobe[6]
port 82 nsew signal input
flabel metal2 s 26514 0 26570 56 0 FreeSans 224 0 0 0 FrameStrobe[7]
port 83 nsew signal input
flabel metal2 s 27618 0 27674 56 0 FreeSans 224 0 0 0 FrameStrobe[8]
port 84 nsew signal input
flabel metal2 s 28722 0 28778 56 0 FreeSans 224 0 0 0 FrameStrobe[9]
port 85 nsew signal input
flabel metal2 s 32494 11194 32550 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[0]
port 86 nsew signal output
flabel metal2 s 35254 11194 35310 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[10]
port 87 nsew signal output
flabel metal2 s 35530 11194 35586 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[11]
port 88 nsew signal output
flabel metal2 s 35806 11194 35862 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[12]
port 89 nsew signal output
flabel metal2 s 36082 11194 36138 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[13]
port 90 nsew signal output
flabel metal2 s 36358 11194 36414 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[14]
port 91 nsew signal output
flabel metal2 s 36634 11194 36690 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[15]
port 92 nsew signal output
flabel metal2 s 36910 11194 36966 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[16]
port 93 nsew signal output
flabel metal2 s 37186 11194 37242 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[17]
port 94 nsew signal output
flabel metal2 s 37462 11194 37518 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[18]
port 95 nsew signal output
flabel metal2 s 37738 11194 37794 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[19]
port 96 nsew signal output
flabel metal2 s 32770 11194 32826 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[1]
port 97 nsew signal output
flabel metal2 s 33046 11194 33102 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[2]
port 98 nsew signal output
flabel metal2 s 33322 11194 33378 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[3]
port 99 nsew signal output
flabel metal2 s 33598 11194 33654 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[4]
port 100 nsew signal output
flabel metal2 s 33874 11194 33930 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[5]
port 101 nsew signal output
flabel metal2 s 34150 11194 34206 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[6]
port 102 nsew signal output
flabel metal2 s 34426 11194 34482 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[7]
port 103 nsew signal output
flabel metal2 s 34702 11194 34758 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[8]
port 104 nsew signal output
flabel metal2 s 34978 11194 35034 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[9]
port 105 nsew signal output
flabel metal2 s 2226 0 2282 56 0 FreeSans 224 0 0 0 HOLD_top
port 106 nsew signal output
flabel metal2 s 3238 11194 3294 11250 0 FreeSans 224 0 0 0 N1BEG[0]
port 107 nsew signal output
flabel metal2 s 3514 11194 3570 11250 0 FreeSans 224 0 0 0 N1BEG[1]
port 108 nsew signal output
flabel metal2 s 3790 11194 3846 11250 0 FreeSans 224 0 0 0 N1BEG[2]
port 109 nsew signal output
flabel metal2 s 4066 11194 4122 11250 0 FreeSans 224 0 0 0 N1BEG[3]
port 110 nsew signal output
flabel metal2 s 4342 11194 4398 11250 0 FreeSans 224 0 0 0 N2BEG[0]
port 111 nsew signal output
flabel metal2 s 4618 11194 4674 11250 0 FreeSans 224 0 0 0 N2BEG[1]
port 112 nsew signal output
flabel metal2 s 4894 11194 4950 11250 0 FreeSans 224 0 0 0 N2BEG[2]
port 113 nsew signal output
flabel metal2 s 5170 11194 5226 11250 0 FreeSans 224 0 0 0 N2BEG[3]
port 114 nsew signal output
flabel metal2 s 5446 11194 5502 11250 0 FreeSans 224 0 0 0 N2BEG[4]
port 115 nsew signal output
flabel metal2 s 5722 11194 5778 11250 0 FreeSans 224 0 0 0 N2BEG[5]
port 116 nsew signal output
flabel metal2 s 5998 11194 6054 11250 0 FreeSans 224 0 0 0 N2BEG[6]
port 117 nsew signal output
flabel metal2 s 6274 11194 6330 11250 0 FreeSans 224 0 0 0 N2BEG[7]
port 118 nsew signal output
flabel metal2 s 6550 11194 6606 11250 0 FreeSans 224 0 0 0 N2BEGb[0]
port 119 nsew signal output
flabel metal2 s 6826 11194 6882 11250 0 FreeSans 224 0 0 0 N2BEGb[1]
port 120 nsew signal output
flabel metal2 s 7102 11194 7158 11250 0 FreeSans 224 0 0 0 N2BEGb[2]
port 121 nsew signal output
flabel metal2 s 7378 11194 7434 11250 0 FreeSans 224 0 0 0 N2BEGb[3]
port 122 nsew signal output
flabel metal2 s 7654 11194 7710 11250 0 FreeSans 224 0 0 0 N2BEGb[4]
port 123 nsew signal output
flabel metal2 s 7930 11194 7986 11250 0 FreeSans 224 0 0 0 N2BEGb[5]
port 124 nsew signal output
flabel metal2 s 8206 11194 8262 11250 0 FreeSans 224 0 0 0 N2BEGb[6]
port 125 nsew signal output
flabel metal2 s 8482 11194 8538 11250 0 FreeSans 224 0 0 0 N2BEGb[7]
port 126 nsew signal output
flabel metal2 s 8758 11194 8814 11250 0 FreeSans 224 0 0 0 N4BEG[0]
port 127 nsew signal output
flabel metal2 s 11518 11194 11574 11250 0 FreeSans 224 0 0 0 N4BEG[10]
port 128 nsew signal output
flabel metal2 s 11794 11194 11850 11250 0 FreeSans 224 0 0 0 N4BEG[11]
port 129 nsew signal output
flabel metal2 s 12070 11194 12126 11250 0 FreeSans 224 0 0 0 N4BEG[12]
port 130 nsew signal output
flabel metal2 s 12346 11194 12402 11250 0 FreeSans 224 0 0 0 N4BEG[13]
port 131 nsew signal output
flabel metal2 s 12622 11194 12678 11250 0 FreeSans 224 0 0 0 N4BEG[14]
port 132 nsew signal output
flabel metal2 s 12898 11194 12954 11250 0 FreeSans 224 0 0 0 N4BEG[15]
port 133 nsew signal output
flabel metal2 s 9034 11194 9090 11250 0 FreeSans 224 0 0 0 N4BEG[1]
port 134 nsew signal output
flabel metal2 s 9310 11194 9366 11250 0 FreeSans 224 0 0 0 N4BEG[2]
port 135 nsew signal output
flabel metal2 s 9586 11194 9642 11250 0 FreeSans 224 0 0 0 N4BEG[3]
port 136 nsew signal output
flabel metal2 s 9862 11194 9918 11250 0 FreeSans 224 0 0 0 N4BEG[4]
port 137 nsew signal output
flabel metal2 s 10138 11194 10194 11250 0 FreeSans 224 0 0 0 N4BEG[5]
port 138 nsew signal output
flabel metal2 s 10414 11194 10470 11250 0 FreeSans 224 0 0 0 N4BEG[6]
port 139 nsew signal output
flabel metal2 s 10690 11194 10746 11250 0 FreeSans 224 0 0 0 N4BEG[7]
port 140 nsew signal output
flabel metal2 s 10966 11194 11022 11250 0 FreeSans 224 0 0 0 N4BEG[8]
port 141 nsew signal output
flabel metal2 s 11242 11194 11298 11250 0 FreeSans 224 0 0 0 N4BEG[9]
port 142 nsew signal output
flabel metal2 s 13174 11194 13230 11250 0 FreeSans 224 0 0 0 NN4BEG[0]
port 143 nsew signal output
flabel metal2 s 15934 11194 15990 11250 0 FreeSans 224 0 0 0 NN4BEG[10]
port 144 nsew signal output
flabel metal2 s 16210 11194 16266 11250 0 FreeSans 224 0 0 0 NN4BEG[11]
port 145 nsew signal output
flabel metal2 s 16486 11194 16542 11250 0 FreeSans 224 0 0 0 NN4BEG[12]
port 146 nsew signal output
flabel metal2 s 16762 11194 16818 11250 0 FreeSans 224 0 0 0 NN4BEG[13]
port 147 nsew signal output
flabel metal2 s 17038 11194 17094 11250 0 FreeSans 224 0 0 0 NN4BEG[14]
port 148 nsew signal output
flabel metal2 s 17314 11194 17370 11250 0 FreeSans 224 0 0 0 NN4BEG[15]
port 149 nsew signal output
flabel metal2 s 13450 11194 13506 11250 0 FreeSans 224 0 0 0 NN4BEG[1]
port 150 nsew signal output
flabel metal2 s 13726 11194 13782 11250 0 FreeSans 224 0 0 0 NN4BEG[2]
port 151 nsew signal output
flabel metal2 s 14002 11194 14058 11250 0 FreeSans 224 0 0 0 NN4BEG[3]
port 152 nsew signal output
flabel metal2 s 14278 11194 14334 11250 0 FreeSans 224 0 0 0 NN4BEG[4]
port 153 nsew signal output
flabel metal2 s 14554 11194 14610 11250 0 FreeSans 224 0 0 0 NN4BEG[5]
port 154 nsew signal output
flabel metal2 s 14830 11194 14886 11250 0 FreeSans 224 0 0 0 NN4BEG[6]
port 155 nsew signal output
flabel metal2 s 15106 11194 15162 11250 0 FreeSans 224 0 0 0 NN4BEG[7]
port 156 nsew signal output
flabel metal2 s 15382 11194 15438 11250 0 FreeSans 224 0 0 0 NN4BEG[8]
port 157 nsew signal output
flabel metal2 s 15658 11194 15714 11250 0 FreeSans 224 0 0 0 NN4BEG[9]
port 158 nsew signal output
flabel metal2 s 3330 0 3386 56 0 FreeSans 224 0 0 0 RESET_top
port 159 nsew signal output
flabel metal2 s 17866 11194 17922 11250 0 FreeSans 224 0 0 0 S1END[0]
port 160 nsew signal input
flabel metal2 s 18142 11194 18198 11250 0 FreeSans 224 0 0 0 S1END[1]
port 161 nsew signal input
flabel metal2 s 18418 11194 18474 11250 0 FreeSans 224 0 0 0 S1END[2]
port 162 nsew signal input
flabel metal2 s 18694 11194 18750 11250 0 FreeSans 224 0 0 0 S1END[3]
port 163 nsew signal input
flabel metal2 s 21178 11194 21234 11250 0 FreeSans 224 0 0 0 S2END[0]
port 164 nsew signal input
flabel metal2 s 21454 11194 21510 11250 0 FreeSans 224 0 0 0 S2END[1]
port 165 nsew signal input
flabel metal2 s 21730 11194 21786 11250 0 FreeSans 224 0 0 0 S2END[2]
port 166 nsew signal input
flabel metal2 s 22006 11194 22062 11250 0 FreeSans 224 0 0 0 S2END[3]
port 167 nsew signal input
flabel metal2 s 22282 11194 22338 11250 0 FreeSans 224 0 0 0 S2END[4]
port 168 nsew signal input
flabel metal2 s 22558 11194 22614 11250 0 FreeSans 224 0 0 0 S2END[5]
port 169 nsew signal input
flabel metal2 s 22834 11194 22890 11250 0 FreeSans 224 0 0 0 S2END[6]
port 170 nsew signal input
flabel metal2 s 23110 11194 23166 11250 0 FreeSans 224 0 0 0 S2END[7]
port 171 nsew signal input
flabel metal2 s 18970 11194 19026 11250 0 FreeSans 224 0 0 0 S2MID[0]
port 172 nsew signal input
flabel metal2 s 19246 11194 19302 11250 0 FreeSans 224 0 0 0 S2MID[1]
port 173 nsew signal input
flabel metal2 s 19522 11194 19578 11250 0 FreeSans 224 0 0 0 S2MID[2]
port 174 nsew signal input
flabel metal2 s 19798 11194 19854 11250 0 FreeSans 224 0 0 0 S2MID[3]
port 175 nsew signal input
flabel metal2 s 20074 11194 20130 11250 0 FreeSans 224 0 0 0 S2MID[4]
port 176 nsew signal input
flabel metal2 s 20350 11194 20406 11250 0 FreeSans 224 0 0 0 S2MID[5]
port 177 nsew signal input
flabel metal2 s 20626 11194 20682 11250 0 FreeSans 224 0 0 0 S2MID[6]
port 178 nsew signal input
flabel metal2 s 20902 11194 20958 11250 0 FreeSans 224 0 0 0 S2MID[7]
port 179 nsew signal input
flabel metal2 s 23386 11194 23442 11250 0 FreeSans 224 0 0 0 S4END[0]
port 180 nsew signal input
flabel metal2 s 26146 11194 26202 11250 0 FreeSans 224 0 0 0 S4END[10]
port 181 nsew signal input
flabel metal2 s 26422 11194 26478 11250 0 FreeSans 224 0 0 0 S4END[11]
port 182 nsew signal input
flabel metal2 s 26698 11194 26754 11250 0 FreeSans 224 0 0 0 S4END[12]
port 183 nsew signal input
flabel metal2 s 26974 11194 27030 11250 0 FreeSans 224 0 0 0 S4END[13]
port 184 nsew signal input
flabel metal2 s 27250 11194 27306 11250 0 FreeSans 224 0 0 0 S4END[14]
port 185 nsew signal input
flabel metal2 s 27526 11194 27582 11250 0 FreeSans 224 0 0 0 S4END[15]
port 186 nsew signal input
flabel metal2 s 23662 11194 23718 11250 0 FreeSans 224 0 0 0 S4END[1]
port 187 nsew signal input
flabel metal2 s 23938 11194 23994 11250 0 FreeSans 224 0 0 0 S4END[2]
port 188 nsew signal input
flabel metal2 s 24214 11194 24270 11250 0 FreeSans 224 0 0 0 S4END[3]
port 189 nsew signal input
flabel metal2 s 24490 11194 24546 11250 0 FreeSans 224 0 0 0 S4END[4]
port 190 nsew signal input
flabel metal2 s 24766 11194 24822 11250 0 FreeSans 224 0 0 0 S4END[5]
port 191 nsew signal input
flabel metal2 s 25042 11194 25098 11250 0 FreeSans 224 0 0 0 S4END[6]
port 192 nsew signal input
flabel metal2 s 25318 11194 25374 11250 0 FreeSans 224 0 0 0 S4END[7]
port 193 nsew signal input
flabel metal2 s 25594 11194 25650 11250 0 FreeSans 224 0 0 0 S4END[8]
port 194 nsew signal input
flabel metal2 s 25870 11194 25926 11250 0 FreeSans 224 0 0 0 S4END[9]
port 195 nsew signal input
flabel metal2 s 27802 11194 27858 11250 0 FreeSans 224 0 0 0 SS4END[0]
port 196 nsew signal input
flabel metal2 s 30562 11194 30618 11250 0 FreeSans 224 0 0 0 SS4END[10]
port 197 nsew signal input
flabel metal2 s 30838 11194 30894 11250 0 FreeSans 224 0 0 0 SS4END[11]
port 198 nsew signal input
flabel metal2 s 31114 11194 31170 11250 0 FreeSans 224 0 0 0 SS4END[12]
port 199 nsew signal input
flabel metal2 s 31390 11194 31446 11250 0 FreeSans 224 0 0 0 SS4END[13]
port 200 nsew signal input
flabel metal2 s 31666 11194 31722 11250 0 FreeSans 224 0 0 0 SS4END[14]
port 201 nsew signal input
flabel metal2 s 31942 11194 31998 11250 0 FreeSans 224 0 0 0 SS4END[15]
port 202 nsew signal input
flabel metal2 s 28078 11194 28134 11250 0 FreeSans 224 0 0 0 SS4END[1]
port 203 nsew signal input
flabel metal2 s 28354 11194 28410 11250 0 FreeSans 224 0 0 0 SS4END[2]
port 204 nsew signal input
flabel metal2 s 28630 11194 28686 11250 0 FreeSans 224 0 0 0 SS4END[3]
port 205 nsew signal input
flabel metal2 s 28906 11194 28962 11250 0 FreeSans 224 0 0 0 SS4END[4]
port 206 nsew signal input
flabel metal2 s 29182 11194 29238 11250 0 FreeSans 224 0 0 0 SS4END[5]
port 207 nsew signal input
flabel metal2 s 29458 11194 29514 11250 0 FreeSans 224 0 0 0 SS4END[6]
port 208 nsew signal input
flabel metal2 s 29734 11194 29790 11250 0 FreeSans 224 0 0 0 SS4END[7]
port 209 nsew signal input
flabel metal2 s 30010 11194 30066 11250 0 FreeSans 224 0 0 0 SS4END[8]
port 210 nsew signal input
flabel metal2 s 30286 11194 30342 11250 0 FreeSans 224 0 0 0 SS4END[9]
port 211 nsew signal input
flabel metal2 s 17682 0 17738 56 0 FreeSans 224 0 0 0 UserCLK
port 212 nsew signal input
flabel metal2 s 32218 11194 32274 11250 0 FreeSans 224 0 0 0 UserCLKo
port 213 nsew signal output
flabel metal2 s 4434 0 4490 56 0 FreeSans 224 0 0 0 VALUE_top0
port 214 nsew signal output
flabel metal2 s 5538 0 5594 56 0 FreeSans 224 0 0 0 VALUE_top1
port 215 nsew signal output
flabel metal2 s 15474 0 15530 56 0 FreeSans 224 0 0 0 VALUE_top10
port 216 nsew signal output
flabel metal2 s 16578 0 16634 56 0 FreeSans 224 0 0 0 VALUE_top11
port 217 nsew signal output
flabel metal2 s 6642 0 6698 56 0 FreeSans 224 0 0 0 VALUE_top2
port 218 nsew signal output
flabel metal2 s 7746 0 7802 56 0 FreeSans 224 0 0 0 VALUE_top3
port 219 nsew signal output
flabel metal2 s 8850 0 8906 56 0 FreeSans 224 0 0 0 VALUE_top4
port 220 nsew signal output
flabel metal2 s 9954 0 10010 56 0 FreeSans 224 0 0 0 VALUE_top5
port 221 nsew signal output
flabel metal2 s 11058 0 11114 56 0 FreeSans 224 0 0 0 VALUE_top6
port 222 nsew signal output
flabel metal2 s 12162 0 12218 56 0 FreeSans 224 0 0 0 VALUE_top7
port 223 nsew signal output
flabel metal2 s 13266 0 13322 56 0 FreeSans 224 0 0 0 VALUE_top8
port 224 nsew signal output
flabel metal2 s 14370 0 14426 56 0 FreeSans 224 0 0 0 VALUE_top9
port 225 nsew signal output
flabel metal4 s 3004 0 3324 11250 0 FreeSans 1920 90 0 0 VGND
port 226 nsew ground bidirectional
flabel metal4 s 3004 0 3324 60 0 FreeSans 480 0 0 0 VGND
port 226 nsew ground bidirectional
flabel metal4 s 3004 11190 3324 11250 0 FreeSans 480 0 0 0 VGND
port 226 nsew ground bidirectional
flabel metal4 s 9004 0 9324 11250 0 FreeSans 1920 90 0 0 VGND
port 226 nsew ground bidirectional
flabel metal4 s 9004 0 9324 60 0 FreeSans 480 0 0 0 VGND
port 226 nsew ground bidirectional
flabel metal4 s 9004 11190 9324 11250 0 FreeSans 480 0 0 0 VGND
port 226 nsew ground bidirectional
flabel metal4 s 15004 0 15324 11250 0 FreeSans 1920 90 0 0 VGND
port 226 nsew ground bidirectional
flabel metal4 s 15004 0 15324 60 0 FreeSans 480 0 0 0 VGND
port 226 nsew ground bidirectional
flabel metal4 s 15004 11190 15324 11250 0 FreeSans 480 0 0 0 VGND
port 226 nsew ground bidirectional
flabel metal4 s 21004 0 21324 11250 0 FreeSans 1920 90 0 0 VGND
port 226 nsew ground bidirectional
flabel metal4 s 21004 0 21324 60 0 FreeSans 480 0 0 0 VGND
port 226 nsew ground bidirectional
flabel metal4 s 21004 11190 21324 11250 0 FreeSans 480 0 0 0 VGND
port 226 nsew ground bidirectional
flabel metal4 s 27004 0 27324 11250 0 FreeSans 1920 90 0 0 VGND
port 226 nsew ground bidirectional
flabel metal4 s 27004 0 27324 60 0 FreeSans 480 0 0 0 VGND
port 226 nsew ground bidirectional
flabel metal4 s 27004 11190 27324 11250 0 FreeSans 480 0 0 0 VGND
port 226 nsew ground bidirectional
flabel metal4 s 33004 0 33324 11250 0 FreeSans 1920 90 0 0 VGND
port 226 nsew ground bidirectional
flabel metal4 s 33004 0 33324 60 0 FreeSans 480 0 0 0 VGND
port 226 nsew ground bidirectional
flabel metal4 s 33004 11190 33324 11250 0 FreeSans 480 0 0 0 VGND
port 226 nsew ground bidirectional
flabel metal4 s 39004 0 39324 11250 0 FreeSans 1920 90 0 0 VGND
port 226 nsew ground bidirectional
flabel metal4 s 39004 0 39324 60 0 FreeSans 480 0 0 0 VGND
port 226 nsew ground bidirectional
flabel metal4 s 39004 11190 39324 11250 0 FreeSans 480 0 0 0 VGND
port 226 nsew ground bidirectional
flabel metal4 s 1944 0 2264 11250 0 FreeSans 1920 90 0 0 VPWR
port 227 nsew power bidirectional
flabel metal4 s 1944 0 2264 60 0 FreeSans 480 0 0 0 VPWR
port 227 nsew power bidirectional
flabel metal4 s 1944 11190 2264 11250 0 FreeSans 480 0 0 0 VPWR
port 227 nsew power bidirectional
flabel metal4 s 7944 0 8264 11250 0 FreeSans 1920 90 0 0 VPWR
port 227 nsew power bidirectional
flabel metal4 s 7944 0 8264 60 0 FreeSans 480 0 0 0 VPWR
port 227 nsew power bidirectional
flabel metal4 s 7944 11190 8264 11250 0 FreeSans 480 0 0 0 VPWR
port 227 nsew power bidirectional
flabel metal4 s 13944 0 14264 11250 0 FreeSans 1920 90 0 0 VPWR
port 227 nsew power bidirectional
flabel metal4 s 13944 0 14264 60 0 FreeSans 480 0 0 0 VPWR
port 227 nsew power bidirectional
flabel metal4 s 13944 11190 14264 11250 0 FreeSans 480 0 0 0 VPWR
port 227 nsew power bidirectional
flabel metal4 s 19944 0 20264 11250 0 FreeSans 1920 90 0 0 VPWR
port 227 nsew power bidirectional
flabel metal4 s 19944 0 20264 60 0 FreeSans 480 0 0 0 VPWR
port 227 nsew power bidirectional
flabel metal4 s 19944 11190 20264 11250 0 FreeSans 480 0 0 0 VPWR
port 227 nsew power bidirectional
flabel metal4 s 25944 0 26264 11250 0 FreeSans 1920 90 0 0 VPWR
port 227 nsew power bidirectional
flabel metal4 s 25944 0 26264 60 0 FreeSans 480 0 0 0 VPWR
port 227 nsew power bidirectional
flabel metal4 s 25944 11190 26264 11250 0 FreeSans 480 0 0 0 VPWR
port 227 nsew power bidirectional
flabel metal4 s 31944 0 32264 11250 0 FreeSans 1920 90 0 0 VPWR
port 227 nsew power bidirectional
flabel metal4 s 31944 0 32264 60 0 FreeSans 480 0 0 0 VPWR
port 227 nsew power bidirectional
flabel metal4 s 31944 11190 32264 11250 0 FreeSans 480 0 0 0 VPWR
port 227 nsew power bidirectional
flabel metal4 s 37944 0 38264 11250 0 FreeSans 1920 90 0 0 VPWR
port 227 nsew power bidirectional
flabel metal4 s 37944 0 38264 60 0 FreeSans 480 0 0 0 VPWR
port 227 nsew power bidirectional
flabel metal4 s 37944 11190 38264 11250 0 FreeSans 480 0 0 0 VPWR
port 227 nsew power bidirectional
rlabel metal1 20470 8704 20470 8704 0 VGND
rlabel metal1 20470 8160 20470 8160 0 VPWR
rlabel metal2 1150 1296 1150 1296 0 CMP_top
rlabel metal3 528 1428 528 1428 0 FrameData[0]
rlabel metal3 252 4148 252 4148 0 FrameData[10]
rlabel metal3 620 4420 620 4420 0 FrameData[11]
rlabel metal3 620 4692 620 4692 0 FrameData[12]
rlabel metal3 712 4964 712 4964 0 FrameData[13]
rlabel metal3 344 5236 344 5236 0 FrameData[14]
rlabel metal3 574 5508 574 5508 0 FrameData[15]
rlabel metal3 298 5780 298 5780 0 FrameData[16]
rlabel metal3 666 6052 666 6052 0 FrameData[17]
rlabel metal3 206 6324 206 6324 0 FrameData[18]
rlabel metal3 528 6596 528 6596 0 FrameData[19]
rlabel metal3 252 1700 252 1700 0 FrameData[1]
rlabel metal3 574 6868 574 6868 0 FrameData[20]
rlabel metal3 436 7140 436 7140 0 FrameData[21]
rlabel metal3 436 7412 436 7412 0 FrameData[22]
rlabel metal3 436 7684 436 7684 0 FrameData[23]
rlabel metal3 666 7956 666 7956 0 FrameData[24]
rlabel metal3 620 8228 620 8228 0 FrameData[25]
rlabel metal3 482 8500 482 8500 0 FrameData[26]
rlabel metal3 160 8772 160 8772 0 FrameData[27]
rlabel metal3 252 9044 252 9044 0 FrameData[28]
rlabel via2 114 9316 114 9316 0 FrameData[29]
rlabel metal3 1218 1972 1218 1972 0 FrameData[2]
rlabel metal3 712 9588 712 9588 0 FrameData[30]
rlabel metal3 1218 9860 1218 9860 0 FrameData[31]
rlabel metal3 712 2244 712 2244 0 FrameData[3]
rlabel metal3 1356 2516 1356 2516 0 FrameData[4]
rlabel metal3 344 2788 344 2788 0 FrameData[5]
rlabel metal3 1402 3060 1402 3060 0 FrameData[6]
rlabel metal3 1402 3332 1402 3332 0 FrameData[7]
rlabel metal3 436 3604 436 3604 0 FrameData[8]
rlabel metal3 436 3876 436 3876 0 FrameData[9]
rlabel metal3 39614 1428 39614 1428 0 FrameData_O[0]
rlabel metal3 40166 4148 40166 4148 0 FrameData_O[10]
rlabel metal3 40396 4420 40396 4420 0 FrameData_O[11]
rlabel metal3 40166 4692 40166 4692 0 FrameData_O[12]
rlabel metal3 39982 4964 39982 4964 0 FrameData_O[13]
rlabel metal3 40166 5236 40166 5236 0 FrameData_O[14]
rlabel metal3 40442 5508 40442 5508 0 FrameData_O[15]
rlabel metal3 40166 5780 40166 5780 0 FrameData_O[16]
rlabel metal3 39890 6052 39890 6052 0 FrameData_O[17]
rlabel metal3 39798 6324 39798 6324 0 FrameData_O[18]
rlabel metal2 39422 6511 39422 6511 0 FrameData_O[19]
rlabel metal3 39430 1700 39430 1700 0 FrameData_O[1]
rlabel metal3 39752 6868 39752 6868 0 FrameData_O[20]
rlabel metal3 40166 7140 40166 7140 0 FrameData_O[21]
rlabel metal3 39936 7412 39936 7412 0 FrameData_O[22]
rlabel metal3 40166 7684 40166 7684 0 FrameData_O[23]
rlabel metal3 40166 7956 40166 7956 0 FrameData_O[24]
rlabel metal3 39982 8228 39982 8228 0 FrameData_O[25]
rlabel metal2 38686 8279 38686 8279 0 FrameData_O[26]
rlabel metal1 39330 7514 39330 7514 0 FrameData_O[27]
rlabel metal1 39468 6630 39468 6630 0 FrameData_O[28]
rlabel metal1 38778 7514 38778 7514 0 FrameData_O[29]
rlabel metal3 39936 1972 39936 1972 0 FrameData_O[2]
rlabel metal1 39192 6630 39192 6630 0 FrameData_O[30]
rlabel metal1 38318 7480 38318 7480 0 FrameData_O[31]
rlabel metal3 40442 2244 40442 2244 0 FrameData_O[3]
rlabel metal3 40166 2516 40166 2516 0 FrameData_O[4]
rlabel metal3 39982 2788 39982 2788 0 FrameData_O[5]
rlabel metal3 40166 3060 40166 3060 0 FrameData_O[6]
rlabel metal3 40442 3332 40442 3332 0 FrameData_O[7]
rlabel metal3 40166 3604 40166 3604 0 FrameData_O[8]
rlabel metal3 39982 3876 39982 3876 0 FrameData_O[9]
rlabel metal2 18814 871 18814 871 0 FrameStrobe[0]
rlabel metal2 35742 1754 35742 1754 0 FrameStrobe[10]
rlabel via2 37306 5763 37306 5763 0 FrameStrobe[11]
rlabel metal2 32062 55 32062 55 0 FrameStrobe[12]
rlabel metal2 33166 55 33166 55 0 FrameStrobe[13]
rlabel metal1 34822 3094 34822 3094 0 FrameStrobe[14]
rlabel metal1 35650 4454 35650 4454 0 FrameStrobe[15]
rlabel metal1 37536 4522 37536 4522 0 FrameStrobe[16]
rlabel metal1 37674 5610 37674 5610 0 FrameStrobe[17]
rlabel metal1 38732 5202 38732 5202 0 FrameStrobe[18]
rlabel metal1 38226 2890 38226 2890 0 FrameStrobe[19]
rlabel metal2 19918 1228 19918 1228 0 FrameStrobe[1]
rlabel metal2 21022 599 21022 599 0 FrameStrobe[2]
rlabel metal1 39146 2958 39146 2958 0 FrameStrobe[3]
rlabel metal1 37628 5202 37628 5202 0 FrameStrobe[4]
rlabel metal1 38548 5678 38548 5678 0 FrameStrobe[5]
rlabel metal2 38502 4216 38502 4216 0 FrameStrobe[6]
rlabel metal1 37858 6290 37858 6290 0 FrameStrobe[7]
rlabel metal2 36662 3519 36662 3519 0 FrameStrobe[8]
rlabel metal2 38042 6477 38042 6477 0 FrameStrobe[9]
rlabel metal1 32798 8500 32798 8500 0 FrameStrobe_O[0]
rlabel metal1 35788 8262 35788 8262 0 FrameStrobe_O[10]
rlabel metal1 35650 8058 35650 8058 0 FrameStrobe_O[11]
rlabel metal1 36248 8602 36248 8602 0 FrameStrobe_O[12]
rlabel metal1 36202 8058 36202 8058 0 FrameStrobe_O[13]
rlabel metal1 37306 8262 37306 8262 0 FrameStrobe_O[14]
rlabel metal1 36754 8058 36754 8058 0 FrameStrobe_O[15]
rlabel metal1 37352 8602 37352 8602 0 FrameStrobe_O[16]
rlabel metal1 37720 8330 37720 8330 0 FrameStrobe_O[17]
rlabel metal1 38502 8568 38502 8568 0 FrameStrobe_O[18]
rlabel metal1 37904 8058 37904 8058 0 FrameStrobe_O[19]
rlabel metal1 32982 8330 32982 8330 0 FrameStrobe_O[1]
rlabel metal1 34040 8602 34040 8602 0 FrameStrobe_O[2]
rlabel metal2 33810 8534 33810 8534 0 FrameStrobe_O[3]
rlabel metal1 33902 8330 33902 8330 0 FrameStrobe_O[4]
rlabel metal1 34822 8568 34822 8568 0 FrameStrobe_O[5]
rlabel metal1 35144 8602 35144 8602 0 FrameStrobe_O[6]
rlabel metal1 34684 8058 34684 8058 0 FrameStrobe_O[7]
rlabel metal1 35144 8330 35144 8330 0 FrameStrobe_O[8]
rlabel metal1 35926 8364 35926 8364 0 FrameStrobe_O[9]
rlabel metal2 2254 1160 2254 1160 0 HOLD_top
rlabel metal1 32936 2278 32936 2278 0 Inst_EF_ADC12.VALID
rlabel metal1 21160 7378 21160 7378 0 Inst_EF_ADC12.curr_state\[0\]
rlabel metal2 16698 8228 16698 8228 0 Inst_EF_ADC12.curr_state\[1\]
rlabel metal2 18630 7956 18630 7956 0 Inst_EF_ADC12.curr_state\[2\]
rlabel metal1 21850 8398 21850 8398 0 Inst_EF_ADC12.curr_state\[3\]
rlabel metal1 20746 8398 20746 8398 0 Inst_EF_ADC12.curr_state\[5\]
rlabel metal1 14214 5882 14214 5882 0 Inst_EF_ADC12.next_bit\[0\]
rlabel metal2 14214 6426 14214 6426 0 Inst_EF_ADC12.next_bit\[10\]
rlabel metal1 10258 4012 10258 4012 0 Inst_EF_ADC12.next_bit\[1\]
rlabel metal2 12926 4692 12926 4692 0 Inst_EF_ADC12.next_bit\[2\]
rlabel metal1 11408 7174 11408 7174 0 Inst_EF_ADC12.next_bit\[3\]
rlabel metal1 10028 7174 10028 7174 0 Inst_EF_ADC12.next_bit\[4\]
rlabel metal2 10166 6460 10166 6460 0 Inst_EF_ADC12.next_bit\[5\]
rlabel metal2 10442 6120 10442 6120 0 Inst_EF_ADC12.next_bit\[6\]
rlabel metal1 12880 6086 12880 6086 0 Inst_EF_ADC12.next_bit\[7\]
rlabel metal1 11914 6834 11914 6834 0 Inst_EF_ADC12.next_bit\[8\]
rlabel metal2 13846 6766 13846 6766 0 Inst_EF_ADC12.next_bit\[9\]
rlabel metal2 32614 7616 32614 7616 0 Inst_EF_ADC12.sample_counter\[0\]
rlabel metal1 30176 7854 30176 7854 0 Inst_EF_ADC12.sample_counter\[1\]
rlabel metal1 29670 7310 29670 7310 0 Inst_EF_ADC12.sample_counter\[2\]
rlabel metal1 29624 6970 29624 6970 0 Inst_EF_ADC12.sample_counter\[3\]
rlabel metal2 14490 4590 14490 4590 0 Inst_EF_ADC12.shift_value\[0\]
rlabel metal2 5566 5916 5566 5916 0 Inst_S_EF_ADC12_ConfigMem.Inst_frame0_bit0.Q
rlabel metal1 18216 5746 18216 5746 0 Inst_S_EF_ADC12_ConfigMem.Inst_frame0_bit1.Q
rlabel metal1 15134 2482 15134 2482 0 Inst_S_EF_ADC12_ConfigMem.Inst_frame0_bit10.Q
rlabel metal2 4738 8228 4738 8228 0 Inst_S_EF_ADC12_ConfigMem.Inst_frame0_bit11.Q
rlabel metal1 7498 7956 7498 7956 0 Inst_S_EF_ADC12_ConfigMem.Inst_frame0_bit12.Q
rlabel metal2 10810 3876 10810 3876 0 Inst_S_EF_ADC12_ConfigMem.Inst_frame0_bit13.Q
rlabel metal1 8832 2822 8832 2822 0 Inst_S_EF_ADC12_ConfigMem.Inst_frame0_bit14.Q
rlabel metal1 2990 5882 2990 5882 0 Inst_S_EF_ADC12_ConfigMem.Inst_frame0_bit15.Q
rlabel metal1 7130 6868 7130 6868 0 Inst_S_EF_ADC12_ConfigMem.Inst_frame0_bit16.Q
rlabel metal2 29670 3162 29670 3162 0 Inst_S_EF_ADC12_ConfigMem.Inst_frame0_bit17.Q
rlabel metal1 17894 5100 17894 5100 0 Inst_S_EF_ADC12_ConfigMem.Inst_frame0_bit18.Q
rlabel metal2 6578 4794 6578 4794 0 Inst_S_EF_ADC12_ConfigMem.Inst_frame0_bit19.Q
rlabel metal1 23690 2924 23690 2924 0 Inst_S_EF_ADC12_ConfigMem.Inst_frame0_bit2.Q
rlabel metal1 33810 6834 33810 6834 0 Inst_S_EF_ADC12_ConfigMem.Inst_frame0_bit20.Q
rlabel metal1 32706 4692 32706 4692 0 Inst_S_EF_ADC12_ConfigMem.Inst_frame0_bit21.Q
rlabel metal2 23138 3876 23138 3876 0 Inst_S_EF_ADC12_ConfigMem.Inst_frame0_bit22.Q
rlabel metal1 25116 3570 25116 3570 0 Inst_S_EF_ADC12_ConfigMem.Inst_frame0_bit23.Q
rlabel metal2 24978 5916 24978 5916 0 Inst_S_EF_ADC12_ConfigMem.Inst_frame0_bit24.Q
rlabel metal2 25254 3604 25254 3604 0 Inst_S_EF_ADC12_ConfigMem.Inst_frame0_bit25.Q
rlabel metal2 30682 3808 30682 3808 0 Inst_S_EF_ADC12_ConfigMem.Inst_frame0_bit26.Q
rlabel metal1 33235 4794 33235 4794 0 Inst_S_EF_ADC12_ConfigMem.Inst_frame0_bit27.Q
rlabel metal1 23276 5202 23276 5202 0 Inst_S_EF_ADC12_ConfigMem.Inst_frame0_bit28.Q
rlabel metal2 28566 3808 28566 3808 0 Inst_S_EF_ADC12_ConfigMem.Inst_frame0_bit29.Q
rlabel metal2 13846 3604 13846 3604 0 Inst_S_EF_ADC12_ConfigMem.Inst_frame0_bit3.Q
rlabel metal2 28934 4420 28934 4420 0 Inst_S_EF_ADC12_ConfigMem.Inst_frame0_bit30.Q
rlabel metal1 29762 5338 29762 5338 0 Inst_S_EF_ADC12_ConfigMem.Inst_frame0_bit31.Q
rlabel metal1 3864 4250 3864 4250 0 Inst_S_EF_ADC12_ConfigMem.Inst_frame0_bit4.Q
rlabel metal2 6946 2890 6946 2890 0 Inst_S_EF_ADC12_ConfigMem.Inst_frame0_bit5.Q
rlabel metal2 20976 4046 20976 4046 0 Inst_S_EF_ADC12_ConfigMem.Inst_frame0_bit6.Q
rlabel metal2 22402 5049 22402 5049 0 Inst_S_EF_ADC12_ConfigMem.Inst_frame0_bit7.Q
rlabel metal1 27554 7344 27554 7344 0 Inst_S_EF_ADC12_ConfigMem.Inst_frame0_bit8.Q
rlabel metal3 27416 2788 27416 2788 0 Inst_S_EF_ADC12_ConfigMem.Inst_frame0_bit9.Q
rlabel metal2 29762 6868 29762 6868 0 Inst_S_EF_ADC12_ConfigMem.Inst_frame1_bit0.Q
rlabel metal1 28796 5746 28796 5746 0 Inst_S_EF_ADC12_ConfigMem.Inst_frame1_bit1.Q
rlabel metal1 13294 2822 13294 2822 0 Inst_S_EF_ADC12_ConfigMem.Inst_frame1_bit10.Q
rlabel metal1 4462 6868 4462 6868 0 Inst_S_EF_ADC12_ConfigMem.Inst_frame1_bit11.Q
rlabel metal2 5198 7718 5198 7718 0 Inst_S_EF_ADC12_ConfigMem.Inst_frame1_bit12.Q
rlabel metal1 11730 2482 11730 2482 0 Inst_S_EF_ADC12_ConfigMem.Inst_frame1_bit13.Q
rlabel metal1 10396 2822 10396 2822 0 Inst_S_EF_ADC12_ConfigMem.Inst_frame1_bit14.Q
rlabel metal1 5014 5100 5014 5100 0 Inst_S_EF_ADC12_ConfigMem.Inst_frame1_bit15.Q
rlabel metal2 17342 6358 17342 6358 0 Inst_S_EF_ADC12_ConfigMem.Inst_frame1_bit16.Q
rlabel metal2 28290 3876 28290 3876 0 Inst_S_EF_ADC12_ConfigMem.Inst_frame1_bit17.Q
rlabel metal1 19090 4080 19090 4080 0 Inst_S_EF_ADC12_ConfigMem.Inst_frame1_bit18.Q
rlabel via2 7774 4709 7774 4709 0 Inst_S_EF_ADC12_ConfigMem.Inst_frame1_bit19.Q
rlabel metal1 18124 2618 18124 2618 0 Inst_S_EF_ADC12_ConfigMem.Inst_frame1_bit2.Q
rlabel metal1 22356 6834 22356 6834 0 Inst_S_EF_ADC12_ConfigMem.Inst_frame1_bit20.Q
rlabel metal1 27232 4794 27232 4794 0 Inst_S_EF_ADC12_ConfigMem.Inst_frame1_bit21.Q
rlabel metal1 16974 2992 16974 2992 0 Inst_S_EF_ADC12_ConfigMem.Inst_frame1_bit22.Q
rlabel metal1 9522 3604 9522 3604 0 Inst_S_EF_ADC12_ConfigMem.Inst_frame1_bit23.Q
rlabel metal1 24610 8364 24610 8364 0 Inst_S_EF_ADC12_ConfigMem.Inst_frame1_bit24.Q
rlabel metal1 21252 2482 21252 2482 0 Inst_S_EF_ADC12_ConfigMem.Inst_frame1_bit25.Q
rlabel metal1 33120 2822 33120 2822 0 Inst_S_EF_ADC12_ConfigMem.Inst_frame1_bit26.Q
rlabel metal1 36570 4012 36570 4012 0 Inst_S_EF_ADC12_ConfigMem.Inst_frame1_bit27.Q
rlabel metal1 36662 6188 36662 6188 0 Inst_S_EF_ADC12_ConfigMem.Inst_frame1_bit28.Q
rlabel metal1 35098 2924 35098 2924 0 Inst_S_EF_ADC12_ConfigMem.Inst_frame1_bit29.Q
rlabel metal2 18814 3111 18814 3111 0 Inst_S_EF_ADC12_ConfigMem.Inst_frame1_bit3.Q
rlabel metal2 33534 4828 33534 4828 0 Inst_S_EF_ADC12_ConfigMem.Inst_frame1_bit30.Q
rlabel metal1 33994 6188 33994 6188 0 Inst_S_EF_ADC12_ConfigMem.Inst_frame1_bit31.Q
rlabel metal1 4922 4012 4922 4012 0 Inst_S_EF_ADC12_ConfigMem.Inst_frame1_bit4.Q
rlabel metal2 5474 4148 5474 4148 0 Inst_S_EF_ADC12_ConfigMem.Inst_frame1_bit5.Q
rlabel metal2 21574 4828 21574 4828 0 Inst_S_EF_ADC12_ConfigMem.Inst_frame1_bit6.Q
rlabel metal1 22218 4658 22218 4658 0 Inst_S_EF_ADC12_ConfigMem.Inst_frame1_bit7.Q
rlabel metal2 27922 5015 27922 5015 0 Inst_S_EF_ADC12_ConfigMem.Inst_frame1_bit8.Q
rlabel metal1 28152 3366 28152 3366 0 Inst_S_EF_ADC12_ConfigMem.Inst_frame1_bit9.Q
rlabel metal1 31004 6834 31004 6834 0 Inst_S_EF_ADC12_ConfigMem.Inst_frame2_bit30.Q
rlabel metal2 31418 6630 31418 6630 0 Inst_S_EF_ADC12_ConfigMem.Inst_frame2_bit31.Q
rlabel metal2 19458 2618 19458 2618 0 Inst_S_EF_ADC12_switch_matrix.N1BEG0
rlabel metal1 5566 4114 5566 4114 0 Inst_S_EF_ADC12_switch_matrix.N1BEG1
rlabel metal1 22954 4794 22954 4794 0 Inst_S_EF_ADC12_switch_matrix.N1BEG2
rlabel metal2 29118 5508 29118 5508 0 Inst_S_EF_ADC12_switch_matrix.N1BEG3
rlabel metal1 13340 2618 13340 2618 0 Inst_S_EF_ADC12_switch_matrix.N2BEG0
rlabel metal1 3266 5236 3266 5236 0 Inst_S_EF_ADC12_switch_matrix.N2BEG1
rlabel metal1 2346 7412 2346 7412 0 Inst_S_EF_ADC12_switch_matrix.N2BEG2
rlabel metal1 10672 2414 10672 2414 0 Inst_S_EF_ADC12_switch_matrix.N2BEG3
rlabel metal1 13938 3536 13938 3536 0 Inst_S_EF_ADC12_switch_matrix.N2BEG4
rlabel metal2 5566 4250 5566 4250 0 Inst_S_EF_ADC12_switch_matrix.N2BEG5
rlabel metal1 18446 4590 18446 4590 0 Inst_S_EF_ADC12_switch_matrix.N2BEG6
rlabel metal1 27554 4080 27554 4080 0 Inst_S_EF_ADC12_switch_matrix.N2BEG7
rlabel metal2 18814 3706 18814 3706 0 Inst_S_EF_ADC12_switch_matrix.N2BEGb0
rlabel metal2 24426 4284 24426 4284 0 Inst_S_EF_ADC12_switch_matrix.N2BEGb1
rlabel metal1 23138 6766 23138 6766 0 Inst_S_EF_ADC12_switch_matrix.N2BEGb2
rlabel metal1 27278 5202 27278 5202 0 Inst_S_EF_ADC12_switch_matrix.N2BEGb3
rlabel metal1 17618 2414 17618 2414 0 Inst_S_EF_ADC12_switch_matrix.N2BEGb4
rlabel metal1 8694 3706 8694 3706 0 Inst_S_EF_ADC12_switch_matrix.N2BEGb5
rlabel metal2 25254 7310 25254 7310 0 Inst_S_EF_ADC12_switch_matrix.N2BEGb6
rlabel metal1 21482 2618 21482 2618 0 Inst_S_EF_ADC12_switch_matrix.N2BEGb7
rlabel metal1 32430 2618 32430 2618 0 Inst_S_EF_ADC12_switch_matrix.N4BEG0
rlabel metal1 35972 3502 35972 3502 0 Inst_S_EF_ADC12_switch_matrix.N4BEG1
rlabel metal1 3542 4590 3542 4590 0 Inst_S_EF_ADC12_switch_matrix.N4BEG10
rlabel metal1 6302 2822 6302 2822 0 Inst_S_EF_ADC12_switch_matrix.N4BEG11
rlabel metal1 20654 3978 20654 3978 0 Inst_S_EF_ADC12_switch_matrix.N4BEG12
rlabel metal1 21712 5338 21712 5338 0 Inst_S_EF_ADC12_switch_matrix.N4BEG13
rlabel metal2 27094 6970 27094 6970 0 Inst_S_EF_ADC12_switch_matrix.N4BEG14
rlabel metal1 26910 2618 26910 2618 0 Inst_S_EF_ADC12_switch_matrix.N4BEG15
rlabel metal2 36110 6596 36110 6596 0 Inst_S_EF_ADC12_switch_matrix.N4BEG2
rlabel metal1 34454 2414 34454 2414 0 Inst_S_EF_ADC12_switch_matrix.N4BEG3
rlabel metal1 32936 4114 32936 4114 0 Inst_S_EF_ADC12_switch_matrix.N4BEG4
rlabel metal2 33442 5882 33442 5882 0 Inst_S_EF_ADC12_switch_matrix.N4BEG5
rlabel metal2 5198 4828 5198 4828 0 Inst_S_EF_ADC12_switch_matrix.N4BEG6
rlabel metal2 18538 4522 18538 4522 0 Inst_S_EF_ADC12_switch_matrix.N4BEG7
rlabel metal1 23184 2414 23184 2414 0 Inst_S_EF_ADC12_switch_matrix.N4BEG8
rlabel metal1 15870 4080 15870 4080 0 Inst_S_EF_ADC12_switch_matrix.N4BEG9
rlabel metal1 15824 2618 15824 2618 0 Inst_S_EF_ADC12_switch_matrix.NN4BEG0
rlabel metal2 2714 7990 2714 7990 0 Inst_S_EF_ADC12_switch_matrix.NN4BEG1
rlabel metal2 34546 7174 34546 7174 0 Inst_S_EF_ADC12_switch_matrix.NN4BEG10
rlabel metal2 32430 4284 32430 4284 0 Inst_S_EF_ADC12_switch_matrix.NN4BEG11
rlabel metal1 23874 4114 23874 4114 0 Inst_S_EF_ADC12_switch_matrix.NN4BEG12
rlabel metal1 24748 3502 24748 3502 0 Inst_S_EF_ADC12_switch_matrix.NN4BEG13
rlabel metal1 24334 5678 24334 5678 0 Inst_S_EF_ADC12_switch_matrix.NN4BEG14
rlabel metal2 25530 3468 25530 3468 0 Inst_S_EF_ADC12_switch_matrix.NN4BEG15
rlabel metal2 1426 8704 1426 8704 0 Inst_S_EF_ADC12_switch_matrix.NN4BEG2
rlabel metal2 11730 3468 11730 3468 0 Inst_S_EF_ADC12_switch_matrix.NN4BEG3
rlabel metal1 9752 2278 9752 2278 0 Inst_S_EF_ADC12_switch_matrix.NN4BEG4
rlabel metal2 2898 5338 2898 5338 0 Inst_S_EF_ADC12_switch_matrix.NN4BEG5
rlabel metal2 5290 5372 5290 5372 0 Inst_S_EF_ADC12_switch_matrix.NN4BEG6
rlabel metal1 30452 3026 30452 3026 0 Inst_S_EF_ADC12_switch_matrix.NN4BEG7
rlabel metal2 19090 4250 19090 4250 0 Inst_S_EF_ADC12_switch_matrix.NN4BEG8
rlabel metal1 7084 4250 7084 4250 0 Inst_S_EF_ADC12_switch_matrix.NN4BEG9
rlabel metal2 3266 11145 3266 11145 0 N1BEG[0]
rlabel metal1 1564 6426 1564 6426 0 N1BEG[1]
rlabel metal1 3634 6630 3634 6630 0 N1BEG[2]
rlabel metal1 4232 5882 4232 5882 0 N1BEG[3]
rlabel metal2 1794 8194 1794 8194 0 N2BEG[0]
rlabel metal1 4048 9690 4048 9690 0 N2BEG[1]
rlabel metal1 4002 8058 4002 8058 0 N2BEG[2]
rlabel metal1 4508 5814 4508 5814 0 N2BEG[3]
rlabel metal1 3220 6630 3220 6630 0 N2BEG[4]
rlabel metal1 5980 3978 5980 3978 0 N2BEG[5]
rlabel metal1 3220 6970 3220 6970 0 N2BEG[6]
rlabel metal1 6164 5338 6164 5338 0 N2BEG[7]
rlabel metal1 3910 6086 3910 6086 0 N2BEGb[0]
rlabel metal1 6900 5882 6900 5882 0 N2BEGb[1]
rlabel metal1 7176 6426 7176 6426 0 N2BEGb[2]
rlabel metal1 7498 5882 7498 5882 0 N2BEGb[3]
rlabel metal2 2714 7463 2714 7463 0 N2BEGb[4]
rlabel metal1 6118 6426 6118 6426 0 N2BEGb[5]
rlabel metal1 4508 6154 4508 6154 0 N2BEGb[6]
rlabel metal2 8510 10433 8510 10433 0 N2BEGb[7]
rlabel metal2 6486 8296 6486 8296 0 N4BEG[0]
rlabel metal1 5198 8364 5198 8364 0 N4BEG[10]
rlabel metal2 6118 9248 6118 9248 0 N4BEG[11]
rlabel metal1 7176 8602 7176 8602 0 N4BEG[12]
rlabel metal1 10488 9758 10488 9758 0 N4BEG[13]
rlabel metal2 12650 10550 12650 10550 0 N4BEG[14]
rlabel via1 12926 11196 12926 11196 0 N4BEG[15]
rlabel metal2 8970 10404 8970 10404 0 N4BEG[1]
rlabel metal2 5198 6681 5198 6681 0 N4BEG[2]
rlabel metal1 8004 5882 8004 5882 0 N4BEG[3]
rlabel metal2 7590 8143 7590 8143 0 N4BEG[4]
rlabel metal2 3542 8823 3542 8823 0 N4BEG[5]
rlabel metal1 4784 6630 4784 6630 0 N4BEG[6]
rlabel metal2 5014 9027 5014 9027 0 N4BEG[7]
rlabel metal1 5796 8602 5796 8602 0 N4BEG[8]
rlabel metal3 10350 10268 10350 10268 0 N4BEG[9]
rlabel metal2 13202 10465 13202 10465 0 NN4BEG[0]
rlabel metal1 15226 8568 15226 8568 0 NN4BEG[10]
rlabel metal1 15916 8602 15916 8602 0 NN4BEG[11]
rlabel metal1 16008 8330 16008 8330 0 NN4BEG[12]
rlabel metal1 16560 8602 16560 8602 0 NN4BEG[13]
rlabel metal1 17572 8602 17572 8602 0 NN4BEG[14]
rlabel metal1 17802 8058 17802 8058 0 NN4BEG[15]
rlabel metal3 14812 10268 14812 10268 0 NN4BEG[1]
rlabel metal2 13754 10584 13754 10584 0 NN4BEG[2]
rlabel metal2 14030 10516 14030 10516 0 NN4BEG[3]
rlabel metal1 13984 7242 13984 7242 0 NN4BEG[4]
rlabel metal2 14582 10958 14582 10958 0 NN4BEG[5]
rlabel metal2 14858 10601 14858 10601 0 NN4BEG[6]
rlabel metal1 14030 8602 14030 8602 0 NN4BEG[7]
rlabel metal1 13386 8364 13386 8364 0 NN4BEG[8]
rlabel metal1 14766 8330 14766 8330 0 NN4BEG[9]
rlabel metal2 3358 599 3358 599 0 RESET_top
rlabel metal2 17894 9853 17894 9853 0 S1END[0]
rlabel metal3 18331 8092 18331 8092 0 S1END[1]
rlabel metal2 18446 11026 18446 11026 0 S1END[2]
rlabel via3 18699 8636 18699 8636 0 S1END[3]
rlabel metal2 21206 10533 21206 10533 0 S2END[0]
rlabel metal2 21482 9836 21482 9836 0 S2END[1]
rlabel metal2 21758 9768 21758 9768 0 S2END[2]
rlabel metal1 22264 6902 22264 6902 0 S2END[3]
rlabel metal1 22954 6970 22954 6970 0 S2END[4]
rlabel metal2 22586 10465 22586 10465 0 S2END[5]
rlabel metal2 22862 10533 22862 10533 0 S2END[6]
rlabel metal2 23138 10261 23138 10261 0 S2END[7]
rlabel metal2 18998 10516 18998 10516 0 S2MID[0]
rlabel metal2 19274 8748 19274 8748 0 S2MID[1]
rlabel metal2 19550 10465 19550 10465 0 S2MID[2]
rlabel metal2 19826 10261 19826 10261 0 S2MID[3]
rlabel metal2 20102 9836 20102 9836 0 S2MID[4]
rlabel metal2 20378 10125 20378 10125 0 S2MID[5]
rlabel metal2 20654 8748 20654 8748 0 S2MID[6]
rlabel metal2 20930 10652 20930 10652 0 S2MID[7]
rlabel metal2 23414 10669 23414 10669 0 S4END[0]
rlabel metal1 29026 7820 29026 7820 0 S4END[10]
rlabel metal2 26450 10669 26450 10669 0 S4END[11]
rlabel metal2 26726 9088 26726 9088 0 S4END[12]
rlabel metal2 27002 10737 27002 10737 0 S4END[13]
rlabel metal2 27278 10533 27278 10533 0 S4END[14]
rlabel metal2 27554 10040 27554 10040 0 S4END[15]
rlabel metal1 25070 9418 25070 9418 0 S4END[1]
rlabel metal2 23966 9445 23966 9445 0 S4END[2]
rlabel metal2 24288 7990 24288 7990 0 S4END[3]
rlabel metal2 24518 10601 24518 10601 0 S4END[4]
rlabel metal1 25254 8262 25254 8262 0 S4END[5]
rlabel metal2 25070 9632 25070 9632 0 S4END[6]
rlabel metal2 25346 10006 25346 10006 0 S4END[7]
rlabel metal2 25622 10040 25622 10040 0 S4END[8]
rlabel metal2 25898 10465 25898 10465 0 S4END[9]
rlabel metal2 32338 8874 32338 8874 0 SS4END[0]
rlabel metal2 34086 9180 34086 9180 0 SS4END[10]
rlabel via2 32062 6749 32062 6749 0 SS4END[11]
rlabel metal2 33534 8857 33534 8857 0 SS4END[12]
rlabel metal1 32016 9350 32016 9350 0 SS4END[13]
rlabel metal2 33718 8755 33718 8755 0 SS4END[14]
rlabel metal2 31970 10210 31970 10210 0 SS4END[15]
rlabel via3 28083 8636 28083 8636 0 SS4END[1]
rlabel metal2 28382 10737 28382 10737 0 SS4END[2]
rlabel metal2 28658 8952 28658 8952 0 SS4END[3]
rlabel metal2 32430 9401 32430 9401 0 SS4END[4]
rlabel metal2 29210 9836 29210 9836 0 SS4END[5]
rlabel metal2 32246 7565 32246 7565 0 SS4END[6]
rlabel metal1 30682 9214 30682 9214 0 SS4END[7]
rlabel metal2 31786 6443 31786 6443 0 SS4END[8]
rlabel metal2 32890 7616 32890 7616 0 SS4END[9]
rlabel metal1 19596 4182 19596 4182 0 UserCLK
rlabel metal1 18722 6358 18722 6358 0 UserCLK_regs
rlabel metal1 34454 7174 34454 7174 0 UserCLKo
rlabel metal2 4462 1160 4462 1160 0 VALUE_top0
rlabel metal2 5566 1160 5566 1160 0 VALUE_top1
rlabel metal2 15502 1160 15502 1160 0 VALUE_top10
rlabel metal2 16606 1160 16606 1160 0 VALUE_top11
rlabel metal2 6670 1160 6670 1160 0 VALUE_top2
rlabel metal2 7774 1160 7774 1160 0 VALUE_top3
rlabel metal2 8878 55 8878 55 0 VALUE_top4
rlabel metal2 9982 1160 9982 1160 0 VALUE_top5
rlabel metal2 11086 1160 11086 1160 0 VALUE_top6
rlabel metal2 12466 1153 12466 1153 0 VALUE_top7
rlabel metal2 13294 1840 13294 1840 0 VALUE_top8
rlabel metal2 14398 1160 14398 1160 0 VALUE_top9
rlabel metal1 21753 7446 21753 7446 0 _000_
rlabel metal1 17332 7378 17332 7378 0 _001_
rlabel metal2 22586 6970 22586 6970 0 _002_
rlabel via1 19085 7378 19085 7378 0 _003_
rlabel metal1 17622 7854 17622 7854 0 _004_
rlabel metal1 23556 7446 23556 7446 0 _005_
rlabel metal1 16330 6222 16330 6222 0 _006_
rlabel metal1 19448 5678 19448 5678 0 _007_
rlabel metal1 16003 4522 16003 4522 0 _008_
rlabel metal2 15594 6086 15594 6086 0 _009_
rlabel metal1 8004 4794 8004 4794 0 _010_
rlabel via1 12185 3434 12185 3434 0 _011_
rlabel metal2 11086 7378 11086 7378 0 _012_
rlabel viali 9231 7854 9231 7854 0 _013_
rlabel metal1 8234 6358 8234 6358 0 _014_
rlabel metal1 9885 4522 9885 4522 0 _015_
rlabel metal1 12047 4522 12047 4522 0 _016_
rlabel via1 12645 7854 12645 7854 0 _017_
rlabel metal1 15210 7786 15210 7786 0 _018_
rlabel metal1 32062 7310 32062 7310 0 _019_
rlabel metal1 31505 7446 31505 7446 0 _020_
rlabel metal1 28929 7446 28929 7446 0 _021_
rlabel metal1 28147 6766 28147 6766 0 _022_
rlabel via1 15690 5270 15690 5270 0 _023_
rlabel metal1 15962 5712 15962 5712 0 _024_
rlabel metal1 8510 4624 8510 4624 0 _025_
rlabel metal2 11362 5168 11362 5168 0 _026_
rlabel metal2 10718 6596 10718 6596 0 _027_
rlabel metal2 8418 7650 8418 7650 0 _028_
rlabel metal2 8694 6494 8694 6494 0 _029_
rlabel metal1 9046 5610 9046 5610 0 _030_
rlabel via1 11909 6290 11909 6290 0 _031_
rlabel metal1 13068 7446 13068 7446 0 _032_
rlabel metal1 14674 7888 14674 7888 0 _033_
rlabel via1 18745 5338 18745 5338 0 _034_
rlabel metal2 18906 7973 18906 7973 0 _035_
rlabel metal1 14260 7854 14260 7854 0 _036_
rlabel metal1 29946 7446 29946 7446 0 _037_
rlabel metal1 21620 3978 21620 3978 0 _038_
rlabel metal2 21482 5406 21482 5406 0 _039_
rlabel metal1 23460 4794 23460 4794 0 _040_
rlabel metal1 23506 5134 23506 5134 0 _041_
rlabel metal2 23138 6052 23138 6052 0 _042_
rlabel metal2 23046 5423 23046 5423 0 _043_
rlabel metal1 18814 8364 18814 8364 0 _044_
rlabel metal1 28566 3944 28566 3944 0 _045_
rlabel metal1 28612 4046 28612 4046 0 _046_
rlabel metal1 26956 3706 26956 3706 0 _047_
rlabel metal2 29210 5576 29210 5576 0 _048_
rlabel metal1 29118 4794 29118 4794 0 _049_
rlabel metal2 18998 8670 18998 8670 0 _050_
rlabel metal2 10902 5950 10902 5950 0 _051_
rlabel metal1 10856 6426 10856 6426 0 _052_
rlabel metal1 15778 3910 15778 3910 0 _053_
rlabel metal1 17401 7514 17401 7514 0 _054_
rlabel metal2 31050 7616 31050 7616 0 _055_
rlabel metal2 30038 7956 30038 7956 0 _056_
rlabel metal1 29808 5814 29808 5814 0 _057_
rlabel metal1 30912 6630 30912 6630 0 _058_
rlabel metal1 24058 8398 24058 8398 0 _059_
rlabel metal1 23092 8330 23092 8330 0 _060_
rlabel metal2 16422 7378 16422 7378 0 _061_
rlabel metal2 15870 7582 15870 7582 0 _062_
rlabel metal1 1978 8500 1978 8500 0 _063_
rlabel metal1 13340 4250 13340 4250 0 _064_
rlabel metal1 16790 5576 16790 5576 0 _065_
rlabel metal2 16146 4148 16146 4148 0 _066_
rlabel metal1 8740 4250 8740 4250 0 _067_
rlabel metal2 11638 4692 11638 4692 0 _068_
rlabel metal1 2415 8330 2415 8330 0 _069_
rlabel metal1 8234 7922 8234 7922 0 _070_
rlabel metal2 8694 3978 8694 3978 0 _071_
rlabel metal1 9154 4012 9154 4012 0 _072_
rlabel metal2 9982 4335 9982 4335 0 _073_
rlabel metal1 10718 3910 10718 3910 0 _074_
rlabel metal1 14398 7820 14398 7820 0 _075_
rlabel metal1 33304 7854 33304 7854 0 _076_
rlabel metal1 29670 8058 29670 8058 0 _077_
rlabel metal2 30222 7412 30222 7412 0 _078_
rlabel metal1 28106 8262 28106 8262 0 _079_
rlabel metal2 28934 8279 28934 8279 0 _080_
rlabel metal2 26266 7616 26266 7616 0 clknet_0_UserCLK
rlabel metal1 22310 6766 22310 6766 0 clknet_0_UserCLK_regs
rlabel metal1 27646 8500 27646 8500 0 clknet_1_0__leaf_UserCLK
rlabel metal2 14766 4930 14766 4930 0 clknet_2_0__leaf_UserCLK_regs
rlabel metal2 8372 8398 8372 8398 0 clknet_2_1__leaf_UserCLK_regs
rlabel metal2 24150 7616 24150 7616 0 clknet_2_2__leaf_UserCLK_regs
rlabel metal1 15272 7378 15272 7378 0 clknet_2_3__leaf_UserCLK_regs
rlabel metal2 7682 1938 7682 1938 0 net1
rlabel metal2 3542 1907 3542 1907 0 net10
rlabel metal1 39422 4114 39422 4114 0 net100
rlabel metal3 2369 6324 2369 6324 0 net101
rlabel metal1 39422 4454 39422 4454 0 net102
rlabel metal1 36386 5134 36386 5134 0 net103
rlabel metal1 31878 5032 31878 5032 0 net104
rlabel metal2 39836 4284 39836 4284 0 net105
rlabel metal2 16514 3213 16514 3213 0 net106
rlabel metal1 32430 3672 32430 3672 0 net107
rlabel metal2 17158 2584 17158 2584 0 net108
rlabel metal1 38778 6154 38778 6154 0 net109
rlabel metal1 2622 3910 2622 3910 0 net11
rlabel metal2 34638 2210 34638 2210 0 net110
rlabel metal1 26496 6426 26496 6426 0 net111
rlabel metal2 35834 5610 35834 5610 0 net112
rlabel metal4 32660 7820 32660 7820 0 net113
rlabel metal1 17158 9384 17158 9384 0 net114
rlabel metal2 38594 8908 38594 8908 0 net115
rlabel metal2 38870 8415 38870 8415 0 net116
rlabel metal1 33902 2414 33902 2414 0 net117
rlabel metal2 36018 5984 36018 5984 0 net118
rlabel metal1 39238 6732 39238 6732 0 net119
rlabel metal1 5980 5678 5980 5678 0 net12
rlabel metal1 36018 2618 36018 2618 0 net120
rlabel metal2 21666 2924 21666 2924 0 net121
rlabel metal1 34454 5882 34454 5882 0 net122
rlabel metal1 32476 5542 32476 5542 0 net123
rlabel metal2 38870 1802 38870 1802 0 net124
rlabel metal2 37490 2210 37490 2210 0 net125
rlabel metal2 17894 1887 17894 1887 0 net126
rlabel metal1 19964 4454 19964 4454 0 net127
rlabel metal2 19366 5151 19366 5151 0 net128
rlabel metal2 37306 3791 37306 3791 0 net129
rlabel metal2 1610 2176 1610 2176 0 net13
rlabel metal2 38870 3876 38870 3876 0 net130
rlabel metal1 30912 2618 30912 2618 0 net131
rlabel metal1 37260 6630 37260 6630 0 net132
rlabel metal1 37490 5814 37490 5814 0 net133
rlabel metal1 37168 5882 37168 5882 0 net134
rlabel metal1 36984 7514 36984 7514 0 net135
rlabel metal1 35650 2890 35650 2890 0 net136
rlabel metal1 37214 4794 37214 4794 0 net137
rlabel metal1 38042 4794 38042 4794 0 net138
rlabel metal1 37904 5882 37904 5882 0 net139
rlabel metal1 2300 5882 2300 5882 0 net14
rlabel metal1 38686 5338 38686 5338 0 net140
rlabel metal1 37122 3162 37122 3162 0 net141
rlabel metal2 25990 2873 25990 2873 0 net142
rlabel metal2 33074 8262 33074 8262 0 net143
rlabel metal1 36662 2822 36662 2822 0 net144
rlabel metal1 36938 5338 36938 5338 0 net145
rlabel metal1 37490 5542 37490 5542 0 net146
rlabel metal1 38364 5338 38364 5338 0 net147
rlabel metal1 37996 6154 37996 6154 0 net148
rlabel metal1 37444 3978 37444 3978 0 net149
rlabel metal1 1564 4794 1564 4794 0 net15
rlabel metal1 38226 6868 38226 6868 0 net150
rlabel metal2 2622 1513 2622 1513 0 net151
rlabel metal2 19274 2329 19274 2329 0 net152
rlabel metal1 4968 4250 4968 4250 0 net153
rlabel metal3 22701 5644 22701 5644 0 net154
rlabel metal1 4646 2482 4646 2482 0 net155
rlabel metal1 2346 6732 2346 6732 0 net156
rlabel metal1 2944 5338 2944 5338 0 net157
rlabel metal2 2530 7650 2530 7650 0 net158
rlabel metal1 9016 2618 9016 2618 0 net159
rlabel metal1 1702 2618 1702 2618 0 net16
rlabel metal2 4922 4828 4922 4828 0 net160
rlabel metal1 5796 3706 5796 3706 0 net161
rlabel metal2 1518 1703 1518 1703 0 net162
rlabel metal3 16560 1632 16560 1632 0 net163
rlabel metal2 4508 2380 4508 2380 0 net164
rlabel metal1 15640 578 15640 578 0 net165
rlabel metal2 7314 8330 7314 8330 0 net166
rlabel metal1 26864 5338 26864 5338 0 net167
rlabel metal2 17526 1853 17526 1853 0 net168
rlabel metal1 7866 3978 7866 3978 0 net169
rlabel metal2 23506 2176 23506 2176 0 net17
rlabel metal2 17434 10064 17434 10064 0 net170
rlabel metal1 20240 3366 20240 3366 0 net171
rlabel metal2 13294 7123 13294 7123 0 net172
rlabel metal1 4140 4794 4140 4794 0 net173
rlabel metal1 5980 8466 5980 8466 0 net174
rlabel metal1 20608 4454 20608 4454 0 net175
rlabel metal1 21436 6086 21436 6086 0 net176
rlabel metal4 7820 9112 7820 9112 0 net177
rlabel metal1 17066 9962 17066 9962 0 net178
rlabel metal2 35834 2125 35834 2125 0 net179
rlabel via2 2622 7837 2622 7837 0 net18
rlabel metal2 17158 9996 17158 9996 0 net180
rlabel metal2 33442 2006 33442 2006 0 net181
rlabel metal2 32798 3553 32798 3553 0 net182
rlabel metal1 12466 9690 12466 9690 0 net183
rlabel metal2 5014 5372 5014 5372 0 net184
rlabel metal1 5980 7174 5980 7174 0 net185
rlabel metal2 16882 9180 16882 9180 0 net186
rlabel metal2 7038 7701 7038 7701 0 net187
rlabel metal2 15686 3553 15686 3553 0 net188
rlabel metal2 15594 8891 15594 8891 0 net189
rlabel metal2 2530 8823 2530 8823 0 net19
rlabel metal2 15778 8959 15778 8959 0 net190
rlabel metal1 19182 8296 19182 8296 0 net191
rlabel metal2 17526 8976 17526 8976 0 net192
rlabel metal2 18262 8704 18262 8704 0 net193
rlabel metal1 18446 7922 18446 7922 0 net194
rlabel metal2 2714 4318 2714 4318 0 net195
rlabel metal2 1610 8738 1610 8738 0 net196
rlabel metal1 11684 3162 11684 3162 0 net197
rlabel metal2 9982 3315 9982 3315 0 net198
rlabel metal2 10350 8908 10350 8908 0 net199
rlabel metal1 3358 2618 3358 2618 0 net2
rlabel via2 1794 5083 1794 5083 0 net20
rlabel metal1 5336 3910 5336 3910 0 net200
rlabel metal1 12880 8466 12880 8466 0 net201
rlabel metal1 18814 3366 18814 3366 0 net202
rlabel metal1 13662 8500 13662 8500 0 net203
rlabel metal1 19918 7718 19918 7718 0 net204
rlabel metal1 28060 8602 28060 8602 0 net205
rlabel metal2 16698 4420 16698 4420 0 net206
rlabel metal1 14720 6086 14720 6086 0 net207
rlabel metal1 4554 8364 4554 8364 0 net208
rlabel metal1 16974 2448 16974 2448 0 net209
rlabel via2 2070 4539 2070 4539 0 net21
rlabel metal1 5290 5270 5290 5270 0 net210
rlabel metal1 8050 2482 8050 2482 0 net211
rlabel metal1 8970 2448 8970 2448 0 net212
rlabel metal1 6808 6834 6808 6834 0 net213
rlabel metal1 9476 3366 9476 3366 0 net214
rlabel metal1 14260 2346 14260 2346 0 net215
rlabel metal1 20838 4046 20838 4046 0 net216
rlabel metal2 7774 7344 7774 7344 0 net217
rlabel metal1 16928 6834 16928 6834 0 net218
rlabel metal1 22724 8398 22724 8398 0 net219
rlabel metal1 2254 5814 2254 5814 0 net22
rlabel metal2 13570 5100 13570 5100 0 net220
rlabel metal1 17894 8500 17894 8500 0 net221
rlabel metal2 14766 8585 14766 8585 0 net222
rlabel metal2 13294 4386 13294 4386 0 net223
rlabel metal2 13110 5916 13110 5916 0 net224
rlabel metal2 8326 5882 8326 5882 0 net225
rlabel metal1 14490 4624 14490 4624 0 net226
rlabel via2 16054 4131 16054 4131 0 net227
rlabel metal2 9706 8823 9706 8823 0 net228
rlabel metal2 2162 8840 2162 8840 0 net229
rlabel metal2 12558 2907 12558 2907 0 net23
rlabel metal1 22908 7514 22908 7514 0 net230
rlabel metal2 9522 6766 9522 6766 0 net231
rlabel metal1 10902 6630 10902 6630 0 net232
rlabel metal1 10902 4998 10902 4998 0 net233
rlabel metal2 16882 5763 16882 5763 0 net234
rlabel metal1 18934 5202 18934 5202 0 net235
rlabel metal1 18814 6256 18814 6256 0 net236
rlabel metal1 33074 7922 33074 7922 0 net237
rlabel metal1 20838 3060 20838 3060 0 net24
rlabel via2 2162 6205 2162 6205 0 net25
rlabel via2 2530 5661 2530 5661 0 net26
rlabel metal2 2898 2142 2898 2142 0 net27
rlabel metal1 2990 4114 2990 4114 0 net28
rlabel metal1 3220 3094 3220 3094 0 net29
rlabel metal1 9062 3060 9062 3060 0 net3
rlabel metal1 19274 4556 19274 4556 0 net30
rlabel metal3 9476 3400 9476 3400 0 net31
rlabel metal2 2806 3723 2806 3723 0 net32
rlabel metal2 1702 8976 1702 8976 0 net33
rlabel metal2 8142 7548 8142 7548 0 net34
rlabel metal1 7866 6324 7866 6324 0 net35
rlabel metal1 6302 7310 6302 7310 0 net36
rlabel metal1 20424 3026 20424 3026 0 net37
rlabel metal1 19780 3026 19780 3026 0 net38
rlabel metal2 19274 3808 19274 3808 0 net39
rlabel metal1 1932 6698 1932 6698 0 net4
rlabel metal2 2714 3842 2714 3842 0 net40
rlabel metal2 14030 3009 14030 3009 0 net41
rlabel metal1 31924 2958 31924 2958 0 net42
rlabel metal2 34822 5644 34822 5644 0 net43
rlabel metal2 9798 3791 9798 3791 0 net44
rlabel metal1 32062 5202 32062 5202 0 net45
rlabel metal2 25898 1938 25898 1938 0 net46
rlabel metal1 17664 5882 17664 5882 0 net47
rlabel metal1 21114 4726 21114 4726 0 net48
rlabel metal1 17112 6630 17112 6630 0 net49
rlabel metal1 3082 6358 3082 6358 0 net5
rlabel metal2 17802 4284 17802 4284 0 net50
rlabel metal1 21390 2278 21390 2278 0 net51
rlabel metal1 24472 8602 24472 8602 0 net52
rlabel metal2 18354 8687 18354 8687 0 net53
rlabel metal2 23874 5032 23874 5032 0 net54
rlabel metal1 27278 5610 27278 5610 0 net55
rlabel metal2 22678 6494 22678 6494 0 net56
rlabel metal1 25254 5338 25254 5338 0 net57
rlabel metal2 22218 4743 22218 4743 0 net58
rlabel metal2 17526 5117 17526 5117 0 net59
rlabel metal1 10442 3502 10442 3502 0 net6
rlabel metal1 19044 6086 19044 6086 0 net60
rlabel metal1 7406 5202 7406 5202 0 net61
rlabel metal1 20792 5746 20792 5746 0 net62
rlabel metal3 14444 2584 14444 2584 0 net63
rlabel metal1 5474 7854 5474 7854 0 net64
rlabel via2 19274 6069 19274 6069 0 net65
rlabel metal1 13800 2414 13800 2414 0 net66
rlabel metal1 27600 2414 27600 2414 0 net67
rlabel metal1 32890 6426 32890 6426 0 net68
rlabel metal1 32982 4522 32982 4522 0 net69
rlabel metal1 7912 3026 7912 3026 0 net7
rlabel metal1 32798 2890 32798 2890 0 net70
rlabel metal1 33810 6358 33810 6358 0 net71
rlabel metal1 35696 4182 35696 4182 0 net72
rlabel metal1 32844 2414 32844 2414 0 net73
rlabel metal1 27094 7514 27094 7514 0 net74
rlabel metal1 25070 5100 25070 5100 0 net75
rlabel metal1 22724 4250 22724 4250 0 net76
rlabel metal1 17158 10030 17158 10030 0 net77
rlabel metal3 20516 7140 20516 7140 0 net78
rlabel metal1 14352 4250 14352 4250 0 net79
rlabel metal1 1978 2924 1978 2924 0 net8
rlabel metal2 29854 9078 29854 9078 0 net80
rlabel metal1 18262 5678 18262 5678 0 net81
rlabel metal1 5336 5678 5336 5678 0 net82
rlabel metal2 25438 5491 25438 5491 0 net83
rlabel metal2 16606 7888 16606 7888 0 net84
rlabel metal2 32430 4012 32430 4012 0 net85
rlabel metal2 33626 7769 33626 7769 0 net86
rlabel metal2 14582 7684 14582 7684 0 net87
rlabel metal1 33672 8058 33672 8058 0 net88
rlabel metal1 31878 2346 31878 2346 0 net89
rlabel metal1 2346 2890 2346 2890 0 net9
rlabel metal1 25346 5678 25346 5678 0 net90
rlabel metal2 29578 5984 29578 5984 0 net91
rlabel metal2 29946 5440 29946 5440 0 net92
rlabel metal2 32522 5882 32522 5882 0 net93
rlabel metal1 30590 5882 30590 5882 0 net94
rlabel metal2 32982 7463 32982 7463 0 net95
rlabel metal2 31878 5661 31878 5661 0 net96
rlabel metal1 30038 3162 30038 3162 0 net97
rlabel metal3 14812 7480 14812 7480 0 net98
rlabel metal2 38134 2142 38134 2142 0 net99
<< properties >>
string FIXED_BBOX 0 0 41000 11250
<< end >>
