module LUT4AB (Ci,
    Co,
    UserCLK,
    UserCLKo,
    E1BEG,
    E1END,
    E2BEG,
    E2BEGb,
    E2END,
    E2MID,
    E6BEG,
    E6END,
    EE4BEG,
    EE4END,
    FrameData,
    FrameData_O,
    FrameStrobe,
    FrameStrobe_O,
    N1BEG,
    N1END,
    N2BEG,
    N2BEGb,
    N2END,
    N2MID,
    N4BEG,
    N4END,
    NN4BEG,
    NN4END,
    S1BEG,
    S1END,
    S2BEG,
    S2BEGb,
    S2END,
    S2MID,
    S4BEG,
    S4END,
    SS4BEG,
    SS4END,
    W1BEG,
    W1END,
    W2BEG,
    W2BEGb,
    W2END,
    W2MID,
    W6BEG,
    W6END,
    WW4BEG,
    WW4END);
 input Ci;
 output Co;
 input UserCLK;
 output UserCLKo;
 output [3:0] E1BEG;
 input [3:0] E1END;
 output [7:0] E2BEG;
 output [7:0] E2BEGb;
 input [7:0] E2END;
 input [7:0] E2MID;
 output [11:0] E6BEG;
 input [11:0] E6END;
 output [15:0] EE4BEG;
 input [15:0] EE4END;
 input [31:0] FrameData;
 output [31:0] FrameData_O;
 input [19:0] FrameStrobe;
 output [19:0] FrameStrobe_O;
 output [3:0] N1BEG;
 input [3:0] N1END;
 output [7:0] N2BEG;
 output [7:0] N2BEGb;
 input [7:0] N2END;
 input [7:0] N2MID;
 output [15:0] N4BEG;
 input [15:0] N4END;
 output [15:0] NN4BEG;
 input [15:0] NN4END;
 output [3:0] S1BEG;
 input [3:0] S1END;
 output [7:0] S2BEG;
 output [7:0] S2BEGb;
 input [7:0] S2END;
 input [7:0] S2MID;
 output [15:0] S4BEG;
 input [15:0] S4END;
 output [15:0] SS4BEG;
 input [15:0] SS4END;
 output [3:0] W1BEG;
 input [3:0] W1END;
 output [7:0] W2BEG;
 output [7:0] W2BEGb;
 input [7:0] W2END;
 input [7:0] W2MID;
 output [11:0] W6BEG;
 input [11:0] W6END;
 output [15:0] WW4BEG;
 input [15:0] WW4END;

 wire A;
 wire B;
 wire C;
 wire net139;
 wire D;
 wire E;
 wire net141;
 wire net399;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net447;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net433;
 wire net431;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net486;
 wire net177;
 wire net450;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire F;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire G;
 wire H;
 wire \Inst_LA_LUT4c_frame_config_dffesr.LUT_flop ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.c_I0mux ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.c_out_mux ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.c_reset_value ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.LUT_flop ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.c_I0mux ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.c_out_mux ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.c_reset_value ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.LUT_flop ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.c_I0mux ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.c_out_mux ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.c_reset_value ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.LUT_flop ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.c_I0mux ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.c_out_mux ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.c_reset_value ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.LUT_flop ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.c_I0mux ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.c_out_mux ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.c_reset_value ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.LUT_flop ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.c_I0mux ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.c_out_mux ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.c_reset_value ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.LUT_flop ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.c_I0mux ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.c_out_mux ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.c_reset_value ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.LUT_flop ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.c_I0mux ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.c_out_mux ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.c_reset_value ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit9.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit9.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit9.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit9.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit9.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit9.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit9.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit9.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit9.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit9.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit9.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit9.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit9.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit9.Q ;
 wire \Inst_LUT4AB_switch_matrix.E1BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.E1BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.E1BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.E1BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.E2BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.E2BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.E2BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.E2BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.E2BEG4 ;
 wire \Inst_LUT4AB_switch_matrix.E2BEG5 ;
 wire \Inst_LUT4AB_switch_matrix.E2BEG6 ;
 wire \Inst_LUT4AB_switch_matrix.E2BEG7 ;
 wire \Inst_LUT4AB_switch_matrix.E6BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.E6BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.EE4BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.EE4BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.EE4BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.EE4BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.JN2BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.JN2BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.JN2BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.JN2BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.JN2BEG4 ;
 wire \Inst_LUT4AB_switch_matrix.JN2BEG5 ;
 wire \Inst_LUT4AB_switch_matrix.JN2BEG6 ;
 wire \Inst_LUT4AB_switch_matrix.JN2BEG7 ;
 wire \Inst_LUT4AB_switch_matrix.JS2BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.JS2BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.JS2BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.JS2BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.JS2BEG4 ;
 wire \Inst_LUT4AB_switch_matrix.JS2BEG5 ;
 wire \Inst_LUT4AB_switch_matrix.JS2BEG6 ;
 wire \Inst_LUT4AB_switch_matrix.JS2BEG7 ;
 wire \Inst_LUT4AB_switch_matrix.JW2BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.JW2BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.JW2BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.JW2BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.JW2BEG4 ;
 wire \Inst_LUT4AB_switch_matrix.JW2BEG5 ;
 wire \Inst_LUT4AB_switch_matrix.JW2BEG6 ;
 wire \Inst_LUT4AB_switch_matrix.JW2BEG7 ;
 wire \Inst_LUT4AB_switch_matrix.M_AB ;
 wire \Inst_LUT4AB_switch_matrix.M_AD ;
 wire \Inst_LUT4AB_switch_matrix.M_AH ;
 wire \Inst_LUT4AB_switch_matrix.M_EF ;
 wire \Inst_LUT4AB_switch_matrix.N1BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.N1BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.N1BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.N1BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.N4BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.N4BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.N4BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.N4BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.NN4BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.NN4BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.NN4BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.NN4BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.S1BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.S1BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.S1BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.S1BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.S4BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.S4BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.S4BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.S4BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.SS4BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.SS4BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.SS4BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.SS4BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.W1BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.W1BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.W1BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.W1BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.W6BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.W6BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.WW4BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.WW4BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.WW4BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.WW4BEG3 ;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net482;
 wire net483;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net485;
 wire net281;
 wire net448;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net480;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net484;
 wire net481;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net424;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net467;
 wire net355;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net446;
 wire net451;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net487;
 wire net382;
 wire net449;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire UserCLK_regs;
 wire clknet_0_UserCLK;
 wire clknet_1_0__leaf_UserCLK;
 wire clknet_0_UserCLK_regs;
 wire clknet_1_0__leaf_UserCLK_regs;
 wire clknet_1_1__leaf_UserCLK_regs;
 wire net396;
 wire net397;
 wire net398;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net432;
 wire net452;
 wire net453;
 wire net454;

 sky130_fd_sc_hd__inv_1 _0697_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit9.Q ),
    .Y(_0548_));
 sky130_fd_sc_hd__inv_2 _0698_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit3.Q ),
    .Y(_0549_));
 sky130_fd_sc_hd__inv_1 _0699_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit1.Q ),
    .Y(_0550_));
 sky130_fd_sc_hd__inv_2 _0700_ (.A(\Inst_LA_LUT4c_frame_config_dffesr.c_I0mux ),
    .Y(_0551_));
 sky130_fd_sc_hd__inv_2 _0701_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit8.Q ),
    .Y(_0552_));
 sky130_fd_sc_hd__inv_1 _0702_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit9.Q ),
    .Y(_0553_));
 sky130_fd_sc_hd__inv_2 _0703_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit5.Q ),
    .Y(_0554_));
 sky130_fd_sc_hd__inv_1 _0704_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit0.Q ),
    .Y(_0555_));
 sky130_fd_sc_hd__inv_1 _0705_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit1.Q ),
    .Y(_0556_));
 sky130_fd_sc_hd__inv_1 _0706_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit8.Q ),
    .Y(_0557_));
 sky130_fd_sc_hd__inv_1 _0707_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit9.Q ),
    .Y(_0558_));
 sky130_fd_sc_hd__inv_2 _0708_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit0.Q ),
    .Y(_0559_));
 sky130_fd_sc_hd__inv_1 _0709_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit1.Q ),
    .Y(_0560_));
 sky130_fd_sc_hd__inv_1 _0710_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit9.Q ),
    .Y(_0561_));
 sky130_fd_sc_hd__inv_1 _0711_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit1.Q ),
    .Y(_0562_));
 sky130_fd_sc_hd__inv_1 _0712_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit21.Q ),
    .Y(_0563_));
 sky130_fd_sc_hd__inv_1 _0713_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit5.Q ),
    .Y(_0564_));
 sky130_fd_sc_hd__inv_1 _0714_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit5.Q ),
    .Y(_0565_));
 sky130_fd_sc_hd__inv_1 _0715_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit13.Q ),
    .Y(_0566_));
 sky130_fd_sc_hd__inv_1 _0716_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit13.Q ),
    .Y(_0567_));
 sky130_fd_sc_hd__inv_1 _0717_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit17.Q ),
    .Y(_0568_));
 sky130_fd_sc_hd__inv_1 _0718_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit17.Q ),
    .Y(_0569_));
 sky130_fd_sc_hd__inv_1 _0719_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit17.Q ),
    .Y(_0570_));
 sky130_fd_sc_hd__inv_1 _0720_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit17.Q ),
    .Y(_0571_));
 sky130_fd_sc_hd__inv_1 _0721_ (.A(\Inst_LE_LUT4c_frame_config_dffesr.c_reset_value ),
    .Y(_0572_));
 sky130_fd_sc_hd__inv_1 _0722_ (.A(\Inst_LF_LUT4c_frame_config_dffesr.c_reset_value ),
    .Y(_0573_));
 sky130_fd_sc_hd__inv_1 _0723_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit21.Q ),
    .Y(_0574_));
 sky130_fd_sc_hd__inv_1 _0724_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit21.Q ),
    .Y(_0575_));
 sky130_fd_sc_hd__inv_1 _0725_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit21.Q ),
    .Y(_0576_));
 sky130_fd_sc_hd__inv_1 _0726_ (.A(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ),
    .Y(_0577_));
 sky130_fd_sc_hd__inv_1 _0727_ (.A(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ),
    .Y(_0578_));
 sky130_fd_sc_hd__inv_1 _0728_ (.A(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ),
    .Y(_0579_));
 sky130_fd_sc_hd__inv_1 _0729_ (.A(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ),
    .Y(_0580_));
 sky130_fd_sc_hd__inv_2 _0730_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit9.Q ),
    .Y(_0581_));
 sky130_fd_sc_hd__inv_1 _0731_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit25.Q ),
    .Y(_0582_));
 sky130_fd_sc_hd__inv_1 _0732_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit25.Q ),
    .Y(_0583_));
 sky130_fd_sc_hd__inv_1 _0733_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit25.Q ),
    .Y(_0584_));
 sky130_fd_sc_hd__inv_1 _0734_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit25.Q ),
    .Y(_0585_));
 sky130_fd_sc_hd__inv_1 _0735_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit25.Q ),
    .Y(_0586_));
 sky130_fd_sc_hd__inv_1 _0736_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit28.Q ),
    .Y(_0587_));
 sky130_fd_sc_hd__inv_1 _0737_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit29.Q ),
    .Y(_0588_));
 sky130_fd_sc_hd__inv_1 _0738_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit28.Q ),
    .Y(_0589_));
 sky130_fd_sc_hd__inv_1 _0739_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit29.Q ),
    .Y(_0590_));
 sky130_fd_sc_hd__inv_2 _0740_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit28.Q ),
    .Y(_0591_));
 sky130_fd_sc_hd__inv_1 _0741_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit29.Q ),
    .Y(_0592_));
 sky130_fd_sc_hd__inv_2 _0742_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit28.Q ),
    .Y(_0593_));
 sky130_fd_sc_hd__inv_1 _0743_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit29.Q ),
    .Y(_0594_));
 sky130_fd_sc_hd__inv_1 _0744_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit16.Q ),
    .Y(_0595_));
 sky130_fd_sc_hd__inv_1 _0745_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit28.Q ),
    .Y(_0596_));
 sky130_fd_sc_hd__inv_2 _0746_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit31.Q ),
    .Y(_0597_));
 sky130_fd_sc_hd__mux4_1 _0747_ (.A0(net663),
    .A1(net635),
    .A2(net651),
    .A3(net644),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit31.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit30.Q ),
    .X(_0598_));
 sky130_fd_sc_hd__or2_1 _0748_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit0.Q ),
    .B(_0598_),
    .X(_0599_));
 sky130_fd_sc_hd__mux4_1 _0749_ (.A0(net640),
    .A1(net629),
    .A2(net626),
    .A3(net623),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit30.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit31.Q ),
    .X(_0600_));
 sky130_fd_sc_hd__o21a_1 _0750_ (.A1(_0555_),
    .A2(_0600_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit1.Q ),
    .X(_0601_));
 sky130_fd_sc_hd__mux4_1 _0751_ (.A0(net57),
    .A1(net63),
    .A2(net79),
    .A3(net8),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit30.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit31.Q ),
    .X(_0602_));
 sky130_fd_sc_hd__mux4_1 _0752_ (.A0(net814),
    .A1(net91),
    .A2(net119),
    .A3(net138),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit30.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit31.Q ),
    .X(_0603_));
 sky130_fd_sc_hd__mux2_1 _0753_ (.A0(_0602_),
    .A1(_0603_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit0.Q ),
    .X(_0604_));
 sky130_fd_sc_hd__a22o_1 _0754_ (.A1(_0601_),
    .A2(_0599_),
    .B1(_0604_),
    .B2(_0556_),
    .X(\Inst_LUT4AB_switch_matrix.E2BEG1 ));
 sky130_fd_sc_hd__mux4_1 _0755_ (.A0(net26),
    .A1(net107),
    .A2(net124),
    .A3(\Inst_LUT4AB_switch_matrix.E2BEG1 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit28.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit29.Q ),
    .X(_0605_));
 sky130_fd_sc_hd__mux4_2 _0756_ (.A0(net81),
    .A1(net91),
    .A2(net8),
    .A3(net119),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit29.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit28.Q ),
    .X(_0606_));
 sky130_fd_sc_hd__or2_1 _0757_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit5.Q ),
    .B(_0606_),
    .X(_0607_));
 sky130_fd_sc_hd__o211a_1 _0758_ (.A1(_0554_),
    .A2(_0605_),
    .B1(_0607_),
    .C1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit6.Q ),
    .X(_0608_));
 sky130_fd_sc_hd__mux4_2 _0759_ (.A0(net659),
    .A1(net654),
    .A2(net649),
    .A3(net644),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit7.Q ),
    .X(_0609_));
 sky130_fd_sc_hd__or2_4 _0760_ (.A(_0609_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit8.Q ),
    .X(_0610_));
 sky130_fd_sc_hd__mux4_1 _0761_ (.A0(net639),
    .A1(net629),
    .A2(net624),
    .A3(net406),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit7.Q ),
    .X(_0611_));
 sky130_fd_sc_hd__o21a_1 _0762_ (.A1(_0552_),
    .A2(_0611_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit9.Q ),
    .X(_0612_));
 sky130_fd_sc_hd__mux4_1 _0763_ (.A0(net814),
    .A1(net93),
    .A2(net121),
    .A3(net133),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit7.Q ),
    .X(_0613_));
 sky130_fd_sc_hd__mux4_1 _0764_ (.A0(net59),
    .A1(net65),
    .A2(net77),
    .A3(net10),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit7.Q ),
    .X(_0614_));
 sky130_fd_sc_hd__mux2_1 _0765_ (.A0(_0613_),
    .A1(_0614_),
    .S(_0552_),
    .X(_0615_));
 sky130_fd_sc_hd__a22o_4 _0766_ (.A1(_0612_),
    .A2(_0610_),
    .B1(_0615_),
    .B2(_0553_),
    .X(\Inst_LUT4AB_switch_matrix.E2BEG3 ));
 sky130_fd_sc_hd__mux4_2 _0767_ (.A0(net16),
    .A1(net99),
    .A2(net127),
    .A3(\Inst_LUT4AB_switch_matrix.E2BEG3 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit28.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit29.Q ),
    .X(_0616_));
 sky130_fd_sc_hd__mux4_2 _0768_ (.A0(net72),
    .A1(net17),
    .A2(net100),
    .A3(net128),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit28.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit29.Q ),
    .X(_0617_));
 sky130_fd_sc_hd__o21ba_1 _0769_ (.A1(_0554_),
    .A2(_0617_),
    .B1_N(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit6.Q ),
    .X(_0618_));
 sky130_fd_sc_hd__o21a_1 _0770_ (.A1(_0616_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit5.Q ),
    .B1(_0618_),
    .X(_0619_));
 sky130_fd_sc_hd__nor2_1 _0771_ (.A(_0608_),
    .B(_0619_),
    .Y(_0620_));
 sky130_fd_sc_hd__mux4_1 _0772_ (.A0(net659),
    .A1(net655),
    .A2(net650),
    .A3(net645),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit7.Q ),
    .X(_0621_));
 sky130_fd_sc_hd__mux4_1 _0773_ (.A0(net640),
    .A1(net630),
    .A2(net625),
    .A3(net622),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit7.Q ),
    .X(_0622_));
 sky130_fd_sc_hd__mux2_4 _0774_ (.A0(_0621_),
    .A1(_0622_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit8.Q ),
    .X(_0623_));
 sky130_fd_sc_hd__mux4_1 _0775_ (.A0(net65),
    .A1(net816),
    .A2(net77),
    .A3(net10),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit7.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit6.Q ),
    .X(_0624_));
 sky130_fd_sc_hd__and2b_1 _0776_ (.A_N(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit8.Q ),
    .B(_0624_),
    .X(_0625_));
 sky130_fd_sc_hd__mux4_1 _0777_ (.A0(net814),
    .A1(net93),
    .A2(net121),
    .A3(net133),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit7.Q ),
    .X(_0626_));
 sky130_fd_sc_hd__a21o_1 _0778_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit8.Q ),
    .A2(_0626_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit9.Q ),
    .X(_0627_));
 sky130_fd_sc_hd__o22a_4 _0779_ (.A1(_0623_),
    .A2(_0548_),
    .B1(_0625_),
    .B2(_0627_),
    .X(\Inst_LUT4AB_switch_matrix.JN2BEG3 ));
 sky130_fd_sc_hd__mux4_2 _0780_ (.A0(net75),
    .A1(net103),
    .A2(net131),
    .A3(\Inst_LUT4AB_switch_matrix.JN2BEG3 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit26.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit27.Q ),
    .X(_0628_));
 sky130_fd_sc_hd__mux4_1 _0781_ (.A0(net76),
    .A1(net21),
    .A2(net104),
    .A3(net132),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit26.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit27.Q ),
    .X(_0629_));
 sky130_fd_sc_hd__o21ba_1 _0782_ (.A1(_0549_),
    .A2(_0629_),
    .B1_N(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit4.Q ),
    .X(_0630_));
 sky130_fd_sc_hd__o21a_1 _0783_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit3.Q ),
    .A2(_0628_),
    .B1(_0630_),
    .X(_0631_));
 sky130_fd_sc_hd__mux4_1 _0784_ (.A0(net659),
    .A1(net634),
    .A2(net649),
    .A3(net645),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit31.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit30.Q ),
    .X(_0632_));
 sky130_fd_sc_hd__mux4_2 _0785_ (.A0(net639),
    .A1(net629),
    .A2(net624),
    .A3(net403),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit30.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit31.Q ),
    .X(_0633_));
 sky130_fd_sc_hd__mux2_4 _0786_ (.A0(_0632_),
    .A1(_0633_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit0.Q ),
    .X(_0634_));
 sky130_fd_sc_hd__mux4_1 _0787_ (.A0(net814),
    .A1(net91),
    .A2(net119),
    .A3(net133),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit30.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit31.Q ),
    .X(_0635_));
 sky130_fd_sc_hd__mux4_1 _0788_ (.A0(net63),
    .A1(net2),
    .A2(net79),
    .A3(net8),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit31.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit30.Q ),
    .X(_0636_));
 sky130_fd_sc_hd__nand2b_1 _0789_ (.A_N(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit0.Q ),
    .B(_0636_),
    .Y(_0637_));
 sky130_fd_sc_hd__a21oi_1 _0790_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit0.Q ),
    .A2(_0635_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit1.Q ),
    .Y(_0638_));
 sky130_fd_sc_hd__o2bb2a_4 _0791_ (.A1_N(_0637_),
    .A2_N(_0638_),
    .B1(_0550_),
    .B2(_0634_),
    .X(\Inst_LUT4AB_switch_matrix.JN2BEG1 ));
 sky130_fd_sc_hd__mux4_2 _0792_ (.A0(net84),
    .A1(net135),
    .A2(net108),
    .A3(\Inst_LUT4AB_switch_matrix.JN2BEG1 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit27.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit26.Q ),
    .X(_0639_));
 sky130_fd_sc_hd__mux4_2 _0793_ (.A0(net67),
    .A1(net112),
    .A2(net12),
    .A3(net123),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit27.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit26.Q ),
    .X(_0640_));
 sky130_fd_sc_hd__mux2_4 _0794_ (.A0(_0639_),
    .A1(_0640_),
    .S(_0549_),
    .X(_0641_));
 sky130_fd_sc_hd__a211o_1 _0795_ (.A1(_0641_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit4.Q ),
    .B1(_0631_),
    .C1(\Inst_LA_LUT4c_frame_config_dffesr.c_I0mux ),
    .X(_0642_));
 sky130_fd_sc_hd__o21ai_4 _0796_ (.A1(_0551_),
    .A2(net1),
    .B1(_0642_),
    .Y(_0643_));
 sky130_fd_sc_hd__mux2_4 _0797_ (.A0(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ),
    .A1(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ),
    .S(_0643_),
    .X(_0644_));
 sky130_fd_sc_hd__mux4_2 _0798_ (.A0(net659),
    .A1(net654),
    .A2(net649),
    .A3(net644),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit7.Q ),
    .X(_0645_));
 sky130_fd_sc_hd__or2_4 _0799_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit8.Q ),
    .B(_0645_),
    .X(_0646_));
 sky130_fd_sc_hd__mux4_2 _0800_ (.A0(net640),
    .A1(net630),
    .A2(net624),
    .A3(net397),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit7.Q ),
    .X(_0647_));
 sky130_fd_sc_hd__o21a_1 _0801_ (.A1(_0557_),
    .A2(_0647_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit9.Q ),
    .X(_0648_));
 sky130_fd_sc_hd__mux4_1 _0802_ (.A0(net65),
    .A1(net816),
    .A2(net10),
    .A3(net814),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit7.Q ),
    .X(_0649_));
 sky130_fd_sc_hd__mux4_1 _0803_ (.A0(net93),
    .A1(net121),
    .A2(net105),
    .A3(net137),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit7.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit6.Q ),
    .X(_0650_));
 sky130_fd_sc_hd__mux2_1 _0804_ (.A0(_0649_),
    .A1(_0650_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit8.Q ),
    .X(_0651_));
 sky130_fd_sc_hd__a22o_1 _0805_ (.A1(_0648_),
    .A2(_0646_),
    .B1(_0651_),
    .B2(_0558_),
    .X(\Inst_LUT4AB_switch_matrix.JS2BEG3 ));
 sky130_fd_sc_hd__mux4_2 _0806_ (.A0(net73),
    .A1(net18),
    .A2(net129),
    .A3(\Inst_LUT4AB_switch_matrix.JS2BEG3 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit30.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit31.Q ),
    .X(_0652_));
 sky130_fd_sc_hd__mux4_2 _0807_ (.A0(net74),
    .A1(net19),
    .A2(net102),
    .A3(net130),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit30.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit31.Q ),
    .X(_0653_));
 sky130_fd_sc_hd__mux4_1 _0808_ (.A0(net426),
    .A1(net634),
    .A2(net649),
    .A3(net644),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit31.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit30.Q ),
    .X(_0654_));
 sky130_fd_sc_hd__or2_1 _0809_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit0.Q ),
    .B(_0654_),
    .X(_0655_));
 sky130_fd_sc_hd__mux4_1 _0810_ (.A0(net639),
    .A1(net629),
    .A2(net624),
    .A3(net622),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit30.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit31.Q ),
    .X(_0656_));
 sky130_fd_sc_hd__o21a_1 _0811_ (.A1(_0559_),
    .A2(_0656_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit1.Q ),
    .X(_0657_));
 sky130_fd_sc_hd__mux4_1 _0812_ (.A0(net107),
    .A1(net111),
    .A2(net119),
    .A3(net133),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit30.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit31.Q ),
    .X(_0658_));
 sky130_fd_sc_hd__mux4_1 _0813_ (.A0(net83),
    .A1(net26),
    .A2(net2),
    .A3(net814),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit31.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit30.Q ),
    .X(_0659_));
 sky130_fd_sc_hd__mux2_1 _0814_ (.A0(_0658_),
    .A1(_0659_),
    .S(_0559_),
    .X(_0660_));
 sky130_fd_sc_hd__a22o_1 _0815_ (.A1(_0657_),
    .A2(_0655_),
    .B1(_0660_),
    .B2(_0560_),
    .X(\Inst_LUT4AB_switch_matrix.JS2BEG1 ));
 sky130_fd_sc_hd__mux4_2 _0816_ (.A0(net78),
    .A1(net813),
    .A2(net134),
    .A3(\Inst_LUT4AB_switch_matrix.JS2BEG1 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit30.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit31.Q ),
    .X(_0661_));
 sky130_fd_sc_hd__mux4_2 _0817_ (.A0(net65),
    .A1(net93),
    .A2(net24),
    .A3(net121),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit31.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit30.Q ),
    .X(_0662_));
 sky130_fd_sc_hd__mux4_2 _0818_ (.A0(_0652_),
    .A1(_0653_),
    .A2(_0662_),
    .A3(_0661_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit7.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit8.Q ),
    .X(_0663_));
 sky130_fd_sc_hd__mux2_4 _0819_ (.A0(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ),
    .A1(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ),
    .S(_0643_),
    .X(_0664_));
 sky130_fd_sc_hd__mux2_1 _0820_ (.A0(_0664_),
    .A1(_0644_),
    .S(_0620_),
    .X(_0665_));
 sky130_fd_sc_hd__mux4_2 _0821_ (.A0(net426),
    .A1(net430),
    .A2(net649),
    .A3(net644),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit7.Q ),
    .X(_0666_));
 sky130_fd_sc_hd__mux4_1 _0822_ (.A0(net639),
    .A1(net629),
    .A2(net624),
    .A3(net623),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit7.Q ),
    .X(_0667_));
 sky130_fd_sc_hd__mux2_4 _0823_ (.A0(_0666_),
    .A1(_0667_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit8.Q ),
    .X(_0668_));
 sky130_fd_sc_hd__mux4_1 _0824_ (.A0(net59),
    .A1(net10),
    .A2(net65),
    .A3(net814),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit7.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit6.Q ),
    .X(_0669_));
 sky130_fd_sc_hd__and2b_1 _0825_ (.A_N(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit8.Q ),
    .B(_0669_),
    .X(_0670_));
 sky130_fd_sc_hd__mux4_1 _0826_ (.A0(net93),
    .A1(net121),
    .A2(net105),
    .A3(net137),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit7.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit6.Q ),
    .X(_0671_));
 sky130_fd_sc_hd__a21o_1 _0827_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit8.Q ),
    .A2(_0671_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit9.Q ),
    .X(_0672_));
 sky130_fd_sc_hd__o22a_4 _0828_ (.A1(_0668_),
    .A2(_0561_),
    .B1(_0670_),
    .B2(_0672_),
    .X(\Inst_LUT4AB_switch_matrix.JW2BEG3 ));
 sky130_fd_sc_hd__mux4_2 _0829_ (.A0(net69),
    .A1(net14),
    .A2(net97),
    .A3(\Inst_LUT4AB_switch_matrix.JW2BEG3 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit0.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit1.Q ),
    .X(_0673_));
 sky130_fd_sc_hd__mux4_1 _0830_ (.A0(net70),
    .A1(net15),
    .A2(net98),
    .A3(net126),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit0.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit1.Q ),
    .X(_0674_));
 sky130_fd_sc_hd__mux4_2 _0831_ (.A0(net426),
    .A1(net634),
    .A2(net649),
    .A3(net644),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit31.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit30.Q ),
    .X(_0675_));
 sky130_fd_sc_hd__mux4_1 _0832_ (.A0(net639),
    .A1(net629),
    .A2(net624),
    .A3(net416),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit30.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit31.Q ),
    .X(_0676_));
 sky130_fd_sc_hd__mux2_4 _0833_ (.A0(_0675_),
    .A1(_0676_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit0.Q ),
    .X(_0677_));
 sky130_fd_sc_hd__mux4_1 _0834_ (.A0(net57),
    .A1(net8),
    .A2(net63),
    .A3(net814),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit31.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit30.Q ),
    .X(_0678_));
 sky130_fd_sc_hd__and2b_1 _0835_ (.A_N(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit0.Q ),
    .B(_0678_),
    .X(_0679_));
 sky130_fd_sc_hd__mux4_1 _0836_ (.A0(net91),
    .A1(net119),
    .A2(net107),
    .A3(net133),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit31.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit30.Q ),
    .X(_0680_));
 sky130_fd_sc_hd__a21o_1 _0837_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit0.Q ),
    .A2(_0680_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit1.Q ),
    .X(_0681_));
 sky130_fd_sc_hd__o22a_4 _0838_ (.A1(_0677_),
    .A2(_0562_),
    .B1(_0679_),
    .B2(_0681_),
    .X(\Inst_LUT4AB_switch_matrix.JW2BEG1 ));
 sky130_fd_sc_hd__mux4_2 _0839_ (.A0(net77),
    .A1(net814),
    .A2(net105),
    .A3(\Inst_LUT4AB_switch_matrix.JW2BEG1 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit0.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit1.Q ),
    .X(_0682_));
 sky130_fd_sc_hd__mux4_2 _0840_ (.A0(net61),
    .A1(net89),
    .A2(net6),
    .A3(net138),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit1.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit0.Q ),
    .X(_0683_));
 sky130_fd_sc_hd__mux4_2 _0841_ (.A0(_0673_),
    .A1(_0674_),
    .A2(_0683_),
    .A3(_0682_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit9.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit10.Q ),
    .X(_0684_));
 sky130_fd_sc_hd__mux2_1 _0842_ (.A0(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ),
    .A1(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ),
    .S(_0643_),
    .X(_0685_));
 sky130_fd_sc_hd__mux2_1 _0843_ (.A0(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ),
    .A1(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ),
    .S(_0643_),
    .X(_0686_));
 sky130_fd_sc_hd__mux2_1 _0844_ (.A0(_0686_),
    .A1(_0685_),
    .S(_0620_),
    .X(_0687_));
 sky130_fd_sc_hd__mux2_1 _0845_ (.A0(_0687_),
    .A1(_0665_),
    .S(_0663_),
    .X(_0688_));
 sky130_fd_sc_hd__mux2_1 _0846_ (.A0(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ),
    .A1(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ),
    .S(_0643_),
    .X(_0689_));
 sky130_fd_sc_hd__mux2_1 _0847_ (.A0(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ),
    .A1(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ),
    .S(_0643_),
    .X(_0690_));
 sky130_fd_sc_hd__mux2_1 _0848_ (.A0(_0690_),
    .A1(_0689_),
    .S(_0620_),
    .X(_0691_));
 sky130_fd_sc_hd__mux2_1 _0849_ (.A0(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ),
    .A1(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ),
    .S(_0643_),
    .X(_0692_));
 sky130_fd_sc_hd__mux2_1 _0850_ (.A0(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ),
    .A1(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ),
    .S(_0643_),
    .X(_0693_));
 sky130_fd_sc_hd__mux2_1 _0851_ (.A0(_0692_),
    .A1(_0693_),
    .S(_0620_),
    .X(_0694_));
 sky130_fd_sc_hd__mux2_1 _0852_ (.A0(_0694_),
    .A1(_0691_),
    .S(_0663_),
    .X(_0695_));
 sky130_fd_sc_hd__mux2_4 _0853_ (.A0(_0695_),
    .A1(_0688_),
    .S(_0684_),
    .X(_0696_));
 sky130_fd_sc_hd__mux2_4 _0854_ (.A0(_0696_),
    .A1(\Inst_LA_LUT4c_frame_config_dffesr.LUT_flop ),
    .S(\Inst_LA_LUT4c_frame_config_dffesr.c_out_mux ),
    .X(A));
 sky130_fd_sc_hd__mux2_4 _0855_ (.A0(_0640_),
    .A1(_0639_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit13.Q ),
    .X(_0008_));
 sky130_fd_sc_hd__mux2_1 _0856_ (.A0(_0628_),
    .A1(_0629_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit13.Q ),
    .X(_0009_));
 sky130_fd_sc_hd__mux2_2 _0857_ (.A0(_0009_),
    .A1(_0008_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit14.Q ),
    .X(_0010_));
 sky130_fd_sc_hd__or2_4 _0858_ (.A(_0663_),
    .B(net1),
    .X(_0011_));
 sky130_fd_sc_hd__a211o_1 _0859_ (.A1(net1),
    .A2(_0663_),
    .B1(_0608_),
    .C1(_0619_),
    .X(_0012_));
 sky130_fd_sc_hd__and2b_1 _0860_ (.A_N(\Inst_LB_LUT4c_frame_config_dffesr.c_I0mux ),
    .B(_0010_),
    .X(_0013_));
 sky130_fd_sc_hd__a31o_1 _0861_ (.A1(_0012_),
    .A2(_0011_),
    .A3(\Inst_LB_LUT4c_frame_config_dffesr.c_I0mux ),
    .B1(_0013_),
    .X(_0014_));
 sky130_fd_sc_hd__mux4_2 _0862_ (.A0(_0673_),
    .A1(_0674_),
    .A2(_0683_),
    .A3(_0682_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit19.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit20.Q ),
    .X(_0015_));
 sky130_fd_sc_hd__mux4_2 _0863_ (.A0(_0652_),
    .A1(_0653_),
    .A2(_0662_),
    .A3(_0661_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit17.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit18.Q ),
    .X(_0016_));
 sky130_fd_sc_hd__mux4_2 _0864_ (.A0(_0616_),
    .A1(_0617_),
    .A2(_0606_),
    .A3(_0605_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit15.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit16.Q ),
    .X(_0017_));
 sky130_fd_sc_hd__nand2b_1 _0865_ (.A_N(_0016_),
    .B(_0017_),
    .Y(_0018_));
 sky130_fd_sc_hd__nand2b_1 _0866_ (.A_N(_0017_),
    .B(_0016_),
    .Y(_0019_));
 sky130_fd_sc_hd__o22a_1 _0867_ (.A1(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ),
    .A2(_0018_),
    .B1(_0019_),
    .B2(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ),
    .X(_0020_));
 sky130_fd_sc_hd__and2_4 _0868_ (.A(_0016_),
    .B(_0017_),
    .X(_0021_));
 sky130_fd_sc_hd__nand2_1 _0869_ (.A(_0016_),
    .B(_0017_),
    .Y(_0022_));
 sky130_fd_sc_hd__or2_2 _0870_ (.A(_0016_),
    .B(_0017_),
    .X(_0023_));
 sky130_fd_sc_hd__o221a_1 _0871_ (.A1(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ),
    .A2(_0022_),
    .B1(_0023_),
    .B2(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ),
    .C1(_0020_),
    .X(_0024_));
 sky130_fd_sc_hd__o22a_1 _0872_ (.A1(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ),
    .A2(_0018_),
    .B1(_0019_),
    .B2(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ),
    .X(_0025_));
 sky130_fd_sc_hd__o221a_1 _0873_ (.A1(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ),
    .A2(_0022_),
    .B1(_0023_),
    .B2(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ),
    .C1(_0025_),
    .X(_0026_));
 sky130_fd_sc_hd__mux2_4 _0874_ (.A0(_0024_),
    .A1(_0026_),
    .S(_0015_),
    .X(_0027_));
 sky130_fd_sc_hd__or2_1 _0875_ (.A(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ),
    .B(_0019_),
    .X(_0028_));
 sky130_fd_sc_hd__o221a_1 _0876_ (.A1(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ),
    .A2(_0022_),
    .B1(_0023_),
    .B2(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ),
    .C1(_0028_),
    .X(_0029_));
 sky130_fd_sc_hd__o211a_1 _0877_ (.A1(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ),
    .A2(_0018_),
    .B1(_0029_),
    .C1(_0015_),
    .X(_0030_));
 sky130_fd_sc_hd__o21ba_1 _0878_ (.A1(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ),
    .A2(_0019_),
    .B1_N(_0015_),
    .X(_0031_));
 sky130_fd_sc_hd__o22a_1 _0879_ (.A1(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ),
    .A2(_0018_),
    .B1(_0022_),
    .B2(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ),
    .X(_0032_));
 sky130_fd_sc_hd__o211a_1 _0880_ (.A1(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ),
    .A2(_0023_),
    .B1(_0031_),
    .C1(_0032_),
    .X(_0033_));
 sky130_fd_sc_hd__or3b_1 _0881_ (.A(_0030_),
    .B(_0033_),
    .C_N(_0014_),
    .X(_0034_));
 sky130_fd_sc_hd__o21a_1 _0882_ (.A1(_0014_),
    .A2(_0027_),
    .B1(_0034_),
    .X(_0035_));
 sky130_fd_sc_hd__mux2_4 _0883_ (.A0(_0035_),
    .A1(\Inst_LB_LUT4c_frame_config_dffesr.LUT_flop ),
    .S(\Inst_LB_LUT4c_frame_config_dffesr.c_out_mux ),
    .X(B));
 sky130_fd_sc_hd__mux4_1 _0884_ (.A0(net661),
    .A1(net658),
    .A2(net638),
    .A3(net648),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit3.Q ),
    .X(_0036_));
 sky130_fd_sc_hd__mux4_1 _0885_ (.A0(net642),
    .A1(net633),
    .A2(H),
    .A3(net405),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit3.Q ),
    .X(_0037_));
 sky130_fd_sc_hd__mux2_4 _0886_ (.A0(_0036_),
    .A1(_0037_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit4.Q ),
    .X(_0038_));
 sky130_fd_sc_hd__mux4_1 _0887_ (.A0(net58),
    .A1(net80),
    .A2(net64),
    .A3(net9),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit3.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit2.Q ),
    .X(_0039_));
 sky130_fd_sc_hd__and2b_1 _0888_ (.A_N(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit4.Q ),
    .B(_0039_),
    .X(_0040_));
 sky130_fd_sc_hd__mux4_1 _0889_ (.A0(net813),
    .A1(net92),
    .A2(net120),
    .A3(net134),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit3.Q ),
    .X(_0041_));
 sky130_fd_sc_hd__a21o_1 _0890_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit4.Q ),
    .A2(_0041_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit5.Q ),
    .X(_0042_));
 sky130_fd_sc_hd__o22a_4 _0891_ (.A1(_0565_),
    .A2(_0038_),
    .B1(_0040_),
    .B2(_0042_),
    .X(\Inst_LUT4AB_switch_matrix.E2BEG2 ));
 sky130_fd_sc_hd__mux4_2 _0892_ (.A0(net79),
    .A1(net8),
    .A2(net124),
    .A3(\Inst_LUT4AB_switch_matrix.E2BEG2 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit4.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit5.Q ),
    .X(_0043_));
 sky130_fd_sc_hd__mux4_2 _0893_ (.A0(net63),
    .A1(net8),
    .A2(net91),
    .A3(net137),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit4.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit5.Q ),
    .X(_0044_));
 sky130_fd_sc_hd__mux4_2 _0894_ (.A0(net661),
    .A1(net656),
    .A2(C),
    .A3(net637),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit10.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit11.Q ),
    .X(_0045_));
 sky130_fd_sc_hd__and2b_1 _0895_ (.A_N(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit12.Q ),
    .B(_0045_),
    .X(_0046_));
 sky130_fd_sc_hd__mux4_1 _0896_ (.A0(net641),
    .A1(net632),
    .A2(H),
    .A3(\Inst_LUT4AB_switch_matrix.M_EF ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit10.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit11.Q ),
    .X(_0047_));
 sky130_fd_sc_hd__a21bo_1 _0897_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit12.Q ),
    .A2(_0047_),
    .B1_N(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit13.Q ),
    .X(_0048_));
 sky130_fd_sc_hd__mux4_1 _0898_ (.A0(net86),
    .A1(net94),
    .A2(net88),
    .A3(net114),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit11.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit10.Q ),
    .X(_0049_));
 sky130_fd_sc_hd__mux4_1 _0899_ (.A0(net58),
    .A1(net66),
    .A2(net3),
    .A3(net11),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit10.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit11.Q ),
    .X(_0050_));
 sky130_fd_sc_hd__mux2_1 _0900_ (.A0(_0050_),
    .A1(_0049_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit12.Q ),
    .X(_0051_));
 sky130_fd_sc_hd__o22a_4 _0901_ (.A1(_0048_),
    .A2(_0046_),
    .B1(_0051_),
    .B2(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit13.Q ),
    .X(\Inst_LUT4AB_switch_matrix.E2BEG4 ));
 sky130_fd_sc_hd__mux4_2 _0902_ (.A0(net71),
    .A1(net127),
    .A2(net16),
    .A3(\Inst_LUT4AB_switch_matrix.E2BEG4 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit5.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit4.Q ),
    .X(_0052_));
 sky130_fd_sc_hd__mux4_2 _0903_ (.A0(net72),
    .A1(net17),
    .A2(net100),
    .A3(net128),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit4.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit5.Q ),
    .X(_0053_));
 sky130_fd_sc_hd__mux4_2 _0904_ (.A0(_0052_),
    .A1(_0053_),
    .A2(_0044_),
    .A3(_0043_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit3.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit4.Q ),
    .X(_0054_));
 sky130_fd_sc_hd__mux4_2 _0905_ (.A0(net659),
    .A1(net655),
    .A2(net635),
    .A3(net648),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit3.Q ),
    .X(_0055_));
 sky130_fd_sc_hd__and2b_1 _0906_ (.A_N(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit4.Q ),
    .B(_0055_),
    .X(_0056_));
 sky130_fd_sc_hd__mux4_1 _0907_ (.A0(net424),
    .A1(net630),
    .A2(net626),
    .A3(net623),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit3.Q ),
    .X(_0057_));
 sky130_fd_sc_hd__a21bo_1 _0908_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit4.Q ),
    .A2(_0057_),
    .B1_N(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit5.Q ),
    .X(_0058_));
 sky130_fd_sc_hd__mux4_1 _0909_ (.A0(net92),
    .A1(net120),
    .A2(net108),
    .A3(net134),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit3.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit2.Q ),
    .X(_0059_));
 sky130_fd_sc_hd__mux4_1 _0910_ (.A0(net84),
    .A1(net3),
    .A2(net9),
    .A3(net813),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit3.Q ),
    .X(_0060_));
 sky130_fd_sc_hd__mux2_1 _0911_ (.A0(_0060_),
    .A1(_0059_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit4.Q ),
    .X(_0061_));
 sky130_fd_sc_hd__o22a_4 _0912_ (.A1(_0058_),
    .A2(_0056_),
    .B1(_0061_),
    .B2(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit5.Q ),
    .X(\Inst_LUT4AB_switch_matrix.JS2BEG2 ));
 sky130_fd_sc_hd__mux4_2 _0913_ (.A0(net82),
    .A1(net25),
    .A2(net106),
    .A3(\Inst_LUT4AB_switch_matrix.JS2BEG2 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit7.Q ),
    .X(_0062_));
 sky130_fd_sc_hd__mux4_2 _0914_ (.A0(net65),
    .A1(net10),
    .A2(net111),
    .A3(net121),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit7.Q ),
    .X(_0063_));
 sky130_fd_sc_hd__mux4_1 _0915_ (.A0(net661),
    .A1(net658),
    .A2(C),
    .A3(net637),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit10.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit11.Q ),
    .X(_0064_));
 sky130_fd_sc_hd__mux4_2 _0916_ (.A0(net641),
    .A1(net631),
    .A2(net410),
    .A3(net427),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit10.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit11.Q ),
    .X(_0065_));
 sky130_fd_sc_hd__mux2_4 _0917_ (.A0(_0064_),
    .A1(_0065_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit12.Q ),
    .X(_0066_));
 sky130_fd_sc_hd__mux4_1 _0918_ (.A0(net58),
    .A1(net66),
    .A2(net3),
    .A3(net11),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit10.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit11.Q ),
    .X(_0067_));
 sky130_fd_sc_hd__and2b_1 _0919_ (.A_N(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit12.Q ),
    .B(_0067_),
    .X(_0068_));
 sky130_fd_sc_hd__mux4_1 _0920_ (.A0(net86),
    .A1(net94),
    .A2(net114),
    .A3(net116),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit10.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit11.Q ),
    .X(_0069_));
 sky130_fd_sc_hd__a21o_1 _0921_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit12.Q ),
    .A2(_0069_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit13.Q ),
    .X(_0070_));
 sky130_fd_sc_hd__o22a_4 _0922_ (.A1(_0066_),
    .A2(_0566_),
    .B1(_0068_),
    .B2(_0070_),
    .X(\Inst_LUT4AB_switch_matrix.JS2BEG4 ));
 sky130_fd_sc_hd__mux4_2 _0923_ (.A0(net73),
    .A1(net18),
    .A2(net101),
    .A3(\Inst_LUT4AB_switch_matrix.JS2BEG4 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit7.Q ),
    .X(_0071_));
 sky130_fd_sc_hd__mux4_1 _0924_ (.A0(net74),
    .A1(net19),
    .A2(net102),
    .A3(net130),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit7.Q ),
    .X(_0072_));
 sky130_fd_sc_hd__mux4_2 _0925_ (.A0(_0071_),
    .A1(_0072_),
    .A2(_0063_),
    .A3(_0062_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit5.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit6.Q ),
    .X(_0073_));
 sky130_fd_sc_hd__or2_4 _0926_ (.A(_0054_),
    .B(_0073_),
    .X(_0074_));
 sky130_fd_sc_hd__nand2_4 _0927_ (.A(_0073_),
    .B(_0054_),
    .Y(_0075_));
 sky130_fd_sc_hd__inv_2 _0928_ (.A(_0075_),
    .Y(_0076_));
 sky130_fd_sc_hd__mux4_2 _0929_ (.A0(_0052_),
    .A1(_0053_),
    .A2(_0044_),
    .A3(_0043_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit25.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit26.Q ),
    .X(_0077_));
 sky130_fd_sc_hd__mux4_2 _0930_ (.A0(_0071_),
    .A1(_0072_),
    .A2(_0063_),
    .A3(_0062_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit27.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit28.Q ),
    .X(_0078_));
 sky130_fd_sc_hd__nor2_2 _0931_ (.A(_0077_),
    .B(_0078_),
    .Y(_0079_));
 sky130_fd_sc_hd__inv_2 _0932_ (.A(_0079_),
    .Y(_0080_));
 sky130_fd_sc_hd__and2_1 _0933_ (.A(_0077_),
    .B(_0078_),
    .X(_0081_));
 sky130_fd_sc_hd__a31o_1 _0934_ (.A1(_0012_),
    .A2(_0011_),
    .A3(_0023_),
    .B1(_0021_),
    .X(_0082_));
 sky130_fd_sc_hd__a311o_1 _0935_ (.A1(_0011_),
    .A2(_0012_),
    .A3(_0023_),
    .B1(_0021_),
    .C1(_0081_),
    .X(_0083_));
 sky130_fd_sc_hd__a31o_1 _0936_ (.A1(_0083_),
    .A2(_0080_),
    .A3(_0074_),
    .B1(_0076_),
    .X(_0084_));
 sky130_fd_sc_hd__mux4_1 _0937_ (.A0(net646),
    .A1(net631),
    .A2(net627),
    .A3(net397),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit15.Q ),
    .X(_0085_));
 sky130_fd_sc_hd__mux4_1 _0938_ (.A0(net662),
    .A1(net656),
    .A2(net653),
    .A3(net636),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit15.Q ),
    .X(_0086_));
 sky130_fd_sc_hd__mux2_2 _0939_ (.A0(_0086_),
    .A1(_0085_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit16.Q ),
    .X(_0087_));
 sky130_fd_sc_hd__mux4_1 _0940_ (.A0(net59),
    .A1(net67),
    .A2(net816),
    .A3(net12),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit15.Q ),
    .X(_0088_));
 sky130_fd_sc_hd__and2b_1 _0941_ (.A_N(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit16.Q ),
    .B(_0088_),
    .X(_0089_));
 sky130_fd_sc_hd__mux4_1 _0942_ (.A0(net87),
    .A1(net113),
    .A2(net95),
    .A3(net666),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit15.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit14.Q ),
    .X(_0090_));
 sky130_fd_sc_hd__a21o_1 _0943_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit16.Q ),
    .A2(_0090_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit17.Q ),
    .X(_0091_));
 sky130_fd_sc_hd__o22a_4 _0944_ (.A1(_0087_),
    .A2(_0568_),
    .B1(_0089_),
    .B2(_0091_),
    .X(\Inst_LUT4AB_switch_matrix.JN2BEG5 ));
 sky130_fd_sc_hd__mux4_1 _0945_ (.A0(net75),
    .A1(net131),
    .A2(net20),
    .A3(\Inst_LUT4AB_switch_matrix.JN2BEG5 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit11.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit10.Q ),
    .X(_0092_));
 sky130_fd_sc_hd__mux4_2 _0946_ (.A0(net76),
    .A1(net21),
    .A2(net104),
    .A3(net132),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit10.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit11.Q ),
    .X(_0093_));
 sky130_fd_sc_hd__mux4_1 _0947_ (.A0(net80),
    .A1(net120),
    .A2(net9),
    .A3(\Inst_LUT4AB_switch_matrix.JN2BEG3 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit11.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit10.Q ),
    .X(_0094_));
 sky130_fd_sc_hd__mux4_2 _0948_ (.A0(net68),
    .A1(net96),
    .A2(net26),
    .A3(net124),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit11.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit10.Q ),
    .X(_0095_));
 sky130_fd_sc_hd__mux4_1 _0949_ (.A0(_0092_),
    .A1(_0093_),
    .A2(_0095_),
    .A3(_0094_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit11.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit12.Q ),
    .X(_0096_));
 sky130_fd_sc_hd__mux2_4 _0950_ (.A0(_0096_),
    .A1(_0084_),
    .S(\Inst_LE_LUT4c_frame_config_dffesr.c_I0mux ),
    .X(_0097_));
 sky130_fd_sc_hd__mux4_2 _0951_ (.A0(net78),
    .A1(net110),
    .A2(net121),
    .A3(\Inst_LUT4AB_switch_matrix.JS2BEG3 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit15.Q ),
    .X(_0098_));
 sky130_fd_sc_hd__mux4_2 _0952_ (.A0(net66),
    .A1(net11),
    .A2(net110),
    .A3(net122),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit15.Q ),
    .X(_0099_));
 sky130_fd_sc_hd__mux4_1 _0953_ (.A0(net660),
    .A1(net657),
    .A2(net652),
    .A3(net637),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit15.Q ),
    .X(_0100_));
 sky130_fd_sc_hd__mux4_2 _0954_ (.A0(net646),
    .A1(net631),
    .A2(net627),
    .A3(net622),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit15.Q ),
    .X(_0101_));
 sky130_fd_sc_hd__mux2_4 _0955_ (.A0(_0100_),
    .A1(_0101_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit16.Q ),
    .X(_0102_));
 sky130_fd_sc_hd__mux4_1 _0956_ (.A0(net59),
    .A1(net67),
    .A2(net816),
    .A3(net12),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit15.Q ),
    .X(_0103_));
 sky130_fd_sc_hd__and2b_1 _0957_ (.A_N(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit16.Q ),
    .B(_0103_),
    .X(_0104_));
 sky130_fd_sc_hd__mux4_1 _0958_ (.A0(net87),
    .A1(net113),
    .A2(net95),
    .A3(net666),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit15.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit14.Q ),
    .X(_0105_));
 sky130_fd_sc_hd__a21o_1 _0959_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit16.Q ),
    .A2(_0105_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit17.Q ),
    .X(_0106_));
 sky130_fd_sc_hd__o22a_1 _0960_ (.A1(_0102_),
    .A2(_0570_),
    .B1(_0104_),
    .B2(_0106_),
    .X(\Inst_LUT4AB_switch_matrix.JS2BEG5 ));
 sky130_fd_sc_hd__mux4_2 _0961_ (.A0(net73),
    .A1(net129),
    .A2(net101),
    .A3(net408),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit15.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit14.Q ),
    .X(_0107_));
 sky130_fd_sc_hd__mux4_1 _0962_ (.A0(net74),
    .A1(net19),
    .A2(net102),
    .A3(net130),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit15.Q ),
    .X(_0108_));
 sky130_fd_sc_hd__mux4_2 _0963_ (.A0(net431),
    .A1(_0108_),
    .A2(_0099_),
    .A3(_0098_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit15.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit16.Q ),
    .X(_0109_));
 sky130_fd_sc_hd__mux4_2 _0964_ (.A0(net83),
    .A1(net107),
    .A2(net8),
    .A3(\Inst_LUT4AB_switch_matrix.E2BEG3 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit13.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit12.Q ),
    .X(_0110_));
 sky130_fd_sc_hd__mux4_2 _0965_ (.A0(net64),
    .A1(net92),
    .A2(net9),
    .A3(net136),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit13.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit12.Q ),
    .X(_0111_));
 sky130_fd_sc_hd__mux4_1 _0966_ (.A0(net662),
    .A1(net656),
    .A2(net653),
    .A3(net636),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit15.Q ),
    .X(_0112_));
 sky130_fd_sc_hd__mux4_2 _0967_ (.A0(net646),
    .A1(net632),
    .A2(net410),
    .A3(net623),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit15.Q ),
    .X(_0113_));
 sky130_fd_sc_hd__mux2_4 _0968_ (.A0(_0112_),
    .A1(_0113_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit16.Q ),
    .X(_0114_));
 sky130_fd_sc_hd__mux4_1 _0969_ (.A0(net59),
    .A1(net67),
    .A2(net816),
    .A3(net12),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit15.Q ),
    .X(_0115_));
 sky130_fd_sc_hd__and2b_1 _0970_ (.A_N(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit16.Q ),
    .B(_0115_),
    .X(_0116_));
 sky130_fd_sc_hd__mux4_1 _0971_ (.A0(net85),
    .A1(net87),
    .A2(net95),
    .A3(net666),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit15.Q ),
    .X(_0117_));
 sky130_fd_sc_hd__a21o_1 _0972_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit16.Q ),
    .A2(_0117_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit17.Q ),
    .X(_0118_));
 sky130_fd_sc_hd__o22a_4 _0973_ (.A1(_0114_),
    .A2(_0569_),
    .B1(_0116_),
    .B2(_0118_),
    .X(\Inst_LUT4AB_switch_matrix.E2BEG5 ));
 sky130_fd_sc_hd__mux4_2 _0974_ (.A0(net71),
    .A1(net99),
    .A2(net16),
    .A3(\Inst_LUT4AB_switch_matrix.E2BEG5 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit13.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit12.Q ),
    .X(_0119_));
 sky130_fd_sc_hd__mux4_2 _0975_ (.A0(net72),
    .A1(net17),
    .A2(net100),
    .A3(net128),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit12.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit13.Q ),
    .X(_0120_));
 sky130_fd_sc_hd__mux4_2 _0976_ (.A0(_0119_),
    .A1(_0120_),
    .A2(_0111_),
    .A3(_0110_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit13.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit14.Q ),
    .X(_0121_));
 sky130_fd_sc_hd__nand2b_1 _0977_ (.A_N(_0109_),
    .B(_0121_),
    .Y(_0122_));
 sky130_fd_sc_hd__and2_1 _0978_ (.A(_0109_),
    .B(_0121_),
    .X(_0123_));
 sky130_fd_sc_hd__nand2_1 _0979_ (.A(_0109_),
    .B(_0121_),
    .Y(_0124_));
 sky130_fd_sc_hd__nand2b_1 _0980_ (.A_N(_0121_),
    .B(_0109_),
    .Y(_0125_));
 sky130_fd_sc_hd__or2_4 _0981_ (.A(_0109_),
    .B(_0121_),
    .X(_0126_));
 sky130_fd_sc_hd__o22a_1 _0982_ (.A1(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ),
    .A2(_0122_),
    .B1(_0125_),
    .B2(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ),
    .X(_0127_));
 sky130_fd_sc_hd__o221a_1 _0983_ (.A1(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ),
    .A2(_0124_),
    .B1(_0126_),
    .B2(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ),
    .C1(_0127_),
    .X(_0128_));
 sky130_fd_sc_hd__mux4_2 _0984_ (.A0(net27),
    .A1(net136),
    .A2(net105),
    .A3(\Inst_LUT4AB_switch_matrix.JW2BEG3 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit17.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit16.Q ),
    .X(_0129_));
 sky130_fd_sc_hd__mux4_2 _0985_ (.A0(net83),
    .A1(net7),
    .A2(net90),
    .A3(net118),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit16.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit17.Q ),
    .X(_0130_));
 sky130_fd_sc_hd__mux4_1 _0986_ (.A0(net660),
    .A1(net656),
    .A2(net652),
    .A3(net636),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit15.Q ),
    .X(_0131_));
 sky130_fd_sc_hd__mux4_2 _0987_ (.A0(net647),
    .A1(net632),
    .A2(net628),
    .A3(net398),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit15.Q ),
    .X(_0132_));
 sky130_fd_sc_hd__mux2_4 _0988_ (.A0(_0131_),
    .A1(_0132_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit16.Q ),
    .X(_0133_));
 sky130_fd_sc_hd__mux4_1 _0989_ (.A0(net85),
    .A1(net87),
    .A2(net95),
    .A3(net666),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit15.Q ),
    .X(_0134_));
 sky130_fd_sc_hd__mux4_1 _0990_ (.A0(net59),
    .A1(net67),
    .A2(net816),
    .A3(net12),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit15.Q ),
    .X(_0135_));
 sky130_fd_sc_hd__and2b_1 _0991_ (.A_N(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit16.Q ),
    .B(_0135_),
    .X(_0136_));
 sky130_fd_sc_hd__a21o_1 _0992_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit16.Q ),
    .A2(_0134_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit17.Q ),
    .X(_0137_));
 sky130_fd_sc_hd__o22a_4 _0993_ (.A1(_0571_),
    .A2(_0133_),
    .B1(_0136_),
    .B2(_0137_),
    .X(\Inst_LUT4AB_switch_matrix.JW2BEG5 ));
 sky130_fd_sc_hd__mux4_2 _0994_ (.A0(net14),
    .A1(net97),
    .A2(net125),
    .A3(\Inst_LUT4AB_switch_matrix.JW2BEG5 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit16.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit17.Q ),
    .X(_0138_));
 sky130_fd_sc_hd__mux4_2 _0995_ (.A0(net70),
    .A1(net15),
    .A2(net98),
    .A3(net126),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit16.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit17.Q ),
    .X(_0139_));
 sky130_fd_sc_hd__mux4_2 _0996_ (.A0(_0138_),
    .A1(_0139_),
    .A2(_0130_),
    .A3(_0129_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit17.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit18.Q ),
    .X(_0140_));
 sky130_fd_sc_hd__o22a_1 _0997_ (.A1(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ),
    .A2(_0122_),
    .B1(_0126_),
    .B2(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ),
    .X(_0141_));
 sky130_fd_sc_hd__or2_1 _0998_ (.A(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ),
    .B(_0125_),
    .X(_0142_));
 sky130_fd_sc_hd__o211a_1 _0999_ (.A1(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ),
    .A2(_0124_),
    .B1(_0141_),
    .C1(_0142_),
    .X(_0143_));
 sky130_fd_sc_hd__mux2_4 _1000_ (.A0(_0128_),
    .A1(_0143_),
    .S(_0097_),
    .X(_0144_));
 sky130_fd_sc_hd__o22a_1 _1001_ (.A1(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ),
    .A2(_0122_),
    .B1(_0125_),
    .B2(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ),
    .X(_0145_));
 sky130_fd_sc_hd__o221a_1 _1002_ (.A1(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ),
    .A2(_0124_),
    .B1(_0126_),
    .B2(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ),
    .C1(_0145_),
    .X(_0146_));
 sky130_fd_sc_hd__o22a_1 _1003_ (.A1(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ),
    .A2(_0122_),
    .B1(_0125_),
    .B2(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ),
    .X(_0147_));
 sky130_fd_sc_hd__o221a_1 _1004_ (.A1(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ),
    .A2(_0124_),
    .B1(_0126_),
    .B2(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ),
    .C1(_0147_),
    .X(_0148_));
 sky130_fd_sc_hd__mux2_1 _1005_ (.A0(_0146_),
    .A1(_0148_),
    .S(_0097_),
    .X(_0149_));
 sky130_fd_sc_hd__mux2_4 _1006_ (.A0(_0149_),
    .A1(_0144_),
    .S(_0140_),
    .X(_0150_));
 sky130_fd_sc_hd__mux2_4 _1007_ (.A0(_0150_),
    .A1(\Inst_LE_LUT4c_frame_config_dffesr.LUT_flop ),
    .S(\Inst_LE_LUT4c_frame_config_dffesr.c_out_mux ),
    .X(E));
 sky130_fd_sc_hd__mux4_1 _1008_ (.A0(net661),
    .A1(net658),
    .A2(net638),
    .A3(net647),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit3.Q ),
    .X(_0151_));
 sky130_fd_sc_hd__mux4_2 _1009_ (.A0(net643),
    .A1(net633),
    .A2(net628),
    .A3(net415),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit3.Q ),
    .X(_0152_));
 sky130_fd_sc_hd__mux2_4 _1010_ (.A0(_0151_),
    .A1(_0152_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit4.Q ),
    .X(_0153_));
 sky130_fd_sc_hd__mux4_1 _1011_ (.A0(net813),
    .A1(net92),
    .A2(net120),
    .A3(net136),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit3.Q ),
    .X(_0154_));
 sky130_fd_sc_hd__mux4_1 _1012_ (.A0(net64),
    .A1(net80),
    .A2(net3),
    .A3(net9),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit3.Q ),
    .X(_0155_));
 sky130_fd_sc_hd__and2b_1 _1013_ (.A_N(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit4.Q ),
    .B(_0155_),
    .X(_0156_));
 sky130_fd_sc_hd__a21o_1 _1014_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit4.Q ),
    .A2(_0154_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit5.Q ),
    .X(_0157_));
 sky130_fd_sc_hd__o22a_4 _1015_ (.A1(_0153_),
    .A2(_0564_),
    .B1(_0156_),
    .B2(_0157_),
    .X(\Inst_LUT4AB_switch_matrix.JN2BEG2 ));
 sky130_fd_sc_hd__mux4_1 _1016_ (.A0(net9),
    .A1(net137),
    .A2(net112),
    .A3(\Inst_LUT4AB_switch_matrix.JN2BEG2 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit3.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit2.Q ),
    .X(_0158_));
 sky130_fd_sc_hd__mux4_2 _1017_ (.A0(net84),
    .A1(net95),
    .A2(net12),
    .A3(net123),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit3.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit2.Q ),
    .X(_0159_));
 sky130_fd_sc_hd__mux4_1 _1018_ (.A0(net662),
    .A1(net656),
    .A2(net653),
    .A3(net636),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit10.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit11.Q ),
    .X(_0160_));
 sky130_fd_sc_hd__and2b_1 _1019_ (.A_N(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit12.Q ),
    .B(_0160_),
    .X(_0161_));
 sky130_fd_sc_hd__mux4_1 _1020_ (.A0(net642),
    .A1(net631),
    .A2(net627),
    .A3(net623),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit10.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit11.Q ),
    .X(_0162_));
 sky130_fd_sc_hd__a21bo_1 _1021_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit12.Q ),
    .A2(_0162_),
    .B1_N(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit13.Q ),
    .X(_0163_));
 sky130_fd_sc_hd__mux4_1 _1022_ (.A0(net58),
    .A1(net66),
    .A2(net3),
    .A3(net11),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit10.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit11.Q ),
    .X(_0164_));
 sky130_fd_sc_hd__mux4_1 _1023_ (.A0(net86),
    .A1(net94),
    .A2(net114),
    .A3(net665),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit10.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit11.Q ),
    .X(_0165_));
 sky130_fd_sc_hd__mux2_1 _1024_ (.A0(_0164_),
    .A1(_0165_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit12.Q ),
    .X(_0166_));
 sky130_fd_sc_hd__o22a_4 _1025_ (.A1(_0161_),
    .A2(_0163_),
    .B1(_0166_),
    .B2(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit13.Q ),
    .X(\Inst_LUT4AB_switch_matrix.JN2BEG4 ));
 sky130_fd_sc_hd__mux4_1 _1026_ (.A0(net20),
    .A1(net131),
    .A2(net103),
    .A3(\Inst_LUT4AB_switch_matrix.JN2BEG4 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit3.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit2.Q ),
    .X(_0167_));
 sky130_fd_sc_hd__mux4_1 _1027_ (.A0(net76),
    .A1(net21),
    .A2(net104),
    .A3(net132),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit3.Q ),
    .X(_0168_));
 sky130_fd_sc_hd__mux4_1 _1028_ (.A0(_0167_),
    .A1(_0168_),
    .A2(_0159_),
    .A3(_0158_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit23.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit24.Q ),
    .X(_0169_));
 sky130_fd_sc_hd__mux2_4 _1029_ (.A0(_0169_),
    .A1(_0082_),
    .S(\Inst_LC_LUT4c_frame_config_dffesr.c_I0mux ),
    .X(_0170_));
 sky130_fd_sc_hd__and2b_1 _1030_ (.A_N(_0077_),
    .B(_0078_),
    .X(_0171_));
 sky130_fd_sc_hd__and2b_1 _1031_ (.A_N(_0078_),
    .B(_0077_),
    .X(_0172_));
 sky130_fd_sc_hd__a22o_1 _1032_ (.A1(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ),
    .A2(_0171_),
    .B1(_0172_),
    .B2(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ),
    .X(_0173_));
 sky130_fd_sc_hd__a221o_1 _1033_ (.A1(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ),
    .A2(_0079_),
    .B1(_0081_),
    .B2(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ),
    .C1(_0173_),
    .X(_0174_));
 sky130_fd_sc_hd__mux4_1 _1034_ (.A0(net424),
    .A1(net399),
    .A2(net626),
    .A3(net432),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit3.Q ),
    .X(_0175_));
 sky130_fd_sc_hd__mux4_2 _1035_ (.A0(net426),
    .A1(net655),
    .A2(net635),
    .A3(net648),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit3.Q ),
    .X(_0176_));
 sky130_fd_sc_hd__and2b_1 _1036_ (.A_N(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit4.Q ),
    .B(_0176_),
    .X(_0177_));
 sky130_fd_sc_hd__a21bo_1 _1037_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit4.Q ),
    .A2(_0175_),
    .B1_N(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit5.Q ),
    .X(_0178_));
 sky130_fd_sc_hd__mux4_1 _1038_ (.A0(net108),
    .A1(net120),
    .A2(net112),
    .A3(net134),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit3.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit2.Q ),
    .X(_0179_));
 sky130_fd_sc_hd__mux4_1 _1039_ (.A0(net58),
    .A1(net64),
    .A2(net27),
    .A3(net813),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit3.Q ),
    .X(_0180_));
 sky130_fd_sc_hd__mux2_1 _1040_ (.A0(_0180_),
    .A1(_0179_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit4.Q ),
    .X(_0181_));
 sky130_fd_sc_hd__o22a_4 _1041_ (.A1(_0177_),
    .A2(_0178_),
    .B1(_0181_),
    .B2(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit5.Q ),
    .X(\Inst_LUT4AB_switch_matrix.JW2BEG2 ));
 sky130_fd_sc_hd__mux4_2 _1042_ (.A0(net77),
    .A1(net133),
    .A2(net109),
    .A3(\Inst_LUT4AB_switch_matrix.JW2BEG2 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit9.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit8.Q ),
    .X(_0182_));
 sky130_fd_sc_hd__mux4_2 _1043_ (.A0(net61),
    .A1(net89),
    .A2(net25),
    .A3(net117),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit9.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit8.Q ),
    .X(_0183_));
 sky130_fd_sc_hd__mux4_1 _1044_ (.A0(net660),
    .A1(net656),
    .A2(net652),
    .A3(net636),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit10.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit11.Q ),
    .X(_0184_));
 sky130_fd_sc_hd__mux4_2 _1045_ (.A0(net641),
    .A1(net631),
    .A2(net627),
    .A3(net402),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit10.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit11.Q ),
    .X(_0185_));
 sky130_fd_sc_hd__mux2_4 _1046_ (.A0(_0184_),
    .A1(_0185_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit12.Q ),
    .X(_0186_));
 sky130_fd_sc_hd__mux4_1 _1047_ (.A0(net58),
    .A1(net66),
    .A2(net3),
    .A3(net11),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit10.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit11.Q ),
    .X(_0187_));
 sky130_fd_sc_hd__and2b_1 _1048_ (.A_N(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit12.Q ),
    .B(_0187_),
    .X(_0188_));
 sky130_fd_sc_hd__mux4_1 _1049_ (.A0(net86),
    .A1(net94),
    .A2(net88),
    .A3(net114),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit11.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit10.Q ),
    .X(_0189_));
 sky130_fd_sc_hd__a21o_1 _1050_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit12.Q ),
    .A2(_0189_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit13.Q ),
    .X(_0190_));
 sky130_fd_sc_hd__o22a_4 _1051_ (.A1(_0567_),
    .A2(_0186_),
    .B1(_0188_),
    .B2(_0190_),
    .X(\Inst_LUT4AB_switch_matrix.JW2BEG4 ));
 sky130_fd_sc_hd__mux4_2 _1052_ (.A0(net69),
    .A1(net97),
    .A2(net125),
    .A3(\Inst_LUT4AB_switch_matrix.JW2BEG4 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit8.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit9.Q ),
    .X(_0191_));
 sky130_fd_sc_hd__mux4_2 _1053_ (.A0(net70),
    .A1(net15),
    .A2(net98),
    .A3(net126),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit8.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit9.Q ),
    .X(_0192_));
 sky130_fd_sc_hd__mux4_1 _1054_ (.A0(_0191_),
    .A1(_0192_),
    .A2(_0183_),
    .A3(_0182_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit29.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit30.Q ),
    .X(_0193_));
 sky130_fd_sc_hd__a22o_1 _1055_ (.A1(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ),
    .A2(_0081_),
    .B1(_0172_),
    .B2(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ),
    .X(_0194_));
 sky130_fd_sc_hd__a22o_1 _1056_ (.A1(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ),
    .A2(_0079_),
    .B1(_0171_),
    .B2(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ),
    .X(_0195_));
 sky130_fd_sc_hd__or2_1 _1057_ (.A(_0194_),
    .B(_0195_),
    .X(_0196_));
 sky130_fd_sc_hd__mux2_4 _1058_ (.A0(_0196_),
    .A1(_0174_),
    .S(_0170_),
    .X(_0197_));
 sky130_fd_sc_hd__a22o_1 _1059_ (.A1(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ),
    .A2(_0079_),
    .B1(_0171_),
    .B2(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ),
    .X(_0198_));
 sky130_fd_sc_hd__a221o_1 _1060_ (.A1(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ),
    .A2(_0081_),
    .B1(_0172_),
    .B2(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ),
    .C1(_0198_),
    .X(_0199_));
 sky130_fd_sc_hd__a22o_1 _1061_ (.A1(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ),
    .A2(_0171_),
    .B1(_0172_),
    .B2(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ),
    .X(_0200_));
 sky130_fd_sc_hd__a221o_1 _1062_ (.A1(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ),
    .A2(_0079_),
    .B1(_0081_),
    .B2(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ),
    .C1(_0200_),
    .X(_0201_));
 sky130_fd_sc_hd__mux2_1 _1063_ (.A0(_0201_),
    .A1(_0199_),
    .S(_0170_),
    .X(_0202_));
 sky130_fd_sc_hd__mux2_4 _1064_ (.A0(_0202_),
    .A1(_0197_),
    .S(_0193_),
    .X(_0203_));
 sky130_fd_sc_hd__mux2_4 _1065_ (.A0(_0203_),
    .A1(\Inst_LC_LUT4c_frame_config_dffesr.LUT_flop ),
    .S(\Inst_LC_LUT4c_frame_config_dffesr.c_out_mux ),
    .X(C));
 sky130_fd_sc_hd__a311o_1 _1066_ (.A1(_0083_),
    .A2(_0080_),
    .A3(_0074_),
    .B1(_0123_),
    .C1(_0076_),
    .X(_0204_));
 sky130_fd_sc_hd__a21bo_1 _1067_ (.A1(_0204_),
    .A2(_0126_),
    .B1_N(\Inst_LF_LUT4c_frame_config_dffesr.c_I0mux ),
    .X(_0205_));
 sky130_fd_sc_hd__mux4_1 _1068_ (.A0(_0092_),
    .A1(_0093_),
    .A2(_0095_),
    .A3(_0094_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit21.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit22.Q ),
    .X(_0206_));
 sky130_fd_sc_hd__o21a_1 _1069_ (.A1(\Inst_LF_LUT4c_frame_config_dffesr.c_I0mux ),
    .A2(_0206_),
    .B1(_0205_),
    .X(_0207_));
 sky130_fd_sc_hd__mux4_2 _1070_ (.A0(net431),
    .A1(_0108_),
    .A2(_0099_),
    .A3(_0098_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit25.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit26.Q ),
    .X(_0208_));
 sky130_fd_sc_hd__mux4_2 _1071_ (.A0(_0119_),
    .A1(_0120_),
    .A2(_0111_),
    .A3(_0110_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit23.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit24.Q ),
    .X(_0209_));
 sky130_fd_sc_hd__nor2_4 _1072_ (.A(_0209_),
    .B(_0208_),
    .Y(_0210_));
 sky130_fd_sc_hd__inv_2 _1073_ (.A(_0210_),
    .Y(_0211_));
 sky130_fd_sc_hd__and2_1 _1074_ (.A(_0208_),
    .B(_0209_),
    .X(_0212_));
 sky130_fd_sc_hd__and2b_1 _1075_ (.A_N(_0209_),
    .B(_0208_),
    .X(_0213_));
 sky130_fd_sc_hd__and2b_1 _1076_ (.A_N(_0208_),
    .B(_0209_),
    .X(_0214_));
 sky130_fd_sc_hd__a22o_1 _1077_ (.A1(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ),
    .A2(_0210_),
    .B1(_0213_),
    .B2(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ),
    .X(_0215_));
 sky130_fd_sc_hd__a22o_1 _1078_ (.A1(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ),
    .A2(_0212_),
    .B1(_0214_),
    .B2(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ),
    .X(_0216_));
 sky130_fd_sc_hd__or2_1 _1079_ (.A(_0215_),
    .B(_0216_),
    .X(_0217_));
 sky130_fd_sc_hd__mux4_2 _1080_ (.A0(_0138_),
    .A1(_0139_),
    .A2(_0130_),
    .A3(_0129_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit27.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit28.Q ),
    .X(_0218_));
 sky130_fd_sc_hd__a22o_1 _1081_ (.A1(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ),
    .A2(_0210_),
    .B1(_0212_),
    .B2(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ),
    .X(_0219_));
 sky130_fd_sc_hd__a22o_1 _1082_ (.A1(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ),
    .A2(_0213_),
    .B1(_0214_),
    .B2(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ),
    .X(_0220_));
 sky130_fd_sc_hd__or2_1 _1083_ (.A(_0219_),
    .B(_0220_),
    .X(_0221_));
 sky130_fd_sc_hd__mux2_4 _1084_ (.A0(_0221_),
    .A1(_0217_),
    .S(_0207_),
    .X(_0222_));
 sky130_fd_sc_hd__a22o_1 _1085_ (.A1(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ),
    .A2(_0213_),
    .B1(_0214_),
    .B2(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ),
    .X(_0223_));
 sky130_fd_sc_hd__a221o_1 _1086_ (.A1(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ),
    .A2(_0210_),
    .B1(_0212_),
    .B2(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ),
    .C1(_0223_),
    .X(_0224_));
 sky130_fd_sc_hd__a22o_1 _1087_ (.A1(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ),
    .A2(_0212_),
    .B1(_0213_),
    .B2(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ),
    .X(_0225_));
 sky130_fd_sc_hd__a221o_1 _1088_ (.A1(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ),
    .A2(_0210_),
    .B1(_0214_),
    .B2(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ),
    .C1(_0225_),
    .X(_0226_));
 sky130_fd_sc_hd__mux2_1 _1089_ (.A0(_0226_),
    .A1(_0224_),
    .S(_0207_),
    .X(_0227_));
 sky130_fd_sc_hd__mux2_4 _1090_ (.A0(_0222_),
    .A1(_0227_),
    .S(_0218_),
    .X(_0228_));
 sky130_fd_sc_hd__mux2_4 _1091_ (.A0(_0228_),
    .A1(\Inst_LF_LUT4c_frame_config_dffesr.LUT_flop ),
    .S(\Inst_LF_LUT4c_frame_config_dffesr.c_out_mux ),
    .X(F));
 sky130_fd_sc_hd__a31o_1 _1092_ (.A1(_0126_),
    .A2(_0204_),
    .A3(_0211_),
    .B1(_0212_),
    .X(_0229_));
 sky130_fd_sc_hd__mux4_2 _1093_ (.A0(net646),
    .A1(net627),
    .A2(net641),
    .A3(\Inst_LUT4AB_switch_matrix.M_AH ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit19.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit18.Q ),
    .X(_0230_));
 sky130_fd_sc_hd__mux4_1 _1094_ (.A0(net660),
    .A1(net656),
    .A2(net652),
    .A3(net636),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit18.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit19.Q ),
    .X(_0231_));
 sky130_fd_sc_hd__mux2_4 _1095_ (.A0(_0231_),
    .A1(_0230_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit20.Q ),
    .X(_0232_));
 sky130_fd_sc_hd__mux4_1 _1096_ (.A0(net88),
    .A1(net114),
    .A2(net96),
    .A3(net665),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit19.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit18.Q ),
    .X(_0233_));
 sky130_fd_sc_hd__mux4_1 _1097_ (.A0(net60),
    .A1(net68),
    .A2(net815),
    .A3(net13),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit18.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit19.Q ),
    .X(_0234_));
 sky130_fd_sc_hd__and2b_1 _1098_ (.A_N(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit20.Q ),
    .B(_0234_),
    .X(_0235_));
 sky130_fd_sc_hd__a211o_1 _1099_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit20.Q ),
    .A2(_0233_),
    .B1(_0235_),
    .C1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit21.Q ),
    .X(_0236_));
 sky130_fd_sc_hd__o21a_4 _1100_ (.A1(_0232_),
    .A2(_0563_),
    .B1(_0236_),
    .X(\Inst_LUT4AB_switch_matrix.JN2BEG6 ));
 sky130_fd_sc_hd__mux4_2 _1101_ (.A0(net75),
    .A1(net103),
    .A2(net20),
    .A3(\Inst_LUT4AB_switch_matrix.JN2BEG6 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit19.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit18.Q ),
    .X(_0237_));
 sky130_fd_sc_hd__mux4_2 _1102_ (.A0(net76),
    .A1(net21),
    .A2(net104),
    .A3(net132),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit18.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit19.Q ),
    .X(_0238_));
 sky130_fd_sc_hd__mux4_2 _1103_ (.A0(net80),
    .A1(net24),
    .A2(net108),
    .A3(\Inst_LUT4AB_switch_matrix.JN2BEG4 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit18.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit19.Q ),
    .X(_0239_));
 sky130_fd_sc_hd__mux4_2 _1104_ (.A0(net68),
    .A1(net13),
    .A2(net96),
    .A3(net135),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit18.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit19.Q ),
    .X(_0240_));
 sky130_fd_sc_hd__mux4_1 _1105_ (.A0(_0237_),
    .A1(_0238_),
    .A2(_0240_),
    .A3(_0239_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit31.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit0.Q ),
    .X(_0241_));
 sky130_fd_sc_hd__mux2_4 _1106_ (.A0(_0241_),
    .A1(_0229_),
    .S(\Inst_LG_LUT4c_frame_config_dffesr.c_I0mux ),
    .X(_0242_));
 sky130_fd_sc_hd__mux4_2 _1107_ (.A0(net23),
    .A1(net106),
    .A2(net138),
    .A3(\Inst_LUT4AB_switch_matrix.JS2BEG4 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit22.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit23.Q ),
    .X(_0243_));
 sky130_fd_sc_hd__mux4_2 _1108_ (.A0(net82),
    .A1(net94),
    .A2(net11),
    .A3(net122),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit23.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit22.Q ),
    .X(_0244_));
 sky130_fd_sc_hd__mux4_1 _1109_ (.A0(net660),
    .A1(net657),
    .A2(net652),
    .A3(net636),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit18.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit19.Q ),
    .X(_0245_));
 sky130_fd_sc_hd__mux4_1 _1110_ (.A0(net646),
    .A1(net627),
    .A2(net642),
    .A3(net623),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit19.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit18.Q ),
    .X(_0246_));
 sky130_fd_sc_hd__mux2_2 _1111_ (.A0(_0245_),
    .A1(_0246_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit20.Q ),
    .X(_0247_));
 sky130_fd_sc_hd__mux4_1 _1112_ (.A0(net60),
    .A1(net68),
    .A2(net5),
    .A3(net13),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit18.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit19.Q ),
    .X(_0248_));
 sky130_fd_sc_hd__and2b_1 _1113_ (.A_N(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit20.Q ),
    .B(_0248_),
    .X(_0249_));
 sky130_fd_sc_hd__mux4_1 _1114_ (.A0(net88),
    .A1(net114),
    .A2(net96),
    .A3(net665),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit19.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit18.Q ),
    .X(_0250_));
 sky130_fd_sc_hd__a21o_1 _1115_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit20.Q ),
    .A2(_0250_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit21.Q ),
    .X(_0251_));
 sky130_fd_sc_hd__o22a_4 _1116_ (.A1(_0575_),
    .A2(_0247_),
    .B1(_0249_),
    .B2(_0251_),
    .X(\Inst_LUT4AB_switch_matrix.JS2BEG6 ));
 sky130_fd_sc_hd__mux4_2 _1117_ (.A0(net18),
    .A1(net129),
    .A2(net101),
    .A3(\Inst_LUT4AB_switch_matrix.JS2BEG6 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit23.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit22.Q ),
    .X(_0252_));
 sky130_fd_sc_hd__mux4_1 _1118_ (.A0(net74),
    .A1(net19),
    .A2(net102),
    .A3(net130),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit22.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit23.Q ),
    .X(_0253_));
 sky130_fd_sc_hd__mux4_2 _1119_ (.A0(_0252_),
    .A1(_0253_),
    .A2(_0244_),
    .A3(_0243_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit3.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit4.Q ),
    .X(_0254_));
 sky130_fd_sc_hd__mux4_2 _1120_ (.A0(net79),
    .A1(net119),
    .A2(net111),
    .A3(\Inst_LUT4AB_switch_matrix.E2BEG4 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit21.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit20.Q ),
    .X(_0255_));
 sky130_fd_sc_hd__mux4_2 _1121_ (.A0(net64),
    .A1(net109),
    .A2(net9),
    .A3(net120),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit21.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit20.Q ),
    .X(_0256_));
 sky130_fd_sc_hd__mux4_2 _1122_ (.A0(net647),
    .A1(net628),
    .A2(net643),
    .A3(net404),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit19.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit18.Q ),
    .X(_0257_));
 sky130_fd_sc_hd__mux4_1 _1123_ (.A0(net661),
    .A1(net658),
    .A2(net653),
    .A3(net638),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit18.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit19.Q ),
    .X(_0258_));
 sky130_fd_sc_hd__mux2_4 _1124_ (.A0(_0258_),
    .A1(_0257_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit20.Q ),
    .X(_0259_));
 sky130_fd_sc_hd__mux4_1 _1125_ (.A0(net86),
    .A1(net88),
    .A2(net96),
    .A3(net665),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit18.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit19.Q ),
    .X(_0260_));
 sky130_fd_sc_hd__mux4_1 _1126_ (.A0(net60),
    .A1(net68),
    .A2(net815),
    .A3(net13),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit18.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit19.Q ),
    .X(_0261_));
 sky130_fd_sc_hd__and2b_1 _1127_ (.A_N(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit20.Q ),
    .B(_0261_),
    .X(_0262_));
 sky130_fd_sc_hd__a211o_1 _1128_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit20.Q ),
    .A2(_0260_),
    .B1(_0262_),
    .C1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit21.Q ),
    .X(_0263_));
 sky130_fd_sc_hd__o21a_4 _1129_ (.A1(_0574_),
    .A2(_0259_),
    .B1(_0263_),
    .X(\Inst_LUT4AB_switch_matrix.E2BEG6 ));
 sky130_fd_sc_hd__mux4_2 _1130_ (.A0(net71),
    .A1(net127),
    .A2(net99),
    .A3(\Inst_LUT4AB_switch_matrix.E2BEG6 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit21.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit20.Q ),
    .X(_0264_));
 sky130_fd_sc_hd__mux4_2 _1131_ (.A0(net72),
    .A1(net17),
    .A2(net100),
    .A3(net128),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit20.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit21.Q ),
    .X(_0265_));
 sky130_fd_sc_hd__mux4_2 _1132_ (.A0(_0264_),
    .A1(_0265_),
    .A2(_0256_),
    .A3(_0255_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit1.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit2.Q ),
    .X(_0266_));
 sky130_fd_sc_hd__or2_4 _1133_ (.A(_0266_),
    .B(_0254_),
    .X(_0267_));
 sky130_fd_sc_hd__nand2_1 _1134_ (.A(_0254_),
    .B(_0266_),
    .Y(_0268_));
 sky130_fd_sc_hd__inv_2 _1135_ (.A(_0268_),
    .Y(_0269_));
 sky130_fd_sc_hd__mux4_1 _1136_ (.A0(_0577_),
    .A1(_0578_),
    .A2(_0579_),
    .A3(_0580_),
    .S0(_0266_),
    .S1(_0254_),
    .X(_0270_));
 sky130_fd_sc_hd__mux4_2 _1137_ (.A0(net81),
    .A1(net117),
    .A2(net22),
    .A3(\Inst_LUT4AB_switch_matrix.JW2BEG4 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit25.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit24.Q ),
    .X(_0271_));
 sky130_fd_sc_hd__mux4_2 _1138_ (.A0(net62),
    .A1(net90),
    .A2(net27),
    .A3(net118),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit25.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit24.Q ),
    .X(_0272_));
 sky130_fd_sc_hd__mux4_1 _1139_ (.A0(net646),
    .A1(net627),
    .A2(net642),
    .A3(net622),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit19.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit18.Q ),
    .X(_0273_));
 sky130_fd_sc_hd__mux4_1 _1140_ (.A0(net662),
    .A1(net656),
    .A2(net652),
    .A3(net636),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit18.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit19.Q ),
    .X(_0274_));
 sky130_fd_sc_hd__mux2_4 _1141_ (.A0(_0274_),
    .A1(_0273_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit20.Q ),
    .X(_0275_));
 sky130_fd_sc_hd__mux4_1 _1142_ (.A0(net86),
    .A1(net88),
    .A2(net96),
    .A3(net665),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit18.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit19.Q ),
    .X(_0276_));
 sky130_fd_sc_hd__mux4_1 _1143_ (.A0(net60),
    .A1(net68),
    .A2(net815),
    .A3(net13),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit18.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit19.Q ),
    .X(_0277_));
 sky130_fd_sc_hd__and2b_1 _1144_ (.A_N(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit20.Q ),
    .B(_0277_),
    .X(_0278_));
 sky130_fd_sc_hd__a21o_1 _1145_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit20.Q ),
    .A2(_0276_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit21.Q ),
    .X(_0279_));
 sky130_fd_sc_hd__o22a_4 _1146_ (.A1(_0275_),
    .A2(_0576_),
    .B1(_0278_),
    .B2(_0279_),
    .X(\Inst_LUT4AB_switch_matrix.JW2BEG6 ));
 sky130_fd_sc_hd__mux4_2 _1147_ (.A0(net69),
    .A1(net14),
    .A2(net125),
    .A3(\Inst_LUT4AB_switch_matrix.JW2BEG6 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit24.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit25.Q ),
    .X(_0280_));
 sky130_fd_sc_hd__mux4_1 _1148_ (.A0(net70),
    .A1(net15),
    .A2(net98),
    .A3(net126),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit24.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit25.Q ),
    .X(_0281_));
 sky130_fd_sc_hd__mux4_2 _1149_ (.A0(_0280_),
    .A1(_0281_),
    .A2(_0272_),
    .A3(_0271_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit5.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit6.Q ),
    .X(_0282_));
 sky130_fd_sc_hd__mux4_1 _1150_ (.A0(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ),
    .A1(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ),
    .A2(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ),
    .A3(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ),
    .S0(_0266_),
    .S1(_0254_),
    .X(_0283_));
 sky130_fd_sc_hd__o21ai_2 _1151_ (.A1(_0283_),
    .A2(_0242_),
    .B1(_0282_),
    .Y(_0284_));
 sky130_fd_sc_hd__a21oi_2 _1152_ (.A1(_0242_),
    .A2(_0270_),
    .B1(_0284_),
    .Y(_0285_));
 sky130_fd_sc_hd__mux4_1 _1153_ (.A0(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ),
    .A1(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ),
    .A2(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ),
    .A3(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ),
    .S0(_0266_),
    .S1(_0254_),
    .X(_0286_));
 sky130_fd_sc_hd__or3b_4 _1154_ (.A(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ),
    .B(_0254_),
    .C_N(_0266_),
    .X(_0287_));
 sky130_fd_sc_hd__or3b_1 _1155_ (.A(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ),
    .B(_0266_),
    .C_N(_0254_),
    .X(_0288_));
 sky130_fd_sc_hd__o22a_1 _1156_ (.A1(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ),
    .A2(_0267_),
    .B1(_0268_),
    .B2(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ),
    .X(_0289_));
 sky130_fd_sc_hd__and3_1 _1157_ (.A(_0287_),
    .B(_0288_),
    .C(_0289_),
    .X(_0290_));
 sky130_fd_sc_hd__mux2_1 _1158_ (.A0(_0286_),
    .A1(_0290_),
    .S(_0242_),
    .X(_0291_));
 sky130_fd_sc_hd__and2b_1 _1159_ (.A_N(_0282_),
    .B(_0291_),
    .X(_0292_));
 sky130_fd_sc_hd__nand2b_1 _1160_ (.A_N(\Inst_LG_LUT4c_frame_config_dffesr.LUT_flop ),
    .B(\Inst_LG_LUT4c_frame_config_dffesr.c_out_mux ),
    .Y(_0293_));
 sky130_fd_sc_hd__o31a_4 _1161_ (.A1(_0292_),
    .A2(_0285_),
    .A3(\Inst_LG_LUT4c_frame_config_dffesr.c_out_mux ),
    .B1(_0293_),
    .X(G));
 sky130_fd_sc_hd__a311o_1 _1162_ (.A1(_0211_),
    .A2(_0204_),
    .A3(_0126_),
    .B1(_0212_),
    .C1(_0269_),
    .X(_0294_));
 sky130_fd_sc_hd__a21o_1 _1163_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit9.Q ),
    .A2(_0238_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit10.Q ),
    .X(_0295_));
 sky130_fd_sc_hd__a21oi_1 _1164_ (.A1(_0581_),
    .A2(_0237_),
    .B1(_0295_),
    .Y(_0296_));
 sky130_fd_sc_hd__nand2_1 _1165_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit9.Q ),
    .B(_0239_),
    .Y(_0297_));
 sky130_fd_sc_hd__nand2_1 _1166_ (.A(_0581_),
    .B(_0240_),
    .Y(_0298_));
 sky130_fd_sc_hd__a311oi_1 _1167_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit10.Q ),
    .A2(_0297_),
    .A3(_0298_),
    .B1(\Inst_LH_LUT4c_frame_config_dffesr.c_I0mux ),
    .C1(_0296_),
    .Y(_0299_));
 sky130_fd_sc_hd__a31o_1 _1168_ (.A1(_0294_),
    .A2(_0267_),
    .A3(\Inst_LH_LUT4c_frame_config_dffesr.c_I0mux ),
    .B1(_0299_),
    .X(_0300_));
 sky130_fd_sc_hd__mux4_2 _1169_ (.A0(_0252_),
    .A1(_0253_),
    .A2(_0244_),
    .A3(_0243_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit13.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit14.Q ),
    .X(_0301_));
 sky130_fd_sc_hd__mux4_2 _1170_ (.A0(_0264_),
    .A1(_0265_),
    .A2(_0256_),
    .A3(_0255_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit11.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit12.Q ),
    .X(_0302_));
 sky130_fd_sc_hd__nand2b_1 _1171_ (.A_N(_0302_),
    .B(_0301_),
    .Y(_0303_));
 sky130_fd_sc_hd__or2_4 _1172_ (.A(_0301_),
    .B(_0302_),
    .X(_0304_));
 sky130_fd_sc_hd__o22a_1 _1173_ (.A1(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ),
    .A2(_0303_),
    .B1(_0304_),
    .B2(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ),
    .X(_0305_));
 sky130_fd_sc_hd__and2_1 _1174_ (.A(_0301_),
    .B(_0302_),
    .X(_0306_));
 sky130_fd_sc_hd__nand2_1 _1175_ (.A(_0301_),
    .B(_0302_),
    .Y(_0307_));
 sky130_fd_sc_hd__nand2b_1 _1176_ (.A_N(_0301_),
    .B(_0302_),
    .Y(_0308_));
 sky130_fd_sc_hd__o22a_1 _1177_ (.A1(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ),
    .A2(_0307_),
    .B1(_0308_),
    .B2(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ),
    .X(_0309_));
 sky130_fd_sc_hd__a21o_1 _1178_ (.A1(_0305_),
    .A2(_0309_),
    .B1(_0300_),
    .X(_0310_));
 sky130_fd_sc_hd__mux4_2 _1179_ (.A0(_0280_),
    .A1(_0281_),
    .A2(_0272_),
    .A3(_0271_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit15.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit16.Q ),
    .X(_0311_));
 sky130_fd_sc_hd__o22a_1 _1180_ (.A1(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ),
    .A2(_0303_),
    .B1(_0304_),
    .B2(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ),
    .X(_0312_));
 sky130_fd_sc_hd__o22a_1 _1181_ (.A1(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ),
    .A2(_0307_),
    .B1(_0308_),
    .B2(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ),
    .X(_0313_));
 sky130_fd_sc_hd__nand2_1 _1182_ (.A(_0312_),
    .B(_0313_),
    .Y(_0314_));
 sky130_fd_sc_hd__a21oi_1 _1183_ (.A1(_0300_),
    .A2(_0314_),
    .B1(_0311_),
    .Y(_0315_));
 sky130_fd_sc_hd__o22a_1 _1184_ (.A1(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ),
    .A2(_0303_),
    .B1(_0307_),
    .B2(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ),
    .X(_0316_));
 sky130_fd_sc_hd__or2_1 _1185_ (.A(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ),
    .B(_0308_),
    .X(_0317_));
 sky130_fd_sc_hd__o211a_1 _1186_ (.A1(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ),
    .A2(_0304_),
    .B1(_0316_),
    .C1(_0317_),
    .X(_0318_));
 sky130_fd_sc_hd__o22a_1 _1187_ (.A1(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ),
    .A2(_0307_),
    .B1(_0308_),
    .B2(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ),
    .X(_0319_));
 sky130_fd_sc_hd__or2_1 _1188_ (.A(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ),
    .B(_0303_),
    .X(_0320_));
 sky130_fd_sc_hd__o211a_1 _1189_ (.A1(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ),
    .A2(_0304_),
    .B1(_0319_),
    .C1(_0320_),
    .X(_0321_));
 sky130_fd_sc_hd__mux2_1 _1190_ (.A0(_0318_),
    .A1(_0321_),
    .S(_0300_),
    .X(_0322_));
 sky130_fd_sc_hd__a22o_1 _1191_ (.A1(_0315_),
    .A2(_0310_),
    .B1(_0322_),
    .B2(_0311_),
    .X(_0323_));
 sky130_fd_sc_hd__mux2_4 _1192_ (.A0(_0323_),
    .A1(\Inst_LH_LUT4c_frame_config_dffesr.LUT_flop ),
    .S(\Inst_LH_LUT4c_frame_config_dffesr.c_out_mux ),
    .X(H));
 sky130_fd_sc_hd__mux2_4 _1193_ (.A0(\Inst_LUT4AB_switch_matrix.JN2BEG6 ),
    .A1(\Inst_LUT4AB_switch_matrix.E2BEG6 ),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit22.Q ),
    .X(_0324_));
 sky130_fd_sc_hd__mux2_1 _1194_ (.A0(\Inst_LUT4AB_switch_matrix.JS2BEG6 ),
    .A1(\Inst_LUT4AB_switch_matrix.JW2BEG6 ),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit22.Q ),
    .X(_0325_));
 sky130_fd_sc_hd__mux2_4 _1195_ (.A0(_0324_),
    .A1(_0325_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit23.Q ),
    .X(_0326_));
 sky130_fd_sc_hd__mux4_2 _1196_ (.A0(\Inst_LUT4AB_switch_matrix.JN2BEG4 ),
    .A1(\Inst_LUT4AB_switch_matrix.JS2BEG4 ),
    .A2(\Inst_LUT4AB_switch_matrix.E2BEG4 ),
    .A3(\Inst_LUT4AB_switch_matrix.JW2BEG4 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit19.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit18.Q ),
    .X(_0327_));
 sky130_fd_sc_hd__mux2_4 _1197_ (.A0(_0326_),
    .A1(net396),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit17.Q ),
    .X(_0328_));
 sky130_fd_sc_hd__mux2_4 _1198_ (.A0(net647),
    .A1(net641),
    .S(_0328_),
    .X(\Inst_LUT4AB_switch_matrix.M_EF ));
 sky130_fd_sc_hd__mux2_1 _1199_ (.A0(_0167_),
    .A1(_0168_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit1.Q ),
    .X(_0329_));
 sky130_fd_sc_hd__mux2_1 _1200_ (.A0(_0159_),
    .A1(_0158_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit1.Q ),
    .X(_0330_));
 sky130_fd_sc_hd__mux2_1 _1201_ (.A0(_0329_),
    .A1(_0330_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit2.Q ),
    .X(_0331_));
 sky130_fd_sc_hd__and2b_1 _1202_ (.A_N(\Inst_LD_LUT4c_frame_config_dffesr.c_I0mux ),
    .B(_0331_),
    .X(_0332_));
 sky130_fd_sc_hd__a31o_1 _1203_ (.A1(\Inst_LD_LUT4c_frame_config_dffesr.c_I0mux ),
    .A2(_0080_),
    .A3(_0083_),
    .B1(_0332_),
    .X(_0333_));
 sky130_fd_sc_hd__nand2b_1 _1204_ (.A_N(_0073_),
    .B(_0054_),
    .Y(_0334_));
 sky130_fd_sc_hd__o22a_1 _1205_ (.A1(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ),
    .A2(_0074_),
    .B1(_0334_),
    .B2(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ),
    .X(_0335_));
 sky130_fd_sc_hd__nand2b_1 _1206_ (.A_N(_0054_),
    .B(_0073_),
    .Y(_0336_));
 sky130_fd_sc_hd__o221a_1 _1207_ (.A1(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ),
    .A2(_0075_),
    .B1(_0336_),
    .B2(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ),
    .C1(_0335_),
    .X(_0337_));
 sky130_fd_sc_hd__mux4_2 _1208_ (.A0(_0191_),
    .A1(_0192_),
    .A2(_0183_),
    .A3(_0182_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit7.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit8.Q ),
    .X(_0338_));
 sky130_fd_sc_hd__o22a_1 _1209_ (.A1(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ),
    .A2(_0334_),
    .B1(_0336_),
    .B2(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ),
    .X(_0339_));
 sky130_fd_sc_hd__o221a_1 _1210_ (.A1(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ),
    .A2(_0074_),
    .B1(_0075_),
    .B2(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ),
    .C1(_0339_),
    .X(_0340_));
 sky130_fd_sc_hd__mux2_1 _1211_ (.A0(_0337_),
    .A1(_0340_),
    .S(_0333_),
    .X(_0341_));
 sky130_fd_sc_hd__o22a_1 _1212_ (.A1(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ),
    .A2(_0075_),
    .B1(_0334_),
    .B2(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ),
    .X(_0342_));
 sky130_fd_sc_hd__o22a_1 _1213_ (.A1(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ),
    .A2(_0074_),
    .B1(_0336_),
    .B2(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ),
    .X(_0343_));
 sky130_fd_sc_hd__nand2_1 _1214_ (.A(_0342_),
    .B(_0343_),
    .Y(_0344_));
 sky130_fd_sc_hd__o22a_1 _1215_ (.A1(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ),
    .A2(_0075_),
    .B1(_0336_),
    .B2(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ),
    .X(_0345_));
 sky130_fd_sc_hd__o22a_1 _1216_ (.A1(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ),
    .A2(_0074_),
    .B1(_0334_),
    .B2(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ),
    .X(_0346_));
 sky130_fd_sc_hd__a21o_1 _1217_ (.A1(_0345_),
    .A2(_0346_),
    .B1(_0333_),
    .X(_0347_));
 sky130_fd_sc_hd__a21oi_1 _1218_ (.A1(_0333_),
    .A2(_0344_),
    .B1(_0338_),
    .Y(_0348_));
 sky130_fd_sc_hd__a22o_1 _1219_ (.A1(_0341_),
    .A2(_0338_),
    .B1(_0347_),
    .B2(_0348_),
    .X(_0349_));
 sky130_fd_sc_hd__mux2_4 _1220_ (.A0(_0349_),
    .A1(\Inst_LD_LUT4c_frame_config_dffesr.LUT_flop ),
    .S(\Inst_LD_LUT4c_frame_config_dffesr.c_out_mux ),
    .X(D));
 sky130_fd_sc_hd__mux2_4 _1221_ (.A0(\Inst_LUT4AB_switch_matrix.JN2BEG5 ),
    .A1(\Inst_LUT4AB_switch_matrix.E2BEG5 ),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit20.Q ),
    .X(_0350_));
 sky130_fd_sc_hd__mux2_4 _1222_ (.A0(\Inst_LUT4AB_switch_matrix.JS2BEG5 ),
    .A1(\Inst_LUT4AB_switch_matrix.JW2BEG5 ),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit20.Q ),
    .X(_0351_));
 sky130_fd_sc_hd__mux2_4 _1223_ (.A0(_0350_),
    .A1(_0351_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit21.Q ),
    .X(_0352_));
 sky130_fd_sc_hd__mux2_4 _1224_ (.A0(_0352_),
    .A1(net396),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit16.Q ),
    .X(_0353_));
 sky130_fd_sc_hd__mux2_4 _1225_ (.A0(net652),
    .A1(net636),
    .S(_0353_),
    .X(_0354_));
 sky130_fd_sc_hd__mux2_4 _1226_ (.A0(net623),
    .A1(_0354_),
    .S(net412),
    .X(_0355_));
 sky130_fd_sc_hd__mux2_4 _1227_ (.A0(_0354_),
    .A1(_0355_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit16.Q ),
    .X(\Inst_LUT4AB_switch_matrix.M_AD ));
 sky130_fd_sc_hd__mux4_1 _1228_ (.A0(net661),
    .A1(net658),
    .A2(net653),
    .A3(net638),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit22.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit23.Q ),
    .X(_0356_));
 sky130_fd_sc_hd__mux4_2 _1229_ (.A0(net647),
    .A1(net633),
    .A2(net643),
    .A3(net414),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit23.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit22.Q ),
    .X(_0357_));
 sky130_fd_sc_hd__mux2_4 _1230_ (.A0(_0356_),
    .A1(_0357_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit24.Q ),
    .X(_0358_));
 sky130_fd_sc_hd__mux4_1 _1231_ (.A0(net57),
    .A1(net61),
    .A2(net2),
    .A3(net6),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit22.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit23.Q ),
    .X(_0359_));
 sky130_fd_sc_hd__nand2b_1 _1232_ (.A_N(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit24.Q ),
    .B(_0359_),
    .Y(_0360_));
 sky130_fd_sc_hd__mux4_1 _1233_ (.A0(net85),
    .A1(net87),
    .A2(net109),
    .A3(net135),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit22.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit23.Q ),
    .X(_0361_));
 sky130_fd_sc_hd__a21oi_1 _1234_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit24.Q ),
    .A2(_0361_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit25.Q ),
    .Y(_0362_));
 sky130_fd_sc_hd__a2bb2o_4 _1235_ (.A1_N(_0583_),
    .A2_N(_0358_),
    .B1(_0360_),
    .B2(_0362_),
    .X(_0363_));
 sky130_fd_sc_hd__inv_6 _1236_ (.A(_0363_),
    .Y(\Inst_LUT4AB_switch_matrix.E2BEG7 ));
 sky130_fd_sc_hd__mux4_1 _1237_ (.A0(net662),
    .A1(net656),
    .A2(net652),
    .A3(net636),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit22.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit23.Q ),
    .X(_0364_));
 sky130_fd_sc_hd__mux4_1 _1238_ (.A0(net646),
    .A1(net631),
    .A2(net641),
    .A3(net432),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit23.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit22.Q ),
    .X(_0365_));
 sky130_fd_sc_hd__mux2_1 _1239_ (.A0(_0364_),
    .A1(_0365_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit24.Q ),
    .X(_0366_));
 sky130_fd_sc_hd__mux4_1 _1240_ (.A0(net57),
    .A1(net61),
    .A2(net2),
    .A3(net24),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit22.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit23.Q ),
    .X(_0367_));
 sky130_fd_sc_hd__and2b_1 _1241_ (.A_N(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit24.Q ),
    .B(_0367_),
    .X(_0368_));
 sky130_fd_sc_hd__mux4_1 _1242_ (.A0(net85),
    .A1(net113),
    .A2(net89),
    .A3(net666),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit23.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit22.Q ),
    .X(_0369_));
 sky130_fd_sc_hd__a21o_1 _1243_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit24.Q ),
    .A2(_0369_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit25.Q ),
    .X(_0370_));
 sky130_fd_sc_hd__o22a_1 _1244_ (.A1(_0582_),
    .A2(_0366_),
    .B1(_0368_),
    .B2(_0370_),
    .X(\Inst_LUT4AB_switch_matrix.JN2BEG7 ));
 sky130_fd_sc_hd__mux4_2 _1245_ (.A0(net646),
    .A1(net631),
    .A2(net641),
    .A3(\Inst_LUT4AB_switch_matrix.M_AB ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit23.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit22.Q ),
    .X(_0371_));
 sky130_fd_sc_hd__mux4_1 _1246_ (.A0(net660),
    .A1(net657),
    .A2(net652),
    .A3(net637),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit22.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit23.Q ),
    .X(_0372_));
 sky130_fd_sc_hd__mux2_4 _1247_ (.A0(_0372_),
    .A1(_0371_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit24.Q ),
    .X(_0373_));
 sky130_fd_sc_hd__mux4_1 _1248_ (.A0(net57),
    .A1(net81),
    .A2(net2),
    .A3(net6),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit22.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit23.Q ),
    .X(_0374_));
 sky130_fd_sc_hd__nand2b_1 _1249_ (.A_N(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit24.Q ),
    .B(_0374_),
    .Y(_0375_));
 sky130_fd_sc_hd__mux4_1 _1250_ (.A0(net85),
    .A1(net87),
    .A2(net89),
    .A3(net113),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit22.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit23.Q ),
    .X(_0376_));
 sky130_fd_sc_hd__a21oi_1 _1251_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit24.Q ),
    .A2(_0376_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit25.Q ),
    .Y(_0377_));
 sky130_fd_sc_hd__a2bb2o_4 _1252_ (.A1_N(_0585_),
    .A2_N(_0373_),
    .B1(_0375_),
    .B2(_0377_),
    .X(_0378_));
 sky130_fd_sc_hd__inv_1 _1253_ (.A(_0378_),
    .Y(\Inst_LUT4AB_switch_matrix.JW2BEG7 ));
 sky130_fd_sc_hd__mux4_2 _1254_ (.A0(net646),
    .A1(net631),
    .A2(net641),
    .A3(\Inst_LUT4AB_switch_matrix.M_AD ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit23.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit22.Q ),
    .X(_0379_));
 sky130_fd_sc_hd__mux4_1 _1255_ (.A0(net660),
    .A1(net657),
    .A2(net652),
    .A3(net637),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit22.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit23.Q ),
    .X(_0380_));
 sky130_fd_sc_hd__mux2_4 _1256_ (.A0(_0380_),
    .A1(_0379_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit24.Q ),
    .X(_0381_));
 sky130_fd_sc_hd__mux4_1 _1257_ (.A0(net57),
    .A1(net61),
    .A2(net2),
    .A3(net6),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit22.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit23.Q ),
    .X(_0382_));
 sky130_fd_sc_hd__and2b_1 _1258_ (.A_N(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit24.Q ),
    .B(_0382_),
    .X(_0383_));
 sky130_fd_sc_hd__mux4_1 _1259_ (.A0(net85),
    .A1(net113),
    .A2(net89),
    .A3(net115),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit23.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit22.Q ),
    .X(_0384_));
 sky130_fd_sc_hd__a21o_1 _1260_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit24.Q ),
    .A2(_0384_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit25.Q ),
    .X(_0385_));
 sky130_fd_sc_hd__o22a_1 _1261_ (.A1(_0381_),
    .A2(_0584_),
    .B1(_0383_),
    .B2(_0385_),
    .X(\Inst_LUT4AB_switch_matrix.JS2BEG7 ));
 sky130_fd_sc_hd__nand2_2 _1262_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit24.Q ),
    .B(_0378_),
    .Y(_0386_));
 sky130_fd_sc_hd__o211a_1 _1263_ (.A1(\Inst_LUT4AB_switch_matrix.JS2BEG7 ),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit24.Q ),
    .B1(_0386_),
    .C1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit25.Q ),
    .X(_0387_));
 sky130_fd_sc_hd__mux2_1 _1264_ (.A0(\Inst_LUT4AB_switch_matrix.JN2BEG7 ),
    .A1(\Inst_LUT4AB_switch_matrix.E2BEG7 ),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit24.Q ),
    .X(_0388_));
 sky130_fd_sc_hd__a21oi_2 _1265_ (.A1(_0586_),
    .A2(_0388_),
    .B1(_0387_),
    .Y(_0389_));
 sky130_fd_sc_hd__inv_2 _1266_ (.A(_0389_),
    .Y(_0390_));
 sky130_fd_sc_hd__mux2_4 _1267_ (.A0(_0390_),
    .A1(net412),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit17.Q ),
    .X(_0391_));
 sky130_fd_sc_hd__mux2_4 _1268_ (.A0(_0391_),
    .A1(_0328_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit16.Q ),
    .X(_0392_));
 sky130_fd_sc_hd__mux2_4 _1269_ (.A0(net632),
    .A1(net627),
    .S(_0392_),
    .X(_0393_));
 sky130_fd_sc_hd__mux2_4 _1270_ (.A0(net432),
    .A1(_0393_),
    .S(_0391_),
    .X(_0394_));
 sky130_fd_sc_hd__mux2_4 _1271_ (.A0(_0393_),
    .A1(_0394_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit16.Q ),
    .X(_0395_));
 sky130_fd_sc_hd__mux2_4 _1272_ (.A0(_0355_),
    .A1(_0394_),
    .S(_0390_),
    .X(_0396_));
 sky130_fd_sc_hd__mux2_4 _1273_ (.A0(_0395_),
    .A1(_0396_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit17.Q ),
    .X(\Inst_LUT4AB_switch_matrix.M_AH ));
 sky130_fd_sc_hd__mux2_4 _1274_ (.A0(net660),
    .A1(net656),
    .S(net407),
    .X(\Inst_LUT4AB_switch_matrix.M_AB ));
 sky130_fd_sc_hd__mux4_1 _1275_ (.A0(net639),
    .A1(net629),
    .A2(net624),
    .A3(net397),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit26.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit27.Q ),
    .X(_0397_));
 sky130_fd_sc_hd__or2_1 _1276_ (.A(_0587_),
    .B(_0397_),
    .X(_0398_));
 sky130_fd_sc_hd__mux4_1 _1277_ (.A0(net654),
    .A1(net634),
    .A2(net649),
    .A3(net644),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit27.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit26.Q ),
    .X(_0399_));
 sky130_fd_sc_hd__o21a_1 _1278_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit28.Q ),
    .A2(_0399_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit29.Q ),
    .X(_0400_));
 sky130_fd_sc_hd__mux4_1 _1279_ (.A0(net60),
    .A1(net7),
    .A2(net62),
    .A3(net813),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit27.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit26.Q ),
    .X(_0401_));
 sky130_fd_sc_hd__mux4_1 _1280_ (.A0(net90),
    .A1(net118),
    .A2(net106),
    .A3(net134),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit27.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit26.Q ),
    .X(_0402_));
 sky130_fd_sc_hd__mux2_1 _1281_ (.A0(_0401_),
    .A1(_0402_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit28.Q ),
    .X(_0403_));
 sky130_fd_sc_hd__a22o_1 _1282_ (.A1(_0398_),
    .A2(_0400_),
    .B1(_0403_),
    .B2(_0588_),
    .X(\Inst_LUT4AB_switch_matrix.JW2BEG0 ));
 sky130_fd_sc_hd__mux4_1 _1283_ (.A0(net430),
    .A1(net411),
    .A2(net649),
    .A3(net644),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit27.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit26.Q ),
    .X(_0404_));
 sky130_fd_sc_hd__mux4_2 _1284_ (.A0(net639),
    .A1(net629),
    .A2(net624),
    .A3(net416),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit26.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit27.Q ),
    .X(_0405_));
 sky130_fd_sc_hd__or2_4 _1285_ (.A(_0405_),
    .B(_0589_),
    .X(_0406_));
 sky130_fd_sc_hd__o21a_1 _1286_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit28.Q ),
    .A2(_0404_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit29.Q ),
    .X(_0407_));
 sky130_fd_sc_hd__mux4_1 _1287_ (.A0(net82),
    .A1(net7),
    .A2(net815),
    .A3(net813),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit27.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit26.Q ),
    .X(_0408_));
 sky130_fd_sc_hd__mux4_1 _1288_ (.A0(net90),
    .A1(net118),
    .A2(net106),
    .A3(net134),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit27.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit26.Q ),
    .X(_0409_));
 sky130_fd_sc_hd__mux2_1 _1289_ (.A0(_0408_),
    .A1(_0409_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit28.Q ),
    .X(_0410_));
 sky130_fd_sc_hd__a22o_4 _1290_ (.A1(_0407_),
    .A2(_0406_),
    .B1(_0410_),
    .B2(_0590_),
    .X(\Inst_LUT4AB_switch_matrix.JS2BEG0 ));
 sky130_fd_sc_hd__mux4_1 _1291_ (.A0(net654),
    .A1(net411),
    .A2(net649),
    .A3(net645),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit27.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit26.Q ),
    .X(_0411_));
 sky130_fd_sc_hd__or2_1 _1292_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit28.Q ),
    .B(_0411_),
    .X(_0412_));
 sky130_fd_sc_hd__mux4_1 _1293_ (.A0(net639),
    .A1(net629),
    .A2(net624),
    .A3(net622),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit26.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit27.Q ),
    .X(_0413_));
 sky130_fd_sc_hd__o21a_1 _1294_ (.A1(_0591_),
    .A2(_0413_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit29.Q ),
    .X(_0414_));
 sky130_fd_sc_hd__mux4_1 _1295_ (.A0(net813),
    .A1(net118),
    .A2(net90),
    .A3(net134),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit27.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit26.Q ),
    .X(_0415_));
 sky130_fd_sc_hd__mux4_1 _1296_ (.A0(net60),
    .A1(net62),
    .A2(net78),
    .A3(net25),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit26.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit27.Q ),
    .X(_0416_));
 sky130_fd_sc_hd__mux2_1 _1297_ (.A0(_0415_),
    .A1(_0416_),
    .S(_0591_),
    .X(_0417_));
 sky130_fd_sc_hd__a22o_1 _1298_ (.A1(_0412_),
    .A2(_0414_),
    .B1(_0417_),
    .B2(_0592_),
    .X(\Inst_LUT4AB_switch_matrix.E2BEG0 ));
 sky130_fd_sc_hd__mux4_1 _1299_ (.A0(net654),
    .A1(net634),
    .A2(net649),
    .A3(net645),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit27.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit26.Q ),
    .X(_0418_));
 sky130_fd_sc_hd__or2_1 _1300_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit28.Q ),
    .B(_0418_),
    .X(_0419_));
 sky130_fd_sc_hd__mux4_1 _1301_ (.A0(net639),
    .A1(net630),
    .A2(net625),
    .A3(net623),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit26.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit27.Q ),
    .X(_0420_));
 sky130_fd_sc_hd__o21a_1 _1302_ (.A1(_0593_),
    .A2(_0420_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit29.Q ),
    .X(_0421_));
 sky130_fd_sc_hd__mux4_1 _1303_ (.A0(net813),
    .A1(net110),
    .A2(net118),
    .A3(net134),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit26.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit27.Q ),
    .X(_0422_));
 sky130_fd_sc_hd__mux4_1 _1304_ (.A0(net62),
    .A1(net815),
    .A2(net78),
    .A3(net7),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit27.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit26.Q ),
    .X(_0423_));
 sky130_fd_sc_hd__mux2_1 _1305_ (.A0(_0422_),
    .A1(_0423_),
    .S(_0593_),
    .X(_0424_));
 sky130_fd_sc_hd__a22o_1 _1306_ (.A1(_0419_),
    .A2(_0421_),
    .B1(_0424_),
    .B2(_0594_),
    .X(\Inst_LUT4AB_switch_matrix.JN2BEG0 ));
 sky130_fd_sc_hd__mux4_2 _1307_ (.A0(_0652_),
    .A1(_0071_),
    .A2(_0107_),
    .A3(_0252_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit30.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit31.Q ),
    .X(_0425_));
 sky130_fd_sc_hd__mux4_1 _1308_ (.A0(net631),
    .A1(net627),
    .A2(net397),
    .A3(net432),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit30.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit31.Q ),
    .X(_0426_));
 sky130_fd_sc_hd__mux2_4 _1309_ (.A0(_0426_),
    .A1(_0425_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit0.Q ),
    .X(_0427_));
 sky130_fd_sc_hd__mux4_1 _1310_ (.A0(net4),
    .A1(net666),
    .A2(net660),
    .A3(net430),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit30.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit31.Q ),
    .X(_0428_));
 sky130_fd_sc_hd__or2_1 _1311_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit0.Q ),
    .B(_0428_),
    .X(_0429_));
 sky130_fd_sc_hd__mux4_1 _1312_ (.A0(net650),
    .A1(net411),
    .A2(net646),
    .A3(net641),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit30.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit31.Q ),
    .X(_0430_));
 sky130_fd_sc_hd__inv_1 _1313_ (.A(_0430_),
    .Y(_0431_));
 sky130_fd_sc_hd__a21oi_1 _1314_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit0.Q ),
    .A2(_0431_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit1.Q ),
    .Y(_0432_));
 sky130_fd_sc_hd__a22o_1 _1315_ (.A1(_0427_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit1.Q ),
    .B1(_0429_),
    .B2(_0432_),
    .X(\Inst_LUT4AB_switch_matrix.W6BEG1 ));
 sky130_fd_sc_hd__mux4_1 _1316_ (.A0(net815),
    .A1(net665),
    .A2(net426),
    .A3(net430),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit26.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit27.Q ),
    .X(_0433_));
 sky130_fd_sc_hd__mux2_1 _1317_ (.A0(net645),
    .A1(net640),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit26.Q ),
    .X(_0434_));
 sky130_fd_sc_hd__mux2_1 _1318_ (.A0(net650),
    .A1(net411),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit26.Q ),
    .X(_0435_));
 sky130_fd_sc_hd__and2b_1 _1319_ (.A_N(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit27.Q ),
    .B(_0435_),
    .X(_0436_));
 sky130_fd_sc_hd__a21bo_1 _1320_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit27.Q ),
    .A2(_0434_),
    .B1_N(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit28.Q ),
    .X(_0437_));
 sky130_fd_sc_hd__o22a_1 _1321_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit28.Q ),
    .A2(_0433_),
    .B1(_0436_),
    .B2(_0437_),
    .X(_0438_));
 sky130_fd_sc_hd__mux4_1 _1322_ (.A0(_0617_),
    .A1(_0053_),
    .A2(_0120_),
    .A3(net664),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit26.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit27.Q ),
    .X(_0439_));
 sky130_fd_sc_hd__mux4_2 _1323_ (.A0(net399),
    .A1(net625),
    .A2(net623),
    .A3(net406),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit26.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit27.Q ),
    .X(_0440_));
 sky130_fd_sc_hd__mux2_4 _1324_ (.A0(_0440_),
    .A1(_0439_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit28.Q ),
    .X(_0441_));
 sky130_fd_sc_hd__mux2_4 _1325_ (.A0(_0438_),
    .A1(_0441_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit29.Q ),
    .X(\Inst_LUT4AB_switch_matrix.W6BEG0 ));
 sky130_fd_sc_hd__mux4_1 _1326_ (.A0(net58),
    .A1(net86),
    .A2(net114),
    .A3(net411),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit23.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit24.Q ),
    .X(_0442_));
 sky130_fd_sc_hd__mux4_1 _1327_ (.A0(net645),
    .A1(net431),
    .A2(_0252_),
    .A3(_0662_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit23.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit24.Q ),
    .X(_0443_));
 sky130_fd_sc_hd__mux2_4 _1328_ (.A0(_0442_),
    .A1(_0443_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit25.Q ),
    .X(\Inst_LUT4AB_switch_matrix.WW4BEG3 ));
 sky130_fd_sc_hd__mux4_1 _1329_ (.A0(net650),
    .A1(_0120_),
    .A2(net664),
    .A3(_0063_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit20.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit21.Q ),
    .X(_0444_));
 sky130_fd_sc_hd__mux4_1 _1330_ (.A0(net57),
    .A1(net113),
    .A2(net85),
    .A3(net430),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit21.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit20.Q ),
    .X(_0445_));
 sky130_fd_sc_hd__mux2_1 _1331_ (.A0(_0445_),
    .A1(_0444_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit22.Q ),
    .X(\Inst_LUT4AB_switch_matrix.WW4BEG2 ));
 sky130_fd_sc_hd__mux4_2 _1332_ (.A0(net627),
    .A1(_0652_),
    .A2(_0071_),
    .A3(_0099_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit17.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit18.Q ),
    .X(_0446_));
 sky130_fd_sc_hd__mux4_1 _1333_ (.A0(net60),
    .A1(net88),
    .A2(net665),
    .A3(net660),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit17.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit18.Q ),
    .X(_0447_));
 sky130_fd_sc_hd__mux2_4 _1334_ (.A0(_0447_),
    .A1(_0446_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit19.Q ),
    .X(\Inst_LUT4AB_switch_matrix.WW4BEG1 ));
 sky130_fd_sc_hd__mux4_1 _1335_ (.A0(net631),
    .A1(_0617_),
    .A2(_0053_),
    .A3(_0244_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit15.Q ),
    .X(_0448_));
 sky130_fd_sc_hd__nand2b_1 _1336_ (.A_N(net87),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit14.Q ),
    .Y(_0449_));
 sky130_fd_sc_hd__o21ba_1 _1337_ (.A1(net59),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit14.Q ),
    .B1_N(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit15.Q ),
    .X(_0450_));
 sky130_fd_sc_hd__mux2_1 _1338_ (.A0(net666),
    .A1(net642),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit14.Q ),
    .X(_0451_));
 sky130_fd_sc_hd__a221o_1 _1339_ (.A1(_0449_),
    .A2(_0450_),
    .B1(_0451_),
    .B2(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit15.Q ),
    .C1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit16.Q ),
    .X(_0452_));
 sky130_fd_sc_hd__o21a_1 _1340_ (.A1(_0595_),
    .A2(_0448_),
    .B1(_0452_),
    .X(\Inst_LUT4AB_switch_matrix.WW4BEG0 ));
 sky130_fd_sc_hd__mux4_1 _1341_ (.A0(net648),
    .A1(net431),
    .A2(_0252_),
    .A3(_0683_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit3.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit4.Q ),
    .X(_0453_));
 sky130_fd_sc_hd__mux4_1 _1342_ (.A0(net58),
    .A1(net3),
    .A2(net114),
    .A3(net635),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit3.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit4.Q ),
    .X(_0454_));
 sky130_fd_sc_hd__mux2_4 _1343_ (.A0(_0454_),
    .A1(_0453_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit5.Q ),
    .X(\Inst_LUT4AB_switch_matrix.SS4BEG3 ));
 sky130_fd_sc_hd__mux4_1 _1344_ (.A0(net651),
    .A1(_0120_),
    .A2(net664),
    .A3(_0183_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit0.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit1.Q ),
    .X(_0455_));
 sky130_fd_sc_hd__mux4_1 _1345_ (.A0(net57),
    .A1(net113),
    .A2(net2),
    .A3(net655),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit1.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit0.Q ),
    .X(_0456_));
 sky130_fd_sc_hd__mux2_4 _1346_ (.A0(_0456_),
    .A1(_0455_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit2.Q ),
    .X(\Inst_LUT4AB_switch_matrix.SS4BEG2 ));
 sky130_fd_sc_hd__mux4_1 _1347_ (.A0(net60),
    .A1(net815),
    .A2(net665),
    .A3(net663),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit29.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit30.Q ),
    .X(_0457_));
 sky130_fd_sc_hd__mux2_4 _1348_ (.A0(_0071_),
    .A1(_0130_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit29.Q ),
    .X(_0458_));
 sky130_fd_sc_hd__mux2_1 _1349_ (.A0(net626),
    .A1(_0652_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit29.Q ),
    .X(_0459_));
 sky130_fd_sc_hd__and2b_1 _1350_ (.A_N(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit30.Q ),
    .B(_0459_),
    .X(_0460_));
 sky130_fd_sc_hd__a21bo_1 _1351_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit30.Q ),
    .A2(_0458_),
    .B1_N(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit31.Q ),
    .X(_0461_));
 sky130_fd_sc_hd__o22a_1 _1352_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit31.Q ),
    .A2(_0457_),
    .B1(_0460_),
    .B2(_0461_),
    .X(\Inst_LUT4AB_switch_matrix.SS4BEG1 ));
 sky130_fd_sc_hd__mux4_1 _1353_ (.A0(net399),
    .A1(_0617_),
    .A2(_0053_),
    .A3(_0272_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit26.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit27.Q ),
    .X(_0462_));
 sky130_fd_sc_hd__nand2b_1 _1354_ (.A_N(net816),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit26.Q ),
    .Y(_0463_));
 sky130_fd_sc_hd__o21ba_1 _1355_ (.A1(net59),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit26.Q ),
    .B1_N(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit27.Q ),
    .X(_0464_));
 sky130_fd_sc_hd__mux2_1 _1356_ (.A0(net666),
    .A1(net424),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit26.Q ),
    .X(_0465_));
 sky130_fd_sc_hd__a221o_1 _1357_ (.A1(_0463_),
    .A2(_0464_),
    .B1(_0465_),
    .B2(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit27.Q ),
    .C1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit28.Q ),
    .X(_0466_));
 sky130_fd_sc_hd__o21a_1 _1358_ (.A1(_0596_),
    .A2(_0462_),
    .B1(_0466_),
    .X(\Inst_LUT4AB_switch_matrix.SS4BEG0 ));
 sky130_fd_sc_hd__mux4_2 _1359_ (.A0(_0652_),
    .A1(_0071_),
    .A2(net431),
    .A3(_0252_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit7.Q ),
    .X(_0467_));
 sky130_fd_sc_hd__mux4_1 _1360_ (.A0(net413),
    .A1(net410),
    .A2(net397),
    .A3(net432),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit7.Q ),
    .X(_0468_));
 sky130_fd_sc_hd__mux2_4 _1361_ (.A0(_0468_),
    .A1(_0467_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit8.Q ),
    .X(_0469_));
 sky130_fd_sc_hd__mux4_1 _1362_ (.A0(net816),
    .A1(net666),
    .A2(net661),
    .A3(net658),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit7.Q ),
    .X(_0470_));
 sky130_fd_sc_hd__or2_1 _1363_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit8.Q ),
    .B(_0470_),
    .X(_0471_));
 sky130_fd_sc_hd__mux4_1 _1364_ (.A0(net653),
    .A1(net638),
    .A2(net647),
    .A3(net642),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit7.Q ),
    .X(_0472_));
 sky130_fd_sc_hd__inv_1 _1365_ (.A(_0472_),
    .Y(_0473_));
 sky130_fd_sc_hd__a21oi_1 _1366_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit8.Q ),
    .A2(_0473_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit9.Q ),
    .Y(_0474_));
 sky130_fd_sc_hd__a22o_1 _1367_ (.A1(_0469_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit9.Q ),
    .B1(_0471_),
    .B2(_0474_),
    .X(\Inst_LUT4AB_switch_matrix.E6BEG1 ));
 sky130_fd_sc_hd__mux4_1 _1368_ (.A0(net815),
    .A1(net665),
    .A2(net661),
    .A3(net658),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit3.Q ),
    .X(_0475_));
 sky130_fd_sc_hd__mux2_1 _1369_ (.A0(net647),
    .A1(net642),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit2.Q ),
    .X(_0476_));
 sky130_fd_sc_hd__mux2_1 _1370_ (.A0(net653),
    .A1(net638),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit2.Q ),
    .X(_0477_));
 sky130_fd_sc_hd__and2b_1 _1371_ (.A_N(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit3.Q ),
    .B(_0477_),
    .X(_0478_));
 sky130_fd_sc_hd__a21bo_1 _1372_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit3.Q ),
    .A2(_0476_),
    .B1_N(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit4.Q ),
    .X(_0479_));
 sky130_fd_sc_hd__o22a_1 _1373_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit4.Q ),
    .A2(_0475_),
    .B1(_0478_),
    .B2(_0479_),
    .X(_0480_));
 sky130_fd_sc_hd__mux4_1 _1374_ (.A0(_0617_),
    .A1(_0053_),
    .A2(_0120_),
    .A3(net664),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit3.Q ),
    .X(_0481_));
 sky130_fd_sc_hd__mux4_2 _1375_ (.A0(net413),
    .A1(net628),
    .A2(net623),
    .A3(net427),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit3.Q ),
    .X(_0482_));
 sky130_fd_sc_hd__mux2_4 _1376_ (.A0(_0482_),
    .A1(_0481_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit4.Q ),
    .X(_0483_));
 sky130_fd_sc_hd__mux2_4 _1377_ (.A0(_0480_),
    .A1(_0483_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit5.Q ),
    .X(\Inst_LUT4AB_switch_matrix.E6BEG0 ));
 sky130_fd_sc_hd__mux4_1 _1378_ (.A0(net58),
    .A1(net3),
    .A2(net86),
    .A3(net638),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit31.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit0.Q ),
    .X(_0484_));
 sky130_fd_sc_hd__mux4_1 _1379_ (.A0(net647),
    .A1(net431),
    .A2(_0252_),
    .A3(_0640_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit31.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit0.Q ),
    .X(_0485_));
 sky130_fd_sc_hd__mux2_4 _1380_ (.A0(_0484_),
    .A1(_0485_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit1.Q ),
    .X(\Inst_LUT4AB_switch_matrix.EE4BEG3 ));
 sky130_fd_sc_hd__mux4_1 _1381_ (.A0(net653),
    .A1(_0120_),
    .A2(net664),
    .A3(_0159_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit28.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit29.Q ),
    .X(_0486_));
 sky130_fd_sc_hd__mux4_1 _1382_ (.A0(net57),
    .A1(net85),
    .A2(net2),
    .A3(net658),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit29.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit28.Q ),
    .X(_0487_));
 sky130_fd_sc_hd__mux2_1 _1383_ (.A0(_0487_),
    .A1(_0486_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit30.Q ),
    .X(\Inst_LUT4AB_switch_matrix.EE4BEG2 ));
 sky130_fd_sc_hd__mux4_1 _1384_ (.A0(net60),
    .A1(net815),
    .A2(net88),
    .A3(net661),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit25.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit26.Q ),
    .X(_0488_));
 sky130_fd_sc_hd__mux2_4 _1385_ (.A0(_0071_),
    .A1(_0095_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit25.Q ),
    .X(_0489_));
 sky130_fd_sc_hd__mux2_1 _1386_ (.A0(net410),
    .A1(_0652_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit25.Q ),
    .X(_0490_));
 sky130_fd_sc_hd__and2b_1 _1387_ (.A_N(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit26.Q ),
    .B(_0490_),
    .X(_0491_));
 sky130_fd_sc_hd__a21bo_1 _1388_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit26.Q ),
    .A2(_0489_),
    .B1_N(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit27.Q ),
    .X(_0492_));
 sky130_fd_sc_hd__o22a_4 _1389_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit27.Q ),
    .A2(_0488_),
    .B1(_0491_),
    .B2(_0492_),
    .X(\Inst_LUT4AB_switch_matrix.EE4BEG1 ));
 sky130_fd_sc_hd__mux4_1 _1390_ (.A0(net413),
    .A1(_0617_),
    .A2(_0053_),
    .A3(_0240_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit22.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit23.Q ),
    .X(_0493_));
 sky130_fd_sc_hd__mux4_1 _1391_ (.A0(net59),
    .A1(net87),
    .A2(net816),
    .A3(net642),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit23.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit22.Q ),
    .X(_0494_));
 sky130_fd_sc_hd__mux2_1 _1392_ (.A0(_0494_),
    .A1(_0493_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit24.Q ),
    .X(\Inst_LUT4AB_switch_matrix.EE4BEG0 ));
 sky130_fd_sc_hd__mux4_1 _1393_ (.A0(net58),
    .A1(net3),
    .A2(net114),
    .A3(net638),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit11.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit12.Q ),
    .X(_0495_));
 sky130_fd_sc_hd__mux4_2 _1394_ (.A0(net647),
    .A1(net431),
    .A2(_0252_),
    .A3(_0606_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit11.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit12.Q ),
    .X(_0496_));
 sky130_fd_sc_hd__mux2_4 _1395_ (.A0(_0495_),
    .A1(_0496_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit13.Q ),
    .X(\Inst_LUT4AB_switch_matrix.NN4BEG3 ));
 sky130_fd_sc_hd__mux4_1 _1396_ (.A0(net653),
    .A1(_0120_),
    .A2(net664),
    .A3(_0044_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit8.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit9.Q ),
    .X(_0497_));
 sky130_fd_sc_hd__mux4_1 _1397_ (.A0(net57),
    .A1(net113),
    .A2(net2),
    .A3(net658),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit9.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit8.Q ),
    .X(_0498_));
 sky130_fd_sc_hd__mux2_1 _1398_ (.A0(_0498_),
    .A1(_0497_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit10.Q ),
    .X(\Inst_LUT4AB_switch_matrix.NN4BEG2 ));
 sky130_fd_sc_hd__mux4_1 _1399_ (.A0(net60),
    .A1(net815),
    .A2(net665),
    .A3(net661),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit5.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit6.Q ),
    .X(_0499_));
 sky130_fd_sc_hd__mux2_1 _1400_ (.A0(net410),
    .A1(_0652_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit5.Q ),
    .X(_0500_));
 sky130_fd_sc_hd__and2b_1 _1401_ (.A_N(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit6.Q ),
    .B(_0500_),
    .X(_0501_));
 sky130_fd_sc_hd__mux2_4 _1402_ (.A0(_0071_),
    .A1(_0111_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit5.Q ),
    .X(_0502_));
 sky130_fd_sc_hd__a21bo_1 _1403_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit6.Q ),
    .A2(_0502_),
    .B1_N(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit7.Q ),
    .X(_0503_));
 sky130_fd_sc_hd__o22a_1 _1404_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit7.Q ),
    .A2(_0499_),
    .B1(_0501_),
    .B2(_0503_),
    .X(\Inst_LUT4AB_switch_matrix.NN4BEG1 ));
 sky130_fd_sc_hd__mux4_1 _1405_ (.A0(net413),
    .A1(_0617_),
    .A2(_0053_),
    .A3(_0256_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit3.Q ),
    .X(_0504_));
 sky130_fd_sc_hd__mux4_1 _1406_ (.A0(net59),
    .A1(net666),
    .A2(net816),
    .A3(net642),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit3.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit2.Q ),
    .X(_0505_));
 sky130_fd_sc_hd__mux2_1 _1407_ (.A0(_0505_),
    .A1(_0504_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit4.Q ),
    .X(\Inst_LUT4AB_switch_matrix.NN4BEG0 ));
 sky130_fd_sc_hd__mux4_2 _1408_ (.A0(net663),
    .A1(_0653_),
    .A2(\Inst_LUT4AB_switch_matrix.JS2BEG2 ),
    .A3(_0639_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit12.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit13.Q ),
    .X(\Inst_LUT4AB_switch_matrix.W1BEG3 ));
 sky130_fd_sc_hd__mux4_2 _1409_ (.A0(net624),
    .A1(\Inst_LUT4AB_switch_matrix.JS2BEG1 ),
    .A2(net664),
    .A3(_0271_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit11.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit10.Q ),
    .X(\Inst_LUT4AB_switch_matrix.W1BEG2 ));
 sky130_fd_sc_hd__mux4_2 _1410_ (.A0(net629),
    .A1(_0093_),
    .A2(\Inst_LUT4AB_switch_matrix.JS2BEG0 ),
    .A3(_0098_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit8.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit9.Q ),
    .X(\Inst_LUT4AB_switch_matrix.W1BEG1 ));
 sky130_fd_sc_hd__mux4_1 _1411_ (.A0(net639),
    .A1(\Inst_LUT4AB_switch_matrix.JS2BEG3 ),
    .A2(_0192_),
    .A3(_0043_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit7.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit6.Q ),
    .X(\Inst_LUT4AB_switch_matrix.W1BEG0 ));
 sky130_fd_sc_hd__mux4_1 _1412_ (.A0(net90),
    .A1(net105),
    .A2(net133),
    .A3(net635),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit24.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit25.Q ),
    .X(\Inst_LUT4AB_switch_matrix.S4BEG3 ));
 sky130_fd_sc_hd__mux4_1 _1413_ (.A0(net89),
    .A1(net134),
    .A2(net108),
    .A3(net651),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit23.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit22.Q ),
    .X(\Inst_LUT4AB_switch_matrix.S4BEG2 ));
 sky130_fd_sc_hd__mux4_1 _1414_ (.A0(net814),
    .A1(net107),
    .A2(net92),
    .A3(net655),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit21.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit20.Q ),
    .X(\Inst_LUT4AB_switch_matrix.S4BEG1 ));
 sky130_fd_sc_hd__mux4_1 _1415_ (.A0(net813),
    .A1(net106),
    .A2(net91),
    .A3(net663),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit19.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit18.Q ),
    .X(\Inst_LUT4AB_switch_matrix.S4BEG0 ));
 sky130_fd_sc_hd__mux4_2 _1416_ (.A0(net626),
    .A1(_0653_),
    .A2(\Inst_LUT4AB_switch_matrix.E2BEG2 ),
    .A3(_0639_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit16.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit17.Q ),
    .X(\Inst_LUT4AB_switch_matrix.S1BEG3 ));
 sky130_fd_sc_hd__mux4_2 _1417_ (.A0(net399),
    .A1(\Inst_LUT4AB_switch_matrix.E2BEG1 ),
    .A2(net664),
    .A3(_0271_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit15.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit14.Q ),
    .X(\Inst_LUT4AB_switch_matrix.S1BEG2 ));
 sky130_fd_sc_hd__mux4_1 _1418_ (.A0(net424),
    .A1(_0093_),
    .A2(\Inst_LUT4AB_switch_matrix.E2BEG0 ),
    .A3(_0098_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit12.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit13.Q ),
    .X(\Inst_LUT4AB_switch_matrix.S1BEG1 ));
 sky130_fd_sc_hd__mux4_2 _1419_ (.A0(net644),
    .A1(\Inst_LUT4AB_switch_matrix.E2BEG3 ),
    .A2(_0192_),
    .A3(_0043_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit11.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit10.Q ),
    .X(\Inst_LUT4AB_switch_matrix.S1BEG0 ));
 sky130_fd_sc_hd__mux4_2 _1420_ (.A0(net399),
    .A1(_0653_),
    .A2(\Inst_LUT4AB_switch_matrix.JN2BEG2 ),
    .A3(_0639_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit20.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit21.Q ),
    .X(\Inst_LUT4AB_switch_matrix.E1BEG3 ));
 sky130_fd_sc_hd__mux4_2 _1421_ (.A0(net424),
    .A1(\Inst_LUT4AB_switch_matrix.JN2BEG1 ),
    .A2(net664),
    .A3(_0271_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit19.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit18.Q ),
    .X(\Inst_LUT4AB_switch_matrix.E1BEG2 ));
 sky130_fd_sc_hd__mux4_1 _1422_ (.A0(net645),
    .A1(_0093_),
    .A2(\Inst_LUT4AB_switch_matrix.JN2BEG0 ),
    .A3(_0098_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit16.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit17.Q ),
    .X(\Inst_LUT4AB_switch_matrix.E1BEG1 ));
 sky130_fd_sc_hd__mux4_2 _1423_ (.A0(net635),
    .A1(\Inst_LUT4AB_switch_matrix.JN2BEG3 ),
    .A2(_0192_),
    .A3(_0043_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit15.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit14.Q ),
    .X(\Inst_LUT4AB_switch_matrix.E1BEG0 ));
 sky130_fd_sc_hd__mux4_1 _1424_ (.A0(net62),
    .A1(net133),
    .A2(net77),
    .A3(net625),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit1.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit0.Q ),
    .X(\Inst_LUT4AB_switch_matrix.N4BEG3 ));
 sky130_fd_sc_hd__mux4_1 _1425_ (.A0(net61),
    .A1(net80),
    .A2(net134),
    .A3(net632),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit30.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit31.Q ),
    .X(\Inst_LUT4AB_switch_matrix.N4BEG2 ));
 sky130_fd_sc_hd__mux4_2 _1426_ (.A0(net64),
    .A1(net79),
    .A2(net22),
    .A3(net641),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit28.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit29.Q ),
    .X(\Inst_LUT4AB_switch_matrix.N4BEG1 ));
 sky130_fd_sc_hd__mux4_1 _1427_ (.A0(net63),
    .A1(net78),
    .A2(net23),
    .A3(net645),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit26.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit27.Q ),
    .X(\Inst_LUT4AB_switch_matrix.N4BEG0 ));
 sky130_fd_sc_hd__mux4_1 _1428_ (.A0(net643),
    .A1(_0653_),
    .A2(\Inst_LUT4AB_switch_matrix.JW2BEG2 ),
    .A3(_0639_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit24.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit25.Q ),
    .X(\Inst_LUT4AB_switch_matrix.N1BEG3 ));
 sky130_fd_sc_hd__mux4_1 _1429_ (.A0(net644),
    .A1(\Inst_LUT4AB_switch_matrix.JW2BEG1 ),
    .A2(net664),
    .A3(_0271_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit23.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit22.Q ),
    .X(\Inst_LUT4AB_switch_matrix.N1BEG2 ));
 sky130_fd_sc_hd__mux4_1 _1430_ (.A0(net637),
    .A1(_0093_),
    .A2(\Inst_LUT4AB_switch_matrix.JW2BEG0 ),
    .A3(_0098_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit20.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit21.Q ),
    .X(\Inst_LUT4AB_switch_matrix.N1BEG1 ));
 sky130_fd_sc_hd__mux4_1 _1431_ (.A0(net650),
    .A1(\Inst_LUT4AB_switch_matrix.JW2BEG3 ),
    .A2(_0192_),
    .A3(_0043_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit19.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit18.Q ),
    .X(\Inst_LUT4AB_switch_matrix.N1BEG0 ));
 sky130_fd_sc_hd__a31o_1 _1432_ (.A1(_0267_),
    .A2(_0294_),
    .A3(_0304_),
    .B1(_0306_),
    .X(net139));
 sky130_fd_sc_hd__mux2_4 _1433_ (.A0(_0280_),
    .A1(_0674_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit29.Q ),
    .X(_0506_));
 sky130_fd_sc_hd__and2b_1 _1434_ (.A_N(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit30.Q ),
    .B(_0506_),
    .X(_0507_));
 sky130_fd_sc_hd__mux2_1 _1435_ (.A0(_0192_),
    .A1(_0139_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit29.Q ),
    .X(_0508_));
 sky130_fd_sc_hd__a211o_1 _1436_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit30.Q ),
    .A2(_0508_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit31.Q ),
    .C1(_0507_),
    .X(_0509_));
 sky130_fd_sc_hd__mux2_1 _1437_ (.A0(\Inst_LUT4AB_switch_matrix.JN2BEG2 ),
    .A1(\Inst_LUT4AB_switch_matrix.E2BEG2 ),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit29.Q ),
    .X(_0510_));
 sky130_fd_sc_hd__mux2_1 _1438_ (.A0(\Inst_LUT4AB_switch_matrix.JS2BEG2 ),
    .A1(\Inst_LUT4AB_switch_matrix.JW2BEG2 ),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit29.Q ),
    .X(_0511_));
 sky130_fd_sc_hd__mux2_1 _1439_ (.A0(_0510_),
    .A1(_0511_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit30.Q ),
    .X(_0512_));
 sky130_fd_sc_hd__o21ai_4 _1440_ (.A1(_0597_),
    .A2(_0512_),
    .B1(_0509_),
    .Y(_0513_));
 sky130_fd_sc_hd__mux2_1 _1441_ (.A0(_0237_),
    .A1(_0629_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q ),
    .X(_0514_));
 sky130_fd_sc_hd__mux2_1 _1442_ (.A0(_0168_),
    .A1(_0093_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q ),
    .X(_0515_));
 sky130_fd_sc_hd__mux2_1 _1443_ (.A0(_0514_),
    .A1(_0515_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit27.Q ),
    .X(_0516_));
 sky130_fd_sc_hd__mux2_1 _1444_ (.A0(\Inst_LUT4AB_switch_matrix.JS2BEG1 ),
    .A1(\Inst_LUT4AB_switch_matrix.JW2BEG1 ),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q ),
    .X(_0517_));
 sky130_fd_sc_hd__mux2_1 _1445_ (.A0(\Inst_LUT4AB_switch_matrix.JN2BEG1 ),
    .A1(\Inst_LUT4AB_switch_matrix.E2BEG1 ),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q ),
    .X(_0518_));
 sky130_fd_sc_hd__inv_1 _1446_ (.A(_0518_),
    .Y(_0519_));
 sky130_fd_sc_hd__o21ai_1 _1447_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit27.Q ),
    .A2(_0519_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit28.Q ),
    .Y(_0520_));
 sky130_fd_sc_hd__a21o_1 _1448_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit27.Q ),
    .A2(_0517_),
    .B1(_0520_),
    .X(_0521_));
 sky130_fd_sc_hd__o21a_4 _1449_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit28.Q ),
    .A2(_0516_),
    .B1(_0521_),
    .X(_0522_));
 sky130_fd_sc_hd__nand2_1 _1450_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit17.Q ),
    .B(_0522_),
    .Y(_0523_));
 sky130_fd_sc_hd__nand2b_1 _1451_ (.A_N(_0323_),
    .B(_0523_),
    .Y(_0524_));
 sky130_fd_sc_hd__o2bb2a_4 _1452_ (.A1_N(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit8.Q ),
    .A2_N(_0513_),
    .B1(_0523_),
    .B2(\Inst_LH_LUT4c_frame_config_dffesr.c_reset_value ),
    .X(_0525_));
 sky130_fd_sc_hd__a32o_1 _1453_ (.A1(net485),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit8.Q ),
    .A3(_0513_),
    .B1(_0524_),
    .B2(_0525_),
    .X(_0000_));
 sky130_fd_sc_hd__nand2_1 _1454_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit11.Q ),
    .B(_0522_),
    .Y(_0526_));
 sky130_fd_sc_hd__nand2_1 _1455_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit2.Q ),
    .B(net467),
    .Y(_0527_));
 sky130_fd_sc_hd__mux2_1 _1456_ (.A0(\Inst_LA_LUT4c_frame_config_dffesr.c_reset_value ),
    .A1(_0696_),
    .S(_0526_),
    .X(_0528_));
 sky130_fd_sc_hd__mux2_1 _1457_ (.A0(net480),
    .A1(_0528_),
    .S(_0527_),
    .X(_0001_));
 sky130_fd_sc_hd__nand2_1 _1458_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit21.Q ),
    .B(_0522_),
    .Y(_0529_));
 sky130_fd_sc_hd__nand2b_1 _1459_ (.A_N(_0035_),
    .B(_0529_),
    .Y(_0530_));
 sky130_fd_sc_hd__o2bb2a_1 _1460_ (.A1_N(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit12.Q ),
    .A2_N(net621),
    .B1(_0529_),
    .B2(\Inst_LB_LUT4c_frame_config_dffesr.c_reset_value ),
    .X(_0531_));
 sky130_fd_sc_hd__a32o_1 _1461_ (.A1(net487),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit12.Q ),
    .A3(net467),
    .B1(_0530_),
    .B2(_0531_),
    .X(_0002_));
 sky130_fd_sc_hd__nand2_1 _1462_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit31.Q ),
    .B(_0522_),
    .Y(_0532_));
 sky130_fd_sc_hd__nand2b_1 _1463_ (.A_N(_0203_),
    .B(_0532_),
    .Y(_0533_));
 sky130_fd_sc_hd__o2bb2a_1 _1464_ (.A1_N(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit22.Q ),
    .A2_N(net621),
    .B1(_0532_),
    .B2(\Inst_LC_LUT4c_frame_config_dffesr.c_reset_value ),
    .X(_0534_));
 sky130_fd_sc_hd__a32o_1 _1465_ (.A1(net486),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit22.Q ),
    .A3(net467),
    .B1(_0533_),
    .B2(_0534_),
    .X(_0003_));
 sky130_fd_sc_hd__nand2_1 _1466_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit9.Q ),
    .B(_0522_),
    .Y(_0535_));
 sky130_fd_sc_hd__nand2b_1 _1467_ (.A_N(_0349_),
    .B(_0535_),
    .Y(_0536_));
 sky130_fd_sc_hd__o2bb2a_1 _1468_ (.A1_N(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit0.Q ),
    .A2_N(net621),
    .B1(_0535_),
    .B2(\Inst_LD_LUT4c_frame_config_dffesr.c_reset_value ),
    .X(_0537_));
 sky130_fd_sc_hd__a32o_1 _1469_ (.A1(net484),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit0.Q ),
    .A3(net467),
    .B1(_0536_),
    .B2(_0537_),
    .X(_0004_));
 sky130_fd_sc_hd__and2_1 _1470_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit10.Q ),
    .B(_0513_),
    .X(_0538_));
 sky130_fd_sc_hd__a21oi_1 _1471_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit19.Q ),
    .A2(_0522_),
    .B1(_0150_),
    .Y(_0539_));
 sky130_fd_sc_hd__a31o_1 _1472_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit19.Q ),
    .A2(_0572_),
    .A3(_0522_),
    .B1(_0538_),
    .X(_0540_));
 sky130_fd_sc_hd__a2bb2o_1 _1473_ (.A1_N(_0539_),
    .A2_N(_0540_),
    .B1(net483),
    .B2(_0538_),
    .X(_0005_));
 sky130_fd_sc_hd__and2_1 _1474_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit20.Q ),
    .B(net621),
    .X(_0541_));
 sky130_fd_sc_hd__a21oi_1 _1475_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit29.Q ),
    .A2(_0522_),
    .B1(_0228_),
    .Y(_0542_));
 sky130_fd_sc_hd__a31o_1 _1476_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit29.Q ),
    .A2(_0573_),
    .A3(_0522_),
    .B1(_0541_),
    .X(_0543_));
 sky130_fd_sc_hd__a2bb2o_1 _1477_ (.A1_N(_0542_),
    .A2_N(_0543_),
    .B1(net482),
    .B2(_0541_),
    .X(_0006_));
 sky130_fd_sc_hd__nand2_1 _1478_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit7.Q ),
    .B(_0522_),
    .Y(_0544_));
 sky130_fd_sc_hd__inv_1 _1479_ (.A(_0544_),
    .Y(_0545_));
 sky130_fd_sc_hd__o2bb2a_1 _1480_ (.A1_N(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit30.Q ),
    .A2_N(net621),
    .B1(_0544_),
    .B2(\Inst_LG_LUT4c_frame_config_dffesr.c_reset_value ),
    .X(_0546_));
 sky130_fd_sc_hd__o31a_1 _1481_ (.A1(_0285_),
    .A2(_0292_),
    .A3(_0545_),
    .B1(_0546_),
    .X(_0547_));
 sky130_fd_sc_hd__a31o_1 _1482_ (.A1(net481),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit30.Q ),
    .A3(net467),
    .B1(_0547_),
    .X(_0007_));
 sky130_fd_sc_hd__dlxtp_1 _1483_ (.D(net779),
    .GATE(net55),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ));
 sky130_fd_sc_hd__dlxtp_1 _1484_ (.D(net777),
    .GATE(net55),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ));
 sky130_fd_sc_hd__dlxtp_1 _1485_ (.D(net774),
    .GATE(net55),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ));
 sky130_fd_sc_hd__dlxtp_1 _1486_ (.D(net771),
    .GATE(net55),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ));
 sky130_fd_sc_hd__dlxtp_1 _1487_ (.D(net769),
    .GATE(net55),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ));
 sky130_fd_sc_hd__dlxtp_1 _1488_ (.D(net767),
    .GATE(net55),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ));
 sky130_fd_sc_hd__dlxtp_1 _1489_ (.D(net763),
    .GATE(net55),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ));
 sky130_fd_sc_hd__dlxtp_1 _1490_ (.D(net761),
    .GATE(net55),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ));
 sky130_fd_sc_hd__dlxtp_1 _1491_ (.D(net811),
    .GATE(net704),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ));
 sky130_fd_sc_hd__dlxtp_1 _1492_ (.D(net789),
    .GATE(net704),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ));
 sky130_fd_sc_hd__dlxtp_1 _1493_ (.D(net766),
    .GATE(net704),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ));
 sky130_fd_sc_hd__dlxtp_1 _1494_ (.D(net760),
    .GATE(net706),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ));
 sky130_fd_sc_hd__dlxtp_1 _1495_ (.D(net757),
    .GATE(net703),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ));
 sky130_fd_sc_hd__dlxtp_1 _1496_ (.D(net755),
    .GATE(net703),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ));
 sky130_fd_sc_hd__dlxtp_1 _1497_ (.D(net753),
    .GATE(net704),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ));
 sky130_fd_sc_hd__dlxtp_1 _1498_ (.D(net751),
    .GATE(net704),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ));
 sky130_fd_sc_hd__dlxtp_1 _1499_ (.D(net749),
    .GATE(net704),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.c_out_mux ));
 sky130_fd_sc_hd__dlxtp_1 _1500_ (.D(net747),
    .GATE(net705),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.c_I0mux ));
 sky130_fd_sc_hd__dlxtp_1 _1501_ (.D(net809),
    .GATE(net703),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.c_reset_value ));
 sky130_fd_sc_hd__dlxtp_1 _1502_ (.D(net807),
    .GATE(net703),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ));
 sky130_fd_sc_hd__dlxtp_1 _1503_ (.D(net806),
    .GATE(net703),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ));
 sky130_fd_sc_hd__dlxtp_1 _1504_ (.D(net804),
    .GATE(net705),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ));
 sky130_fd_sc_hd__dlxtp_1 _1505_ (.D(net801),
    .GATE(net705),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ));
 sky130_fd_sc_hd__dlxtp_1 _1506_ (.D(net799),
    .GATE(net705),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ));
 sky130_fd_sc_hd__dlxtp_1 _1507_ (.D(net798),
    .GATE(net703),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ));
 sky130_fd_sc_hd__dlxtp_1 _1508_ (.D(net796),
    .GATE(net703),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ));
 sky130_fd_sc_hd__dlxtp_1 _1509_ (.D(net793),
    .GATE(net705),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ));
 sky130_fd_sc_hd__dlxtp_1 _1510_ (.D(net791),
    .GATE(net705),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ));
 sky130_fd_sc_hd__dlxtp_1 _1511_ (.D(net787),
    .GATE(net704),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ));
 sky130_fd_sc_hd__dlxtp_1 _1512_ (.D(net785),
    .GATE(net705),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ));
 sky130_fd_sc_hd__dlxtp_1 _1513_ (.D(net784),
    .GATE(net705),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ));
 sky130_fd_sc_hd__dlxtp_1 _1514_ (.D(net782),
    .GATE(net705),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ));
 sky130_fd_sc_hd__dlxtp_1 _1515_ (.D(net779),
    .GATE(net703),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ));
 sky130_fd_sc_hd__dlxtp_1 _1516_ (.D(net777),
    .GATE(net703),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ));
 sky130_fd_sc_hd__dlxtp_1 _1517_ (.D(net774),
    .GATE(net703),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ));
 sky130_fd_sc_hd__dlxtp_1 _1518_ (.D(net771),
    .GATE(net704),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.c_out_mux ));
 sky130_fd_sc_hd__dlxtp_1 _1519_ (.D(net769),
    .GATE(net705),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.c_I0mux ));
 sky130_fd_sc_hd__dlxtp_1 _1520_ (.D(net767),
    .GATE(net704),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.c_reset_value ));
 sky130_fd_sc_hd__dlxtp_1 _1521_ (.D(net763),
    .GATE(net706),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ));
 sky130_fd_sc_hd__dlxtp_1 _1522_ (.D(net761),
    .GATE(net706),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ));
 sky130_fd_sc_hd__dlxtp_1 _1523_ (.D(net811),
    .GATE(net708),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ));
 sky130_fd_sc_hd__dlxtp_1 _1524_ (.D(net789),
    .GATE(net707),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ));
 sky130_fd_sc_hd__dlxtp_1 _1525_ (.D(net766),
    .GATE(net708),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ));
 sky130_fd_sc_hd__dlxtp_1 _1526_ (.D(net760),
    .GATE(net707),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ));
 sky130_fd_sc_hd__dlxtp_1 _1527_ (.D(net757),
    .GATE(net707),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ));
 sky130_fd_sc_hd__dlxtp_1 _1528_ (.D(net755),
    .GATE(net707),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ));
 sky130_fd_sc_hd__dlxtp_1 _1529_ (.D(net753),
    .GATE(net707),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ));
 sky130_fd_sc_hd__dlxtp_1 _1530_ (.D(net751),
    .GATE(net707),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ));
 sky130_fd_sc_hd__dlxtp_1 _1531_ (.D(net749),
    .GATE(net707),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ));
 sky130_fd_sc_hd__dlxtp_1 _1532_ (.D(net747),
    .GATE(net708),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ));
 sky130_fd_sc_hd__dlxtp_1 _1533_ (.D(net809),
    .GATE(net707),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ));
 sky130_fd_sc_hd__dlxtp_1 _1534_ (.D(net807),
    .GATE(net708),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ));
 sky130_fd_sc_hd__dlxtp_1 _1535_ (.D(net806),
    .GATE(net707),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ));
 sky130_fd_sc_hd__dlxtp_1 _1536_ (.D(net804),
    .GATE(net707),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ));
 sky130_fd_sc_hd__dlxtp_1 _1537_ (.D(net801),
    .GATE(net711),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.c_out_mux ));
 sky130_fd_sc_hd__dlxtp_1 _1538_ (.D(net799),
    .GATE(net708),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.c_I0mux ));
 sky130_fd_sc_hd__dlxtp_1 _1539_ (.D(net798),
    .GATE(net711),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.c_reset_value ));
 sky130_fd_sc_hd__dlxtp_1 _1540_ (.D(net796),
    .GATE(net709),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ));
 sky130_fd_sc_hd__dlxtp_1 _1541_ (.D(net793),
    .GATE(net709),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ));
 sky130_fd_sc_hd__dlxtp_1 _1542_ (.D(net791),
    .GATE(net709),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ));
 sky130_fd_sc_hd__dlxtp_1 _1543_ (.D(net787),
    .GATE(net709),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ));
 sky130_fd_sc_hd__dlxtp_1 _1544_ (.D(net785),
    .GATE(net709),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ));
 sky130_fd_sc_hd__dlxtp_1 _1545_ (.D(net784),
    .GATE(net709),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ));
 sky130_fd_sc_hd__dlxtp_1 _1546_ (.D(net782),
    .GATE(net709),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ));
 sky130_fd_sc_hd__dlxtp_1 _1547_ (.D(net779),
    .GATE(net709),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ));
 sky130_fd_sc_hd__dlxtp_1 _1548_ (.D(net777),
    .GATE(net709),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ));
 sky130_fd_sc_hd__dlxtp_1 _1549_ (.D(net775),
    .GATE(net710),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ));
 sky130_fd_sc_hd__dlxtp_1 _1550_ (.D(net772),
    .GATE(net710),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ));
 sky130_fd_sc_hd__dlxtp_1 _1551_ (.D(net44),
    .GATE(net710),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ));
 sky130_fd_sc_hd__dlxtp_1 _1552_ (.D(net768),
    .GATE(net710),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ));
 sky130_fd_sc_hd__dlxtp_1 _1553_ (.D(net46),
    .GATE(net710),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ));
 sky130_fd_sc_hd__dlxtp_1 _1554_ (.D(net762),
    .GATE(net710),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ));
 sky130_fd_sc_hd__dlxtp_1 _1555_ (.D(net811),
    .GATE(net715),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ));
 sky130_fd_sc_hd__dlxtp_1 _1556_ (.D(net789),
    .GATE(net715),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.c_out_mux ));
 sky130_fd_sc_hd__dlxtp_1 _1557_ (.D(net765),
    .GATE(net715),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.c_I0mux ));
 sky130_fd_sc_hd__dlxtp_1 _1558_ (.D(net760),
    .GATE(net715),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.c_reset_value ));
 sky130_fd_sc_hd__dlxtp_1 _1559_ (.D(net758),
    .GATE(net712),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ));
 sky130_fd_sc_hd__dlxtp_1 _1560_ (.D(net756),
    .GATE(net712),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ));
 sky130_fd_sc_hd__dlxtp_1 _1561_ (.D(net753),
    .GATE(net713),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ));
 sky130_fd_sc_hd__dlxtp_1 _1562_ (.D(net751),
    .GATE(net713),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ));
 sky130_fd_sc_hd__dlxtp_1 _1563_ (.D(net749),
    .GATE(net713),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ));
 sky130_fd_sc_hd__dlxtp_1 _1564_ (.D(net747),
    .GATE(net713),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ));
 sky130_fd_sc_hd__dlxtp_1 _1565_ (.D(net809),
    .GATE(net712),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ));
 sky130_fd_sc_hd__dlxtp_1 _1566_ (.D(net807),
    .GATE(net712),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ));
 sky130_fd_sc_hd__dlxtp_1 _1567_ (.D(net806),
    .GATE(net712),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ));
 sky130_fd_sc_hd__dlxtp_1 _1568_ (.D(net804),
    .GATE(net712),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ));
 sky130_fd_sc_hd__dlxtp_1 _1569_ (.D(net801),
    .GATE(net713),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ));
 sky130_fd_sc_hd__dlxtp_1 _1570_ (.D(net799),
    .GATE(net712),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ));
 sky130_fd_sc_hd__dlxtp_1 _1571_ (.D(net798),
    .GATE(net713),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ));
 sky130_fd_sc_hd__dlxtp_1 _1572_ (.D(net796),
    .GATE(net712),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ));
 sky130_fd_sc_hd__dlxtp_1 _1573_ (.D(net793),
    .GATE(net712),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ));
 sky130_fd_sc_hd__dlxtp_1 _1574_ (.D(net791),
    .GATE(net712),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ));
 sky130_fd_sc_hd__dlxtp_1 _1575_ (.D(net787),
    .GATE(net714),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.c_out_mux ));
 sky130_fd_sc_hd__dlxtp_1 _1576_ (.D(net785),
    .GATE(net714),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.c_I0mux ));
 sky130_fd_sc_hd__dlxtp_1 _1577_ (.D(net784),
    .GATE(net714),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.c_reset_value ));
 sky130_fd_sc_hd__dlxtp_1 _1578_ (.D(net782),
    .GATE(net716),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ));
 sky130_fd_sc_hd__dlxtp_1 _1579_ (.D(net779),
    .GATE(net716),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ));
 sky130_fd_sc_hd__dlxtp_1 _1580_ (.D(net777),
    .GATE(net716),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ));
 sky130_fd_sc_hd__dlxtp_1 _1581_ (.D(net775),
    .GATE(net716),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ));
 sky130_fd_sc_hd__dlxtp_1 _1582_ (.D(net771),
    .GATE(net716),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ));
 sky130_fd_sc_hd__dlxtp_1 _1583_ (.D(net769),
    .GATE(net716),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ));
 sky130_fd_sc_hd__dlxtp_1 _1584_ (.D(net45),
    .GATE(net716),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ));
 sky130_fd_sc_hd__dlxtp_1 _1585_ (.D(net764),
    .GATE(net716),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ));
 sky130_fd_sc_hd__dlxtp_1 _1586_ (.D(net762),
    .GATE(net716),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ));
 sky130_fd_sc_hd__dlxtp_1 _1587_ (.D(net811),
    .GATE(net720),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ));
 sky130_fd_sc_hd__dlxtp_1 _1588_ (.D(net39),
    .GATE(net720),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ));
 sky130_fd_sc_hd__dlxtp_1 _1589_ (.D(net766),
    .GATE(net717),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ));
 sky130_fd_sc_hd__dlxtp_1 _1590_ (.D(net760),
    .GATE(net717),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ));
 sky130_fd_sc_hd__dlxtp_1 _1591_ (.D(net758),
    .GATE(net717),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ));
 sky130_fd_sc_hd__dlxtp_1 _1592_ (.D(net756),
    .GATE(net717),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ));
 sky130_fd_sc_hd__dlxtp_1 _1593_ (.D(net753),
    .GATE(net717),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ));
 sky130_fd_sc_hd__dlxtp_1 _1594_ (.D(net751),
    .GATE(net717),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.c_out_mux ));
 sky130_fd_sc_hd__dlxtp_1 _1595_ (.D(net749),
    .GATE(net717),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.c_I0mux ));
 sky130_fd_sc_hd__dlxtp_1 _1596_ (.D(net747),
    .GATE(net717),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.c_reset_value ));
 sky130_fd_sc_hd__dlxtp_1 _1597_ (.D(net809),
    .GATE(net718),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ));
 sky130_fd_sc_hd__dlxtp_1 _1598_ (.D(net807),
    .GATE(net717),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ));
 sky130_fd_sc_hd__dlxtp_1 _1599_ (.D(net31),
    .GATE(net718),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ));
 sky130_fd_sc_hd__dlxtp_1 _1600_ (.D(net32),
    .GATE(net719),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ));
 sky130_fd_sc_hd__dlxtp_1 _1601_ (.D(net801),
    .GATE(net718),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ));
 sky130_fd_sc_hd__dlxtp_1 _1602_ (.D(net799),
    .GATE(net719),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ));
 sky130_fd_sc_hd__dlxtp_1 _1603_ (.D(net798),
    .GATE(net718),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ));
 sky130_fd_sc_hd__dlxtp_1 _1604_ (.D(net796),
    .GATE(net717),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ));
 sky130_fd_sc_hd__dlxtp_1 _1605_ (.D(net793),
    .GATE(net718),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ));
 sky130_fd_sc_hd__dlxtp_1 _1606_ (.D(net791),
    .GATE(net719),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ));
 sky130_fd_sc_hd__dlxtp_1 _1607_ (.D(net787),
    .GATE(net718),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ));
 sky130_fd_sc_hd__dlxtp_1 _1608_ (.D(net785),
    .GATE(net718),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ));
 sky130_fd_sc_hd__dlxtp_1 _1609_ (.D(net784),
    .GATE(net718),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ));
 sky130_fd_sc_hd__dlxtp_1 _1610_ (.D(net782),
    .GATE(net718),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ));
 sky130_fd_sc_hd__dlxtp_1 _1611_ (.D(net779),
    .GATE(net718),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ));
 sky130_fd_sc_hd__dlxtp_1 _1612_ (.D(net777),
    .GATE(net720),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ));
 sky130_fd_sc_hd__dlxtp_1 _1613_ (.D(net775),
    .GATE(net719),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.c_out_mux ));
 sky130_fd_sc_hd__dlxtp_1 _1614_ (.D(net772),
    .GATE(net720),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.c_I0mux ));
 sky130_fd_sc_hd__dlxtp_1 _1615_ (.D(net44),
    .GATE(net719),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.c_reset_value ));
 sky130_fd_sc_hd__dlxtp_1 _1616_ (.D(net767),
    .GATE(net719),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ));
 sky130_fd_sc_hd__dlxtp_1 _1617_ (.D(net764),
    .GATE(net719),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ));
 sky130_fd_sc_hd__dlxtp_1 _1618_ (.D(net762),
    .GATE(net719),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ));
 sky130_fd_sc_hd__dlxtp_1 _1619_ (.D(net811),
    .GATE(net723),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ));
 sky130_fd_sc_hd__dlxtp_1 _1620_ (.D(net789),
    .GATE(net723),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ));
 sky130_fd_sc_hd__dlxtp_1 _1621_ (.D(net765),
    .GATE(net723),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ));
 sky130_fd_sc_hd__dlxtp_1 _1622_ (.D(net760),
    .GATE(net723),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ));
 sky130_fd_sc_hd__dlxtp_1 _1623_ (.D(net758),
    .GATE(net723),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ));
 sky130_fd_sc_hd__dlxtp_1 _1624_ (.D(net756),
    .GATE(net723),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ));
 sky130_fd_sc_hd__dlxtp_1 _1625_ (.D(net753),
    .GATE(net723),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ));
 sky130_fd_sc_hd__dlxtp_1 _1626_ (.D(net751),
    .GATE(net723),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ));
 sky130_fd_sc_hd__dlxtp_1 _1627_ (.D(net749),
    .GATE(net724),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ));
 sky130_fd_sc_hd__dlxtp_1 _1628_ (.D(net747),
    .GATE(net724),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ));
 sky130_fd_sc_hd__dlxtp_1 _1629_ (.D(net809),
    .GATE(net724),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ));
 sky130_fd_sc_hd__dlxtp_1 _1630_ (.D(net807),
    .GATE(net723),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ));
 sky130_fd_sc_hd__dlxtp_1 _1631_ (.D(net805),
    .GATE(net723),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ));
 sky130_fd_sc_hd__dlxtp_1 _1632_ (.D(net803),
    .GATE(net725),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.c_out_mux ));
 sky130_fd_sc_hd__dlxtp_1 _1633_ (.D(net801),
    .GATE(net724),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.c_I0mux ));
 sky130_fd_sc_hd__dlxtp_1 _1634_ (.D(net799),
    .GATE(net724),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.c_reset_value ));
 sky130_fd_sc_hd__dlxtp_1 _1635_ (.D(net797),
    .GATE(net722),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1636_ (.D(net795),
    .GATE(net722),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1637_ (.D(net794),
    .GATE(net721),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1638_ (.D(net792),
    .GATE(net721),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1639_ (.D(net788),
    .GATE(net721),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1640_ (.D(net786),
    .GATE(net721),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1641_ (.D(net783),
    .GATE(net721),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1642_ (.D(net781),
    .GATE(net721),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1643_ (.D(net780),
    .GATE(net721),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1644_ (.D(net778),
    .GATE(net721),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1645_ (.D(net776),
    .GATE(net721),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1646_ (.D(net773),
    .GATE(net721),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1647_ (.D(net770),
    .GATE(net722),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1648_ (.D(net768),
    .GATE(net722),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1649_ (.D(net764),
    .GATE(net722),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1650_ (.D(net47),
    .GATE(net722),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1651_ (.D(net812),
    .GATE(net728),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1652_ (.D(net790),
    .GATE(net728),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1653_ (.D(net765),
    .GATE(net727),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1654_ (.D(net759),
    .GATE(net726),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1655_ (.D(net758),
    .GATE(net727),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1656_ (.D(net756),
    .GATE(net726),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1657_ (.D(net754),
    .GATE(net726),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1658_ (.D(net752),
    .GATE(net726),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1659_ (.D(net750),
    .GATE(net727),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1660_ (.D(net748),
    .GATE(net726),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1661_ (.D(net810),
    .GATE(net727),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1662_ (.D(net808),
    .GATE(net726),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1663_ (.D(net805),
    .GATE(net726),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1664_ (.D(net803),
    .GATE(net726),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1665_ (.D(net801),
    .GATE(net728),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1666_ (.D(net799),
    .GATE(net728),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1667_ (.D(net797),
    .GATE(net728),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1668_ (.D(net795),
    .GATE(net728),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1669_ (.D(net793),
    .GATE(net728),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1670_ (.D(net791),
    .GATE(net728),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1671_ (.D(net787),
    .GATE(net728),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1672_ (.D(net785),
    .GATE(net728),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1673_ (.D(net784),
    .GATE(net727),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1674_ (.D(net782),
    .GATE(net727),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1675_ (.D(net779),
    .GATE(net727),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1676_ (.D(net43),
    .GATE(net726),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1677_ (.D(net775),
    .GATE(net726),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1678_ (.D(net772),
    .GATE(net727),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1679_ (.D(net769),
    .GATE(net729),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1680_ (.D(net767),
    .GATE(net729),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1681_ (.D(net764),
    .GATE(net729),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1682_ (.D(net762),
    .GATE(net729),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1683_ (.D(net28),
    .GATE(net734),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1684_ (.D(net789),
    .GATE(net733),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1685_ (.D(net765),
    .GATE(net733),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1686_ (.D(net760),
    .GATE(net733),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1687_ (.D(net758),
    .GATE(net733),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1688_ (.D(net756),
    .GATE(net733),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1689_ (.D(net50),
    .GATE(net733),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1690_ (.D(net51),
    .GATE(net733),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1691_ (.D(net52),
    .GATE(net733),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1692_ (.D(net53),
    .GATE(net733),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1693_ (.D(net810),
    .GATE(net732),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1694_ (.D(net808),
    .GATE(net732),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1695_ (.D(net806),
    .GATE(net730),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1696_ (.D(net804),
    .GATE(net730),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1697_ (.D(net802),
    .GATE(net730),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1698_ (.D(net800),
    .GATE(net730),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1699_ (.D(net797),
    .GATE(net730),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1700_ (.D(net795),
    .GATE(net730),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1701_ (.D(net794),
    .GATE(net730),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1702_ (.D(net792),
    .GATE(net730),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1703_ (.D(net787),
    .GATE(net730),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1704_ (.D(net785),
    .GATE(net730),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1705_ (.D(net784),
    .GATE(net732),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1706_ (.D(net782),
    .GATE(net732),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1707_ (.D(net779),
    .GATE(net731),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1708_ (.D(net777),
    .GATE(net731),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1709_ (.D(net774),
    .GATE(net734),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1710_ (.D(net771),
    .GATE(net731),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1711_ (.D(net769),
    .GATE(net734),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1712_ (.D(net767),
    .GATE(net731),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1713_ (.D(net763),
    .GATE(net731),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1714_ (.D(net762),
    .GATE(net731),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1715_ (.D(net811),
    .GATE(net738),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1716_ (.D(net789),
    .GATE(net738),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1717_ (.D(net766),
    .GATE(net738),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1718_ (.D(net48),
    .GATE(net738),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1719_ (.D(net757),
    .GATE(net738),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1720_ (.D(net755),
    .GATE(net738),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1721_ (.D(net754),
    .GATE(net737),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1722_ (.D(net752),
    .GATE(net737),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1723_ (.D(net750),
    .GATE(net737),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1724_ (.D(net748),
    .GATE(net737),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1725_ (.D(net810),
    .GATE(net737),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1726_ (.D(net808),
    .GATE(net737),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1727_ (.D(net806),
    .GATE(net738),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1728_ (.D(net804),
    .GATE(net738),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1729_ (.D(net802),
    .GATE(net737),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1730_ (.D(net800),
    .GATE(net737),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1731_ (.D(net798),
    .GATE(net737),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1732_ (.D(net795),
    .GATE(net736),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1733_ (.D(net794),
    .GATE(net736),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1734_ (.D(net792),
    .GATE(net736),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1735_ (.D(net788),
    .GATE(net735),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1736_ (.D(net786),
    .GATE(net735),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1737_ (.D(net783),
    .GATE(net735),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1738_ (.D(net781),
    .GATE(net736),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1739_ (.D(net780),
    .GATE(net735),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1740_ (.D(net778),
    .GATE(net736),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1741_ (.D(net776),
    .GATE(net735),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1742_ (.D(net773),
    .GATE(net735),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1743_ (.D(net770),
    .GATE(net735),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1744_ (.D(net768),
    .GATE(net735),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1745_ (.D(net764),
    .GATE(net735),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1746_ (.D(net47),
    .GATE(net735),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1747_ (.D(net812),
    .GATE(net54),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1748_ (.D(net790),
    .GATE(net54),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1749_ (.D(net766),
    .GATE(net739),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1750_ (.D(net760),
    .GATE(net742),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1751_ (.D(net757),
    .GATE(net740),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1752_ (.D(net755),
    .GATE(net740),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1753_ (.D(net753),
    .GATE(net740),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1754_ (.D(net751),
    .GATE(net741),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1755_ (.D(net749),
    .GATE(net741),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1756_ (.D(net747),
    .GATE(net739),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1757_ (.D(net809),
    .GATE(net739),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1758_ (.D(net807),
    .GATE(net739),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1759_ (.D(net806),
    .GATE(net739),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1760_ (.D(net804),
    .GATE(net742),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1761_ (.D(net801),
    .GATE(net742),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1762_ (.D(net799),
    .GATE(net740),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1763_ (.D(net798),
    .GATE(net741),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1764_ (.D(net796),
    .GATE(net741),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1765_ (.D(net793),
    .GATE(net741),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1766_ (.D(net791),
    .GATE(net740),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1767_ (.D(net787),
    .GATE(net740),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1768_ (.D(net785),
    .GATE(net739),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1769_ (.D(net784),
    .GATE(net739),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1770_ (.D(net782),
    .GATE(net742),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1771_ (.D(net779),
    .GATE(net742),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1772_ (.D(net777),
    .GATE(net742),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1773_ (.D(net774),
    .GATE(net742),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1774_ (.D(net771),
    .GATE(net54),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1775_ (.D(net769),
    .GATE(net742),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1776_ (.D(net767),
    .GATE(net739),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1777_ (.D(net764),
    .GATE(net739),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1778_ (.D(net761),
    .GATE(net739),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1779_ (.D(net811),
    .GATE(net670),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1780_ (.D(net789),
    .GATE(net670),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1781_ (.D(net765),
    .GATE(net670),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1782_ (.D(net759),
    .GATE(net670),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1783_ (.D(net757),
    .GATE(net670),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1784_ (.D(net756),
    .GATE(net670),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1785_ (.D(net753),
    .GATE(net670),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1786_ (.D(net751),
    .GATE(net670),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1787_ (.D(net749),
    .GATE(net670),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1788_ (.D(net747),
    .GATE(net669),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1789_ (.D(net809),
    .GATE(net668),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1790_ (.D(net807),
    .GATE(net667),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1791_ (.D(net805),
    .GATE(net667),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1792_ (.D(net803),
    .GATE(net668),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1793_ (.D(net801),
    .GATE(net668),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1794_ (.D(net799),
    .GATE(net668),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1795_ (.D(net35),
    .GATE(net669),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1796_ (.D(net36),
    .GATE(net667),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1797_ (.D(net793),
    .GATE(net667),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1798_ (.D(net791),
    .GATE(net668),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1799_ (.D(net787),
    .GATE(net668),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1800_ (.D(net785),
    .GATE(net667),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1801_ (.D(net784),
    .GATE(net667),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1802_ (.D(net782),
    .GATE(net667),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1803_ (.D(net42),
    .GATE(net667),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1804_ (.D(net777),
    .GATE(net668),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1805_ (.D(net774),
    .GATE(net668),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1806_ (.D(net772),
    .GATE(net667),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1807_ (.D(net770),
    .GATE(net667),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1808_ (.D(net45),
    .GATE(net668),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1809_ (.D(net764),
    .GATE(net669),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1810_ (.D(net762),
    .GATE(net669),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1811_ (.D(net811),
    .GATE(net671),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1812_ (.D(net789),
    .GATE(net671),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1813_ (.D(net765),
    .GATE(net671),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1814_ (.D(net760),
    .GATE(net672),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1815_ (.D(net758),
    .GATE(net672),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1816_ (.D(net755),
    .GATE(net674),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1817_ (.D(net753),
    .GATE(net674),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1818_ (.D(net751),
    .GATE(net671),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1819_ (.D(net749),
    .GATE(net671),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1820_ (.D(net747),
    .GATE(net671),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1821_ (.D(net809),
    .GATE(net671),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1822_ (.D(net807),
    .GATE(net671),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1823_ (.D(net806),
    .GATE(net671),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1824_ (.D(net804),
    .GATE(net672),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1825_ (.D(net801),
    .GATE(net672),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1826_ (.D(net799),
    .GATE(net674),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1827_ (.D(net798),
    .GATE(net674),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1828_ (.D(net796),
    .GATE(net672),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1829_ (.D(net794),
    .GATE(net673),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1830_ (.D(net792),
    .GATE(net673),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1831_ (.D(net788),
    .GATE(net673),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1832_ (.D(net786),
    .GATE(net673),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1833_ (.D(net783),
    .GATE(net673),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1834_ (.D(net781),
    .GATE(net673),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1835_ (.D(net780),
    .GATE(net673),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1836_ (.D(net778),
    .GATE(net673),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1837_ (.D(net774),
    .GATE(net674),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1838_ (.D(net771),
    .GATE(net674),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1839_ (.D(net769),
    .GATE(net674),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1840_ (.D(net767),
    .GATE(net674),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1841_ (.D(net763),
    .GATE(net674),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1842_ (.D(net761),
    .GATE(net674),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1843_ (.D(net812),
    .GATE(net675),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1844_ (.D(net790),
    .GATE(net675),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1845_ (.D(net765),
    .GATE(net676),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1846_ (.D(net759),
    .GATE(net676),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1847_ (.D(net758),
    .GATE(net678),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1848_ (.D(net49),
    .GATE(net678),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1849_ (.D(net754),
    .GATE(net677),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1850_ (.D(net752),
    .GATE(net677),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1851_ (.D(net750),
    .GATE(net675),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1852_ (.D(net748),
    .GATE(net675),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1853_ (.D(net810),
    .GATE(net677),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1854_ (.D(net808),
    .GATE(net677),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1855_ (.D(net805),
    .GATE(net676),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1856_ (.D(net803),
    .GATE(net676),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1857_ (.D(net802),
    .GATE(net677),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1858_ (.D(net800),
    .GATE(net677),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1859_ (.D(net797),
    .GATE(net675),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1860_ (.D(net795),
    .GATE(net675),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1861_ (.D(net793),
    .GATE(net677),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1862_ (.D(net791),
    .GATE(net676),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1863_ (.D(net787),
    .GATE(net676),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1864_ (.D(net785),
    .GATE(net676),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1865_ (.D(net783),
    .GATE(net677),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1866_ (.D(net781),
    .GATE(net677),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1867_ (.D(net780),
    .GATE(net675),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1868_ (.D(net778),
    .GATE(net675),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1869_ (.D(net774),
    .GATE(net678),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1870_ (.D(net771),
    .GATE(net678),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1871_ (.D(net770),
    .GATE(net675),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1872_ (.D(net768),
    .GATE(net675),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1873_ (.D(net46),
    .GATE(net676),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1874_ (.D(net762),
    .GATE(net676),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1875_ (.D(net811),
    .GATE(net680),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1876_ (.D(net789),
    .GATE(net680),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1877_ (.D(net766),
    .GATE(net681),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1878_ (.D(net759),
    .GATE(net681),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1879_ (.D(net757),
    .GATE(net679),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1880_ (.D(net755),
    .GATE(net679),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1881_ (.D(net753),
    .GATE(net681),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1882_ (.D(net751),
    .GATE(net681),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1883_ (.D(net750),
    .GATE(net679),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1884_ (.D(net748),
    .GATE(net679),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1885_ (.D(net809),
    .GATE(net682),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1886_ (.D(net807),
    .GATE(net682),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1887_ (.D(net806),
    .GATE(net679),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1888_ (.D(net804),
    .GATE(net679),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1889_ (.D(net33),
    .GATE(net681),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1890_ (.D(net34),
    .GATE(net681),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1891_ (.D(net798),
    .GATE(net680),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1892_ (.D(net796),
    .GATE(net680),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1893_ (.D(net793),
    .GATE(net681),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1894_ (.D(net791),
    .GATE(net681),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1895_ (.D(net788),
    .GATE(net679),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1896_ (.D(net786),
    .GATE(net679),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1897_ (.D(net784),
    .GATE(net682),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1898_ (.D(net782),
    .GATE(net681),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1899_ (.D(net779),
    .GATE(net680),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1900_ (.D(net777),
    .GATE(net680),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1901_ (.D(net774),
    .GATE(net682),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1902_ (.D(net772),
    .GATE(net682),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1903_ (.D(net770),
    .GATE(net679),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1904_ (.D(net768),
    .GATE(net679),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1905_ (.D(net763),
    .GATE(net682),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1906_ (.D(net761),
    .GATE(net682),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1907_ (.D(net812),
    .GATE(net684),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1908_ (.D(net790),
    .GATE(net684),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1909_ (.D(net765),
    .GATE(net686),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1910_ (.D(net759),
    .GATE(net686),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1911_ (.D(net757),
    .GATE(net684),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1912_ (.D(net755),
    .GATE(net684),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1913_ (.D(net754),
    .GATE(net684),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1914_ (.D(net752),
    .GATE(net684),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1915_ (.D(net750),
    .GATE(net683),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1916_ (.D(net748),
    .GATE(net683),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1917_ (.D(net810),
    .GATE(net685),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1918_ (.D(net808),
    .GATE(net686),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1919_ (.D(net805),
    .GATE(net685),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1920_ (.D(net803),
    .GATE(net685),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1921_ (.D(net802),
    .GATE(net685),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1922_ (.D(net800),
    .GATE(net685),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1923_ (.D(net797),
    .GATE(net683),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1924_ (.D(net795),
    .GATE(net683),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1925_ (.D(net794),
    .GATE(net685),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1926_ (.D(net792),
    .GATE(net685),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1927_ (.D(net40),
    .GATE(net686),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1928_ (.D(net41),
    .GATE(net686),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1929_ (.D(net783),
    .GATE(net685),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1930_ (.D(net781),
    .GATE(net685),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1931_ (.D(net780),
    .GATE(net683),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1932_ (.D(net778),
    .GATE(net683),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1933_ (.D(net776),
    .GATE(net683),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1934_ (.D(net773),
    .GATE(net683),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1935_ (.D(net770),
    .GATE(net684),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1936_ (.D(net768),
    .GATE(net684),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1937_ (.D(net763),
    .GATE(net683),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1938_ (.D(net761),
    .GATE(net683),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1939_ (.D(net812),
    .GATE(net687),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1940_ (.D(net790),
    .GATE(net687),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1941_ (.D(net765),
    .GATE(net690),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1942_ (.D(net759),
    .GATE(net690),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1943_ (.D(net758),
    .GATE(net690),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1944_ (.D(net756),
    .GATE(net690),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1945_ (.D(net754),
    .GATE(net56),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1946_ (.D(net752),
    .GATE(net56),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1947_ (.D(net750),
    .GATE(net687),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1948_ (.D(net748),
    .GATE(net687),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1949_ (.D(net810),
    .GATE(net688),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1950_ (.D(net808),
    .GATE(net688),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1951_ (.D(net805),
    .GATE(net688),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1952_ (.D(net803),
    .GATE(net688),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1953_ (.D(net802),
    .GATE(net688),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1954_ (.D(net800),
    .GATE(net688),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1955_ (.D(net797),
    .GATE(net688),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1956_ (.D(net795),
    .GATE(net688),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1957_ (.D(net794),
    .GATE(net688),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1958_ (.D(net792),
    .GATE(net688),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1959_ (.D(net788),
    .GATE(net689),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1960_ (.D(net786),
    .GATE(net689),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1961_ (.D(net783),
    .GATE(net689),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1962_ (.D(net781),
    .GATE(net689),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1963_ (.D(net780),
    .GATE(net689),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1964_ (.D(net778),
    .GATE(net689),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1965_ (.D(net776),
    .GATE(net687),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1966_ (.D(net773),
    .GATE(net687),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1967_ (.D(net770),
    .GATE(net687),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1968_ (.D(net768),
    .GATE(net687),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1969_ (.D(net763),
    .GATE(net687),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1970_ (.D(net761),
    .GATE(net687),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1971_ (.D(net812),
    .GATE(net694),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1972_ (.D(net790),
    .GATE(net694),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1973_ (.D(net765),
    .GATE(net694),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1974_ (.D(net759),
    .GATE(net694),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1975_ (.D(net758),
    .GATE(net693),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1976_ (.D(net756),
    .GATE(net693),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1977_ (.D(net754),
    .GATE(net691),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1978_ (.D(net752),
    .GATE(net691),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1979_ (.D(net750),
    .GATE(net691),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1980_ (.D(net748),
    .GATE(net691),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1981_ (.D(net810),
    .GATE(net693),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1982_ (.D(net808),
    .GATE(net692),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1983_ (.D(net805),
    .GATE(net692),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1984_ (.D(net803),
    .GATE(net692),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1985_ (.D(net802),
    .GATE(net692),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1986_ (.D(net800),
    .GATE(net692),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1987_ (.D(net797),
    .GATE(net692),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1988_ (.D(net795),
    .GATE(net692),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1989_ (.D(net794),
    .GATE(net692),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1990_ (.D(net792),
    .GATE(net692),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1991_ (.D(net788),
    .GATE(net692),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1992_ (.D(net786),
    .GATE(net693),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1993_ (.D(net783),
    .GATE(net693),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1994_ (.D(net781),
    .GATE(net693),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1995_ (.D(net42),
    .GATE(net693),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1996_ (.D(net43),
    .GATE(net693),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1997_ (.D(net776),
    .GATE(net691),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1998_ (.D(net773),
    .GATE(net691),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1999_ (.D(net770),
    .GATE(net691),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2000_ (.D(net768),
    .GATE(net691),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2001_ (.D(net763),
    .GATE(net691),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2002_ (.D(net761),
    .GATE(net691),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2003_ (.D(net812),
    .GATE(net695),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2004_ (.D(net790),
    .GATE(net695),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2005_ (.D(net766),
    .GATE(net696),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2006_ (.D(net759),
    .GATE(net696),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2007_ (.D(net757),
    .GATE(net696),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2008_ (.D(net755),
    .GATE(net696),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2009_ (.D(net754),
    .GATE(net696),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2010_ (.D(net752),
    .GATE(net696),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2011_ (.D(net750),
    .GATE(net695),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2012_ (.D(net748),
    .GATE(net695),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2013_ (.D(net810),
    .GATE(net698),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2014_ (.D(net808),
    .GATE(net698),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2015_ (.D(net805),
    .GATE(net697),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2016_ (.D(net803),
    .GATE(net697),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2017_ (.D(net802),
    .GATE(net697),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2018_ (.D(net800),
    .GATE(net697),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2019_ (.D(net797),
    .GATE(net697),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2020_ (.D(net796),
    .GATE(net697),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2021_ (.D(net794),
    .GATE(net698),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2022_ (.D(net792),
    .GATE(net698),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2023_ (.D(net788),
    .GATE(net698),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2024_ (.D(net786),
    .GATE(net698),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2025_ (.D(net783),
    .GATE(net697),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2026_ (.D(net781),
    .GATE(net697),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2027_ (.D(net780),
    .GATE(net697),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2028_ (.D(net778),
    .GATE(net697),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2029_ (.D(net776),
    .GATE(net695),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2030_ (.D(net773),
    .GATE(net695),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2031_ (.D(net770),
    .GATE(net695),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2032_ (.D(net768),
    .GATE(net695),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2033_ (.D(net763),
    .GATE(net695),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2034_ (.D(net761),
    .GATE(net695),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2035_ (.D(net812),
    .GATE(net699),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2036_ (.D(net790),
    .GATE(net699),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2037_ (.D(net766),
    .GATE(net699),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2038_ (.D(net759),
    .GATE(net699),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2039_ (.D(net757),
    .GATE(net700),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2040_ (.D(net755),
    .GATE(net700),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2041_ (.D(net754),
    .GATE(net699),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2042_ (.D(net752),
    .GATE(net699),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2043_ (.D(net750),
    .GATE(net699),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2044_ (.D(net748),
    .GATE(net699),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2045_ (.D(net810),
    .GATE(net701),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2046_ (.D(net808),
    .GATE(net701),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2047_ (.D(net805),
    .GATE(net702),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2048_ (.D(net803),
    .GATE(net702),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2049_ (.D(net802),
    .GATE(net701),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2050_ (.D(net800),
    .GATE(net701),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2051_ (.D(net797),
    .GATE(net701),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2052_ (.D(net795),
    .GATE(net701),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2053_ (.D(net794),
    .GATE(net701),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2054_ (.D(net792),
    .GATE(net701),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2055_ (.D(net788),
    .GATE(net701),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2056_ (.D(net786),
    .GATE(net701),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2057_ (.D(net783),
    .GATE(net702),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2058_ (.D(net781),
    .GATE(net702),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2059_ (.D(net780),
    .GATE(net702),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2060_ (.D(net778),
    .GATE(net702),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2061_ (.D(net774),
    .GATE(net700),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2062_ (.D(net771),
    .GATE(net700),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2063_ (.D(net769),
    .GATE(net700),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2064_ (.D(net767),
    .GATE(net700),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2065_ (.D(net763),
    .GATE(net699),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2066_ (.D(net761),
    .GATE(net699),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2067_ (.D(net812),
    .GATE(net744),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2068_ (.D(net790),
    .GATE(net744),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2069_ (.D(net766),
    .GATE(net745),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2070_ (.D(net759),
    .GATE(net745),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2071_ (.D(net757),
    .GATE(net743),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2072_ (.D(net755),
    .GATE(net743),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2073_ (.D(net754),
    .GATE(net745),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2074_ (.D(net752),
    .GATE(net745),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2075_ (.D(net749),
    .GATE(net744),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2076_ (.D(net747),
    .GATE(net744),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2077_ (.D(net29),
    .GATE(net746),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2078_ (.D(net30),
    .GATE(net746),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2079_ (.D(net806),
    .GATE(net743),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2080_ (.D(net804),
    .GATE(net743),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2081_ (.D(net802),
    .GATE(net743),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2082_ (.D(net800),
    .GATE(net743),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2083_ (.D(net797),
    .GATE(net743),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2084_ (.D(net795),
    .GATE(net743),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2085_ (.D(net37),
    .GATE(net746),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2086_ (.D(net38),
    .GATE(net746),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2087_ (.D(net788),
    .GATE(net746),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2088_ (.D(net786),
    .GATE(net746),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2089_ (.D(net783),
    .GATE(net746),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2090_ (.D(net781),
    .GATE(net746),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2091_ (.D(net780),
    .GATE(net743),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2092_ (.D(net778),
    .GATE(net743),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2093_ (.D(net774),
    .GATE(net744),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2094_ (.D(net771),
    .GATE(net744),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2095_ (.D(net769),
    .GATE(net744),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2096_ (.D(net767),
    .GATE(net744),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2097_ (.D(net764),
    .GATE(net744),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2098_ (.D(net762),
    .GATE(net744),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit31.Q ));
 sky130_fd_sc_hd__dfxtp_1 _2099_ (.CLK(clknet_1_1__leaf_UserCLK_regs),
    .D(_0000_),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.LUT_flop ));
 sky130_fd_sc_hd__dfxtp_1 _2100_ (.CLK(clknet_1_0__leaf_UserCLK_regs),
    .D(_0001_),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.LUT_flop ));
 sky130_fd_sc_hd__dfxtp_1 _2101_ (.CLK(clknet_1_0__leaf_UserCLK_regs),
    .D(_0002_),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.LUT_flop ));
 sky130_fd_sc_hd__dfxtp_1 _2102_ (.CLK(clknet_1_0__leaf_UserCLK_regs),
    .D(_0003_),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.LUT_flop ));
 sky130_fd_sc_hd__dfxtp_1 _2103_ (.CLK(clknet_1_0__leaf_UserCLK_regs),
    .D(_0004_),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.LUT_flop ));
 sky130_fd_sc_hd__dfxtp_1 _2104_ (.CLK(clknet_1_1__leaf_UserCLK_regs),
    .D(_0005_),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.LUT_flop ));
 sky130_fd_sc_hd__dfxtp_1 _2105_ (.CLK(clknet_1_1__leaf_UserCLK_regs),
    .D(_0006_),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.LUT_flop ));
 sky130_fd_sc_hd__dfxtp_1 _2106_ (.CLK(clknet_1_1__leaf_UserCLK_regs),
    .D(_0007_),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.LUT_flop ));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(E6END[6]));
 sky130_fd_sc_hd__buf_4 _2108_ (.A(\Inst_LUT4AB_switch_matrix.E1BEG1 ),
    .X(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(net155));
 sky130_fd_sc_hd__dlymetal6s2s_1 clone7 (.A(G),
    .X(net399));
 sky130_fd_sc_hd__buf_4 _2111_ (.A(\Inst_LUT4AB_switch_matrix.E2BEG0 ),
    .X(net144));
 sky130_fd_sc_hd__buf_4 _2112_ (.A(\Inst_LUT4AB_switch_matrix.E2BEG1 ),
    .X(net145));
 sky130_fd_sc_hd__clkbuf_2 _2113_ (.A(\Inst_LUT4AB_switch_matrix.E2BEG2 ),
    .X(net146));
 sky130_fd_sc_hd__buf_2 _2114_ (.A(\Inst_LUT4AB_switch_matrix.E2BEG3 ),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_2 _2115_ (.A(\Inst_LUT4AB_switch_matrix.E2BEG4 ),
    .X(net148));
 sky130_fd_sc_hd__buf_1 _2116_ (.A(\Inst_LUT4AB_switch_matrix.E2BEG5 ),
    .X(net149));
 sky130_fd_sc_hd__buf_6 _2117_ (.A(\Inst_LUT4AB_switch_matrix.E2BEG6 ),
    .X(net150));
 sky130_fd_sc_hd__buf_6 rebuffer55 (.A(net448),
    .X(net447));
 sky130_fd_sc_hd__clkbuf_2 _2119_ (.A(net14),
    .X(net152));
 sky130_fd_sc_hd__buf_1 _2120_ (.A(net15),
    .X(net153));
 sky130_fd_sc_hd__buf_1 _2121_ (.A(net16),
    .X(net154));
 sky130_fd_sc_hd__clkbuf_2 _2122_ (.A(net17),
    .X(net155));
 sky130_fd_sc_hd__clkbuf_2 _2123_ (.A(net18),
    .X(net156));
 sky130_fd_sc_hd__clkbuf_1 _2124_ (.A(net19),
    .X(net157));
 sky130_fd_sc_hd__buf_1 _2125_ (.A(net20),
    .X(net158));
 sky130_fd_sc_hd__buf_1 _2126_ (.A(net21),
    .X(net159));
 sky130_fd_sc_hd__clkbuf_1 _2127_ (.A(E6END[2]),
    .X(net160));
 sky130_fd_sc_hd__buf_1 _2128_ (.A(E6END[3]),
    .X(net163));
 sky130_fd_sc_hd__buf_1 _2129_ (.A(E6END[4]),
    .X(net164));
 sky130_fd_sc_hd__buf_1 _2130_ (.A(E6END[5]),
    .X(net165));
 sky130_fd_sc_hd__buf_1 _2131_ (.A(E6END[6]),
    .X(net166));
 sky130_fd_sc_hd__buf_1 _2132_ (.A(E6END[7]),
    .X(net167));
 sky130_fd_sc_hd__buf_1 _2133_ (.A(E6END[8]),
    .X(net168));
 sky130_fd_sc_hd__buf_1 _2134_ (.A(E6END[9]),
    .X(net169));
 sky130_fd_sc_hd__clkbuf_2 _2135_ (.A(E6END[10]),
    .X(net170));
 sky130_fd_sc_hd__clkbuf_2 _2136_ (.A(E6END[11]),
    .X(net171));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer41 (.A(net454),
    .X(net433));
 sky130_fd_sc_hd__buf_6 rebuffer39 (.A(_0107_),
    .X(net431));
 sky130_fd_sc_hd__clkbuf_1 _2139_ (.A(EE4END[4]),
    .X(net172));
 sky130_fd_sc_hd__clkbuf_1 _2140_ (.A(EE4END[5]),
    .X(net179));
 sky130_fd_sc_hd__clkbuf_1 _2141_ (.A(EE4END[6]),
    .X(net180));
 sky130_fd_sc_hd__clkbuf_1 _2142_ (.A(EE4END[7]),
    .X(net181));
 sky130_fd_sc_hd__clkbuf_1 _2143_ (.A(EE4END[8]),
    .X(net182));
 sky130_fd_sc_hd__clkbuf_1 _2144_ (.A(EE4END[9]),
    .X(net183));
 sky130_fd_sc_hd__clkbuf_1 _2145_ (.A(EE4END[10]),
    .X(net184));
 sky130_fd_sc_hd__clkbuf_1 _2146_ (.A(EE4END[11]),
    .X(net185));
 sky130_fd_sc_hd__clkbuf_1 _2147_ (.A(EE4END[12]),
    .X(net186));
 sky130_fd_sc_hd__buf_1 _2148_ (.A(EE4END[13]),
    .X(net187));
 sky130_fd_sc_hd__buf_1 _2149_ (.A(EE4END[14]),
    .X(net173));
 sky130_fd_sc_hd__buf_1 _2150_ (.A(EE4END[15]),
    .X(net174));
 sky130_fd_sc_hd__clkbuf_1 _2151_ (.A(\Inst_LUT4AB_switch_matrix.EE4BEG0 ),
    .X(net175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(\Inst_LC_LUT4c_frame_config_dffesr.LUT_flop ),
    .X(net486));
 sky130_fd_sc_hd__buf_1 _2153_ (.A(\Inst_LUT4AB_switch_matrix.EE4BEG2 ),
    .X(net177));
 sky130_fd_sc_hd__buf_6 rebuffer58 (.A(net451),
    .X(net450));
 sky130_fd_sc_hd__buf_1 _2155_ (.A(net811),
    .X(net188));
 sky130_fd_sc_hd__buf_1 _2156_ (.A(net789),
    .X(net199));
 sky130_fd_sc_hd__buf_1 _2157_ (.A(FrameData[2]),
    .X(net210));
 sky130_fd_sc_hd__buf_1 _2158_ (.A(net760),
    .X(net213));
 sky130_fd_sc_hd__clkbuf_1 _2159_ (.A(net758),
    .X(net214));
 sky130_fd_sc_hd__clkbuf_1 _2160_ (.A(net756),
    .X(net215));
 sky130_fd_sc_hd__buf_1 _2161_ (.A(net753),
    .X(net216));
 sky130_fd_sc_hd__buf_1 _2162_ (.A(net751),
    .X(net217));
 sky130_fd_sc_hd__buf_1 _2163_ (.A(net749),
    .X(net218));
 sky130_fd_sc_hd__buf_1 _2164_ (.A(net747),
    .X(net219));
 sky130_fd_sc_hd__buf_1 _2165_ (.A(net809),
    .X(net189));
 sky130_fd_sc_hd__buf_1 _2166_ (.A(net807),
    .X(net190));
 sky130_fd_sc_hd__buf_1 _2167_ (.A(net805),
    .X(net191));
 sky130_fd_sc_hd__buf_1 _2168_ (.A(net803),
    .X(net192));
 sky130_fd_sc_hd__buf_1 _2169_ (.A(net801),
    .X(net193));
 sky130_fd_sc_hd__buf_1 _2170_ (.A(net799),
    .X(net194));
 sky130_fd_sc_hd__clkbuf_1 _2171_ (.A(net798),
    .X(net195));
 sky130_fd_sc_hd__buf_1 _2172_ (.A(net796),
    .X(net196));
 sky130_fd_sc_hd__clkbuf_1 _2173_ (.A(net793),
    .X(net197));
 sky130_fd_sc_hd__buf_1 _2174_ (.A(net791),
    .X(net198));
 sky130_fd_sc_hd__clkbuf_1 _2175_ (.A(net787),
    .X(net200));
 sky130_fd_sc_hd__buf_1 _2176_ (.A(net785),
    .X(net201));
 sky130_fd_sc_hd__clkbuf_2 _2177_ (.A(net784),
    .X(net202));
 sky130_fd_sc_hd__buf_1 _2178_ (.A(net782),
    .X(net203));
 sky130_fd_sc_hd__clkbuf_1 _2179_ (.A(net779),
    .X(net204));
 sky130_fd_sc_hd__buf_1 _2180_ (.A(net777),
    .X(net205));
 sky130_fd_sc_hd__clkbuf_1 _2181_ (.A(net775),
    .X(net206));
 sky130_fd_sc_hd__clkbuf_2 _2182_ (.A(net771),
    .X(net207));
 sky130_fd_sc_hd__clkbuf_2 _2183_ (.A(net769),
    .X(net208));
 sky130_fd_sc_hd__clkbuf_1 _2184_ (.A(net767),
    .X(net209));
 sky130_fd_sc_hd__buf_1 _2185_ (.A(net764),
    .X(net211));
 sky130_fd_sc_hd__clkbuf_2 _2186_ (.A(net762),
    .X(net212));
 sky130_fd_sc_hd__clkbuf_2 _2187_ (.A(net746),
    .X(net220));
 sky130_fd_sc_hd__clkbuf_2 _2188_ (.A(FrameStrobe[1]),
    .X(net231));
 sky130_fd_sc_hd__clkbuf_2 _2189_ (.A(FrameStrobe[2]),
    .X(net232));
 sky130_fd_sc_hd__buf_1 _2190_ (.A(net693),
    .X(net233));
 sky130_fd_sc_hd__clkbuf_2 _2191_ (.A(net690),
    .X(net234));
 sky130_fd_sc_hd__buf_1 _2192_ (.A(net685),
    .X(net235));
 sky130_fd_sc_hd__buf_1 _2193_ (.A(net681),
    .X(net236));
 sky130_fd_sc_hd__buf_1 _2194_ (.A(net676),
    .X(net237));
 sky130_fd_sc_hd__clkbuf_1 _2195_ (.A(net671),
    .X(net238));
 sky130_fd_sc_hd__buf_1 _2196_ (.A(net669),
    .X(net239));
 sky130_fd_sc_hd__buf_1 _2197_ (.A(net742),
    .X(net221));
 sky130_fd_sc_hd__clkbuf_2 _2198_ (.A(net738),
    .X(net222));
 sky130_fd_sc_hd__buf_1 _2199_ (.A(net733),
    .X(net223));
 sky130_fd_sc_hd__buf_1 _2200_ (.A(net727),
    .X(net224));
 sky130_fd_sc_hd__clkbuf_1 _2201_ (.A(net725),
    .X(net225));
 sky130_fd_sc_hd__clkbuf_1 _2202_ (.A(net719),
    .X(net226));
 sky130_fd_sc_hd__buf_1 _2203_ (.A(FrameStrobe[16]),
    .X(net227));
 sky130_fd_sc_hd__buf_1 _2204_ (.A(net709),
    .X(net228));
 sky130_fd_sc_hd__buf_1 _2205_ (.A(net706),
    .X(net229));
 sky130_fd_sc_hd__clkbuf_2 _2206_ (.A(net55),
    .X(net230));
 sky130_fd_sc_hd__clkbuf_2 _2207_ (.A(\Inst_LUT4AB_switch_matrix.N1BEG0 ),
    .X(net240));
 sky130_fd_sc_hd__buf_4 _2208_ (.A(\Inst_LUT4AB_switch_matrix.N1BEG1 ),
    .X(net241));
 sky130_fd_sc_hd__clkbuf_2 _2209_ (.A(\Inst_LUT4AB_switch_matrix.N1BEG2 ),
    .X(net242));
 sky130_fd_sc_hd__buf_4 _2210_ (.A(\Inst_LUT4AB_switch_matrix.N1BEG3 ),
    .X(net243));
 sky130_fd_sc_hd__buf_4 _2211_ (.A(\Inst_LUT4AB_switch_matrix.JN2BEG0 ),
    .X(net244));
 sky130_fd_sc_hd__buf_8 _2212_ (.A(\Inst_LUT4AB_switch_matrix.JN2BEG1 ),
    .X(net245));
 sky130_fd_sc_hd__buf_8 _2213_ (.A(\Inst_LUT4AB_switch_matrix.JN2BEG2 ),
    .X(net246));
 sky130_fd_sc_hd__buf_6 _2214_ (.A(\Inst_LUT4AB_switch_matrix.JN2BEG3 ),
    .X(net247));
 sky130_fd_sc_hd__buf_4 _2215_ (.A(\Inst_LUT4AB_switch_matrix.JN2BEG4 ),
    .X(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(net141));
 sky130_fd_sc_hd__buf_1 _2217_ (.A(\Inst_LUT4AB_switch_matrix.JN2BEG6 ),
    .X(net250));
 sky130_fd_sc_hd__clkbuf_1 _2218_ (.A(\Inst_LUT4AB_switch_matrix.JN2BEG7 ),
    .X(net251));
 sky130_fd_sc_hd__buf_1 _2219_ (.A(net69),
    .X(net252));
 sky130_fd_sc_hd__buf_4 _2220_ (.A(net70),
    .X(net253));
 sky130_fd_sc_hd__clkbuf_2 _2221_ (.A(net71),
    .X(net254));
 sky130_fd_sc_hd__buf_4 _2222_ (.A(net72),
    .X(net255));
 sky130_fd_sc_hd__buf_1 _2223_ (.A(net73),
    .X(net256));
 sky130_fd_sc_hd__clkbuf_2 _2224_ (.A(net74),
    .X(net257));
 sky130_fd_sc_hd__clkbuf_2 _2225_ (.A(net75),
    .X(net258));
 sky130_fd_sc_hd__clkbuf_2 _2226_ (.A(net76),
    .X(net259));
 sky130_fd_sc_hd__clkbuf_1 _2227_ (.A(N4END[4]),
    .X(net260));
 sky130_fd_sc_hd__clkbuf_1 _2228_ (.A(N4END[5]),
    .X(net267));
 sky130_fd_sc_hd__clkbuf_1 _2229_ (.A(N4END[6]),
    .X(net268));
 sky130_fd_sc_hd__clkbuf_1 _2230_ (.A(N4END[7]),
    .X(net269));
 sky130_fd_sc_hd__clkbuf_1 _2231_ (.A(N4END[8]),
    .X(net270));
 sky130_fd_sc_hd__clkbuf_1 _2232_ (.A(N4END[9]),
    .X(net271));
 sky130_fd_sc_hd__clkbuf_1 _2233_ (.A(N4END[10]),
    .X(net272));
 sky130_fd_sc_hd__clkbuf_1 _2234_ (.A(N4END[11]),
    .X(net273));
 sky130_fd_sc_hd__clkbuf_1 _2235_ (.A(N4END[12]),
    .X(net274));
 sky130_fd_sc_hd__buf_1 _2236_ (.A(N4END[13]),
    .X(net275));
 sky130_fd_sc_hd__buf_1 _2237_ (.A(N4END[14]),
    .X(net261));
 sky130_fd_sc_hd__buf_1 _2238_ (.A(N4END[15]),
    .X(net262));
 sky130_fd_sc_hd__buf_4 _2239_ (.A(\Inst_LUT4AB_switch_matrix.N4BEG0 ),
    .X(net263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(\Inst_LF_LUT4c_frame_config_dffesr.LUT_flop ),
    .X(net482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(\Inst_LE_LUT4c_frame_config_dffesr.LUT_flop ),
    .X(net483));
 sky130_fd_sc_hd__clkbuf_2 _2242_ (.A(\Inst_LUT4AB_switch_matrix.N4BEG3 ),
    .X(net266));
 sky130_fd_sc_hd__buf_1 _2243_ (.A(NN4END[4]),
    .X(net276));
 sky130_fd_sc_hd__clkbuf_1 _2244_ (.A(NN4END[5]),
    .X(net283));
 sky130_fd_sc_hd__clkbuf_1 _2245_ (.A(NN4END[6]),
    .X(net284));
 sky130_fd_sc_hd__clkbuf_1 _2246_ (.A(NN4END[7]),
    .X(net285));
 sky130_fd_sc_hd__buf_1 _2247_ (.A(NN4END[8]),
    .X(net286));
 sky130_fd_sc_hd__buf_1 _2248_ (.A(NN4END[9]),
    .X(net287));
 sky130_fd_sc_hd__buf_1 _2249_ (.A(NN4END[10]),
    .X(net288));
 sky130_fd_sc_hd__buf_1 _2250_ (.A(NN4END[11]),
    .X(net289));
 sky130_fd_sc_hd__buf_1 _2251_ (.A(NN4END[12]),
    .X(net290));
 sky130_fd_sc_hd__buf_1 _2252_ (.A(NN4END[13]),
    .X(net291));
 sky130_fd_sc_hd__buf_1 _2253_ (.A(NN4END[14]),
    .X(net277));
 sky130_fd_sc_hd__buf_1 _2254_ (.A(NN4END[15]),
    .X(net278));
 sky130_fd_sc_hd__buf_1 _2255_ (.A(\Inst_LUT4AB_switch_matrix.NN4BEG0 ),
    .X(net279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(\Inst_LH_LUT4c_frame_config_dffesr.LUT_flop ),
    .X(net485));
 sky130_fd_sc_hd__clkbuf_1 _2257_ (.A(\Inst_LUT4AB_switch_matrix.NN4BEG2 ),
    .X(net281));
 sky130_fd_sc_hd__buf_6 rebuffer56 (.A(net449),
    .X(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(E6END[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(E6END[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(net171));
 sky130_fd_sc_hd__buf_6 _2263_ (.A(\Inst_LUT4AB_switch_matrix.JS2BEG0 ),
    .X(net296));
 sky130_fd_sc_hd__clkbuf_2 _2264_ (.A(\Inst_LUT4AB_switch_matrix.JS2BEG1 ),
    .X(net297));
 sky130_fd_sc_hd__clkbuf_2 _2265_ (.A(\Inst_LUT4AB_switch_matrix.JS2BEG2 ),
    .X(net298));
 sky130_fd_sc_hd__clkbuf_2 _2266_ (.A(\Inst_LUT4AB_switch_matrix.JS2BEG3 ),
    .X(net299));
 sky130_fd_sc_hd__clkbuf_2 _2267_ (.A(\Inst_LUT4AB_switch_matrix.JS2BEG4 ),
    .X(net300));
 sky130_fd_sc_hd__buf_2 _2268_ (.A(net408),
    .X(net301));
 sky130_fd_sc_hd__buf_4 _2269_ (.A(\Inst_LUT4AB_switch_matrix.JS2BEG6 ),
    .X(net302));
 sky130_fd_sc_hd__buf_6 _2270_ (.A(net400),
    .X(net303));
 sky130_fd_sc_hd__buf_1 _2271_ (.A(net97),
    .X(net304));
 sky130_fd_sc_hd__clkbuf_1 _2272_ (.A(net98),
    .X(net305));
 sky130_fd_sc_hd__buf_1 _2273_ (.A(net99),
    .X(net306));
 sky130_fd_sc_hd__clkbuf_1 _2274_ (.A(net100),
    .X(net307));
 sky130_fd_sc_hd__clkbuf_2 _2275_ (.A(net101),
    .X(net308));
 sky130_fd_sc_hd__buf_1 _2276_ (.A(net102),
    .X(net309));
 sky130_fd_sc_hd__buf_1 _2277_ (.A(net103),
    .X(net310));
 sky130_fd_sc_hd__buf_1 _2278_ (.A(net104),
    .X(net311));
 sky130_fd_sc_hd__clkbuf_2 _2279_ (.A(S4END[4]),
    .X(net312));
 sky130_fd_sc_hd__buf_2 _2280_ (.A(S4END[5]),
    .X(net319));
 sky130_fd_sc_hd__clkbuf_2 _2281_ (.A(S4END[6]),
    .X(net320));
 sky130_fd_sc_hd__clkbuf_2 _2282_ (.A(S4END[7]),
    .X(net321));
 sky130_fd_sc_hd__clkbuf_2 _2283_ (.A(S4END[8]),
    .X(net322));
 sky130_fd_sc_hd__clkbuf_2 _2284_ (.A(S4END[9]),
    .X(net323));
 sky130_fd_sc_hd__clkbuf_2 _2285_ (.A(S4END[10]),
    .X(net324));
 sky130_fd_sc_hd__clkbuf_2 _2286_ (.A(S4END[11]),
    .X(net325));
 sky130_fd_sc_hd__clkbuf_2 _2287_ (.A(S4END[12]),
    .X(net326));
 sky130_fd_sc_hd__clkbuf_2 _2288_ (.A(S4END[13]),
    .X(net327));
 sky130_fd_sc_hd__clkbuf_2 _2289_ (.A(S4END[14]),
    .X(net313));
 sky130_fd_sc_hd__clkbuf_2 _2290_ (.A(S4END[15]),
    .X(net314));
 sky130_fd_sc_hd__clkbuf_2 _2291_ (.A(\Inst_LUT4AB_switch_matrix.S4BEG0 ),
    .X(net315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(\Inst_LA_LUT4c_frame_config_dffesr.LUT_flop ),
    .X(net480));
 sky130_fd_sc_hd__buf_1 _2293_ (.A(\Inst_LUT4AB_switch_matrix.S4BEG2 ),
    .X(net317));
 sky130_fd_sc_hd__clkbuf_1 _2294_ (.A(\Inst_LUT4AB_switch_matrix.S4BEG3 ),
    .X(net318));
 sky130_fd_sc_hd__clkbuf_2 _2295_ (.A(SS4END[4]),
    .X(net328));
 sky130_fd_sc_hd__clkbuf_2 _2296_ (.A(SS4END[5]),
    .X(net335));
 sky130_fd_sc_hd__clkbuf_2 _2297_ (.A(SS4END[6]),
    .X(net336));
 sky130_fd_sc_hd__clkbuf_2 _2298_ (.A(SS4END[7]),
    .X(net337));
 sky130_fd_sc_hd__clkbuf_2 _2299_ (.A(SS4END[8]),
    .X(net338));
 sky130_fd_sc_hd__clkbuf_2 _2300_ (.A(SS4END[9]),
    .X(net339));
 sky130_fd_sc_hd__clkbuf_2 _2301_ (.A(SS4END[10]),
    .X(net340));
 sky130_fd_sc_hd__clkbuf_2 _2302_ (.A(SS4END[11]),
    .X(net341));
 sky130_fd_sc_hd__clkbuf_2 _2303_ (.A(SS4END[12]),
    .X(net342));
 sky130_fd_sc_hd__clkbuf_2 _2304_ (.A(SS4END[13]),
    .X(net343));
 sky130_fd_sc_hd__clkbuf_2 _2305_ (.A(SS4END[14]),
    .X(net329));
 sky130_fd_sc_hd__clkbuf_2 _2306_ (.A(SS4END[15]),
    .X(net330));
 sky130_fd_sc_hd__buf_1 _2307_ (.A(\Inst_LUT4AB_switch_matrix.SS4BEG0 ),
    .X(net331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(\Inst_LD_LUT4c_frame_config_dffesr.LUT_flop ),
    .X(net484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(\Inst_LG_LUT4c_frame_config_dffesr.LUT_flop ),
    .X(net481));
 sky130_fd_sc_hd__buf_6 _2310_ (.A(\Inst_LUT4AB_switch_matrix.SS4BEG3 ),
    .X(net334));
 sky130_fd_sc_hd__buf_2 _2311_ (.A(clknet_1_0__leaf_UserCLK),
    .X(net344));
 sky130_fd_sc_hd__buf_1 _2312_ (.A(\Inst_LUT4AB_switch_matrix.W1BEG0 ),
    .X(net345));
 sky130_fd_sc_hd__clkbuf_1 clone32 (.A(net643),
    .X(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(E6END[4]));
 sky130_fd_sc_hd__clkbuf_1 _2316_ (.A(\Inst_LUT4AB_switch_matrix.JW2BEG0 ),
    .X(net349));
 sky130_fd_sc_hd__clkbuf_1 _2317_ (.A(\Inst_LUT4AB_switch_matrix.JW2BEG1 ),
    .X(net350));
 sky130_fd_sc_hd__buf_6 _2318_ (.A(\Inst_LUT4AB_switch_matrix.JW2BEG2 ),
    .X(net351));
 sky130_fd_sc_hd__clkbuf_1 _2319_ (.A(\Inst_LUT4AB_switch_matrix.JW2BEG3 ),
    .X(net352));
 sky130_fd_sc_hd__buf_6 _2320_ (.A(\Inst_LUT4AB_switch_matrix.JW2BEG4 ),
    .X(net353));
 sky130_fd_sc_hd__buf_6 clone75 (.A(_0513_),
    .X(net467));
 sky130_fd_sc_hd__buf_6 _2322_ (.A(\Inst_LUT4AB_switch_matrix.JW2BEG6 ),
    .X(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(E6END[3]));
 sky130_fd_sc_hd__buf_1 _2324_ (.A(net125),
    .X(net357));
 sky130_fd_sc_hd__clkbuf_2 _2325_ (.A(net126),
    .X(net358));
 sky130_fd_sc_hd__clkbuf_2 _2326_ (.A(net127),
    .X(net359));
 sky130_fd_sc_hd__clkbuf_2 _2327_ (.A(net128),
    .X(net360));
 sky130_fd_sc_hd__buf_1 _2328_ (.A(net129),
    .X(net361));
 sky130_fd_sc_hd__clkbuf_2 _2329_ (.A(net130),
    .X(net362));
 sky130_fd_sc_hd__clkbuf_2 _2330_ (.A(net131),
    .X(net363));
 sky130_fd_sc_hd__clkbuf_2 _2331_ (.A(net132),
    .X(net364));
 sky130_fd_sc_hd__clkbuf_2 _2332_ (.A(W6END[2]),
    .X(net365));
 sky130_fd_sc_hd__clkbuf_2 _2333_ (.A(W6END[3]),
    .X(net368));
 sky130_fd_sc_hd__clkbuf_2 _2334_ (.A(W6END[4]),
    .X(net369));
 sky130_fd_sc_hd__clkbuf_2 _2335_ (.A(W6END[5]),
    .X(net370));
 sky130_fd_sc_hd__clkbuf_2 _2336_ (.A(W6END[6]),
    .X(net371));
 sky130_fd_sc_hd__clkbuf_2 _2337_ (.A(W6END[7]),
    .X(net372));
 sky130_fd_sc_hd__clkbuf_2 _2338_ (.A(W6END[8]),
    .X(net373));
 sky130_fd_sc_hd__clkbuf_2 _2339_ (.A(W6END[9]),
    .X(net374));
 sky130_fd_sc_hd__buf_4 _2340_ (.A(W6END[10]),
    .X(net375));
 sky130_fd_sc_hd__buf_4 _2341_ (.A(W6END[11]),
    .X(net376));
 sky130_fd_sc_hd__buf_6 rebuffer54 (.A(net447),
    .X(net446));
 sky130_fd_sc_hd__buf_6 rebuffer59 (.A(net452),
    .X(net451));
 sky130_fd_sc_hd__clkbuf_2 _2344_ (.A(WW4END[4]),
    .X(net377));
 sky130_fd_sc_hd__clkbuf_2 _2345_ (.A(WW4END[5]),
    .X(net384));
 sky130_fd_sc_hd__clkbuf_2 _2346_ (.A(WW4END[6]),
    .X(net385));
 sky130_fd_sc_hd__clkbuf_2 _2347_ (.A(WW4END[7]),
    .X(net386));
 sky130_fd_sc_hd__clkbuf_2 _2348_ (.A(WW4END[8]),
    .X(net387));
 sky130_fd_sc_hd__clkbuf_2 _2349_ (.A(WW4END[9]),
    .X(net388));
 sky130_fd_sc_hd__clkbuf_2 _2350_ (.A(WW4END[10]),
    .X(net389));
 sky130_fd_sc_hd__clkbuf_2 _2351_ (.A(WW4END[11]),
    .X(net390));
 sky130_fd_sc_hd__clkbuf_2 _2352_ (.A(WW4END[12]),
    .X(net391));
 sky130_fd_sc_hd__clkbuf_2 _2353_ (.A(WW4END[13]),
    .X(net392));
 sky130_fd_sc_hd__clkbuf_2 _2354_ (.A(WW4END[14]),
    .X(net378));
 sky130_fd_sc_hd__clkbuf_2 _2355_ (.A(WW4END[15]),
    .X(net379));
 sky130_fd_sc_hd__clkbuf_2 _2356_ (.A(\Inst_LUT4AB_switch_matrix.WW4BEG0 ),
    .X(net380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(\Inst_LB_LUT4c_frame_config_dffesr.LUT_flop ),
    .X(net487));
 sky130_fd_sc_hd__clkbuf_1 _2358_ (.A(\Inst_LUT4AB_switch_matrix.WW4BEG2 ),
    .X(net382));
 sky130_fd_sc_hd__buf_6 rebuffer57 (.A(net450),
    .X(net449));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_679 ();
 sky130_fd_sc_hd__buf_6 fanout621 (.A(_0513_),
    .X(net621));
 sky130_fd_sc_hd__buf_12 fanout622 (.A(\Inst_LUT4AB_switch_matrix.M_EF ),
    .X(net622));
 sky130_fd_sc_hd__buf_6 fanout623 (.A(\Inst_LUT4AB_switch_matrix.M_AB ),
    .X(net623));
 sky130_fd_sc_hd__buf_2 fanout624 (.A(net625),
    .X(net624));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout625 (.A(net626),
    .X(net625));
 sky130_fd_sc_hd__buf_2 fanout626 (.A(H),
    .X(net626));
 sky130_fd_sc_hd__buf_6 fanout627 (.A(net628),
    .X(net627));
 sky130_fd_sc_hd__buf_8 fanout628 (.A(H),
    .X(net628));
 sky130_fd_sc_hd__buf_2 fanout629 (.A(net630),
    .X(net629));
 sky130_fd_sc_hd__buf_8 fanout630 (.A(G),
    .X(net630));
 sky130_fd_sc_hd__buf_2 fanout631 (.A(net633),
    .X(net631));
 sky130_fd_sc_hd__buf_8 fanout632 (.A(net633),
    .X(net632));
 sky130_fd_sc_hd__buf_8 fanout633 (.A(G),
    .X(net633));
 sky130_fd_sc_hd__buf_8 fanout634 (.A(D),
    .X(net634));
 sky130_fd_sc_hd__buf_2 fanout635 (.A(D),
    .X(net635));
 sky130_fd_sc_hd__buf_2 fanout636 (.A(net637),
    .X(net636));
 sky130_fd_sc_hd__buf_4 fanout637 (.A(net638),
    .X(net637));
 sky130_fd_sc_hd__buf_6 fanout638 (.A(D),
    .X(net638));
 sky130_fd_sc_hd__buf_6 fanout639 (.A(net640),
    .X(net639));
 sky130_fd_sc_hd__buf_8 fanout640 (.A(net643),
    .X(net640));
 sky130_fd_sc_hd__buf_8 fanout641 (.A(net642),
    .X(net641));
 sky130_fd_sc_hd__buf_8 fanout642 (.A(net643),
    .X(net642));
 sky130_fd_sc_hd__buf_8 fanout643 (.A(F),
    .X(net643));
 sky130_fd_sc_hd__buf_4 fanout644 (.A(net645),
    .X(net644));
 sky130_fd_sc_hd__buf_2 fanout645 (.A(net648),
    .X(net645));
 sky130_fd_sc_hd__buf_2 fanout646 (.A(net647),
    .X(net646));
 sky130_fd_sc_hd__clkbuf_4 fanout647 (.A(net648),
    .X(net647));
 sky130_fd_sc_hd__buf_6 fanout648 (.A(E),
    .X(net648));
 sky130_fd_sc_hd__buf_4 fanout649 (.A(net651),
    .X(net649));
 sky130_fd_sc_hd__buf_1 fanout650 (.A(net651),
    .X(net650));
 sky130_fd_sc_hd__clkbuf_2 fanout651 (.A(C),
    .X(net651));
 sky130_fd_sc_hd__buf_2 fanout652 (.A(net653),
    .X(net652));
 sky130_fd_sc_hd__buf_2 fanout653 (.A(C),
    .X(net653));
 sky130_fd_sc_hd__buf_8 fanout654 (.A(net655),
    .X(net654));
 sky130_fd_sc_hd__buf_8 fanout655 (.A(B),
    .X(net655));
 sky130_fd_sc_hd__buf_2 fanout656 (.A(net657),
    .X(net656));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout657 (.A(net658),
    .X(net657));
 sky130_fd_sc_hd__clkbuf_4 fanout658 (.A(B),
    .X(net658));
 sky130_fd_sc_hd__buf_8 fanout659 (.A(net663),
    .X(net659));
 sky130_fd_sc_hd__buf_2 fanout660 (.A(net662),
    .X(net660));
 sky130_fd_sc_hd__buf_2 fanout661 (.A(net662),
    .X(net661));
 sky130_fd_sc_hd__clkbuf_2 fanout662 (.A(net663),
    .X(net662));
 sky130_fd_sc_hd__buf_8 fanout663 (.A(A),
    .X(net663));
 sky130_fd_sc_hd__clkbuf_4 fanout664 (.A(_0265_),
    .X(net664));
 sky130_fd_sc_hd__clkbuf_4 fanout665 (.A(net116),
    .X(net665));
 sky130_fd_sc_hd__clkbuf_4 fanout666 (.A(net115),
    .X(net666));
 sky130_fd_sc_hd__clkbuf_2 fanout667 (.A(net668),
    .X(net667));
 sky130_fd_sc_hd__clkbuf_2 fanout668 (.A(net669),
    .X(net668));
 sky130_fd_sc_hd__clkbuf_2 fanout669 (.A(net670),
    .X(net669));
 sky130_fd_sc_hd__buf_2 fanout670 (.A(FrameStrobe[9]),
    .X(net670));
 sky130_fd_sc_hd__clkbuf_2 fanout671 (.A(net672),
    .X(net671));
 sky130_fd_sc_hd__buf_1 fanout672 (.A(net673),
    .X(net672));
 sky130_fd_sc_hd__clkbuf_4 fanout673 (.A(FrameStrobe[8]),
    .X(net673));
 sky130_fd_sc_hd__buf_2 fanout674 (.A(FrameStrobe[8]),
    .X(net674));
 sky130_fd_sc_hd__buf_2 fanout675 (.A(net678),
    .X(net675));
 sky130_fd_sc_hd__clkbuf_2 fanout676 (.A(net677),
    .X(net676));
 sky130_fd_sc_hd__buf_2 fanout677 (.A(net678),
    .X(net677));
 sky130_fd_sc_hd__clkbuf_2 fanout678 (.A(FrameStrobe[7]),
    .X(net678));
 sky130_fd_sc_hd__clkbuf_2 fanout679 (.A(FrameStrobe[6]),
    .X(net679));
 sky130_fd_sc_hd__buf_1 fanout680 (.A(FrameStrobe[6]),
    .X(net680));
 sky130_fd_sc_hd__clkbuf_2 fanout681 (.A(net682),
    .X(net681));
 sky130_fd_sc_hd__clkbuf_4 fanout682 (.A(FrameStrobe[6]),
    .X(net682));
 sky130_fd_sc_hd__clkbuf_2 fanout683 (.A(net686),
    .X(net683));
 sky130_fd_sc_hd__buf_2 fanout684 (.A(net686),
    .X(net684));
 sky130_fd_sc_hd__buf_2 fanout685 (.A(net686),
    .X(net685));
 sky130_fd_sc_hd__clkbuf_2 fanout686 (.A(FrameStrobe[5]),
    .X(net686));
 sky130_fd_sc_hd__buf_2 fanout687 (.A(net56),
    .X(net687));
 sky130_fd_sc_hd__clkbuf_2 fanout688 (.A(net690),
    .X(net688));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout689 (.A(net690),
    .X(net689));
 sky130_fd_sc_hd__buf_2 fanout690 (.A(net56),
    .X(net690));
 sky130_fd_sc_hd__clkbuf_2 fanout691 (.A(net694),
    .X(net691));
 sky130_fd_sc_hd__clkbuf_2 fanout692 (.A(net693),
    .X(net692));
 sky130_fd_sc_hd__buf_2 fanout693 (.A(net694),
    .X(net693));
 sky130_fd_sc_hd__clkbuf_2 fanout694 (.A(FrameStrobe[3]),
    .X(net694));
 sky130_fd_sc_hd__clkbuf_2 fanout695 (.A(net696),
    .X(net695));
 sky130_fd_sc_hd__clkbuf_2 fanout696 (.A(FrameStrobe[2]),
    .X(net696));
 sky130_fd_sc_hd__buf_2 fanout697 (.A(net698),
    .X(net697));
 sky130_fd_sc_hd__clkbuf_2 fanout698 (.A(FrameStrobe[2]),
    .X(net698));
 sky130_fd_sc_hd__buf_2 fanout699 (.A(FrameStrobe[1]),
    .X(net699));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout700 (.A(FrameStrobe[1]),
    .X(net700));
 sky130_fd_sc_hd__clkbuf_2 fanout701 (.A(net702),
    .X(net701));
 sky130_fd_sc_hd__clkbuf_2 fanout702 (.A(FrameStrobe[1]),
    .X(net702));
 sky130_fd_sc_hd__clkbuf_2 fanout703 (.A(net704),
    .X(net703));
 sky130_fd_sc_hd__clkbuf_2 fanout704 (.A(FrameStrobe[18]),
    .X(net704));
 sky130_fd_sc_hd__clkbuf_2 fanout705 (.A(net706),
    .X(net705));
 sky130_fd_sc_hd__buf_1 fanout706 (.A(FrameStrobe[18]),
    .X(net706));
 sky130_fd_sc_hd__clkbuf_2 fanout707 (.A(net708),
    .X(net707));
 sky130_fd_sc_hd__clkbuf_1 fanout708 (.A(net711),
    .X(net708));
 sky130_fd_sc_hd__clkbuf_2 fanout709 (.A(net711),
    .X(net709));
 sky130_fd_sc_hd__clkbuf_1 fanout710 (.A(net711),
    .X(net710));
 sky130_fd_sc_hd__buf_1 fanout711 (.A(FrameStrobe[17]),
    .X(net711));
 sky130_fd_sc_hd__clkbuf_2 fanout712 (.A(net714),
    .X(net712));
 sky130_fd_sc_hd__buf_1 fanout713 (.A(net714),
    .X(net713));
 sky130_fd_sc_hd__buf_1 fanout714 (.A(net715),
    .X(net714));
 sky130_fd_sc_hd__buf_1 fanout715 (.A(net716),
    .X(net715));
 sky130_fd_sc_hd__clkbuf_2 fanout716 (.A(FrameStrobe[16]),
    .X(net716));
 sky130_fd_sc_hd__clkbuf_2 fanout717 (.A(net720),
    .X(net717));
 sky130_fd_sc_hd__clkbuf_2 fanout718 (.A(net719),
    .X(net718));
 sky130_fd_sc_hd__clkbuf_2 fanout719 (.A(net720),
    .X(net719));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout720 (.A(FrameStrobe[15]),
    .X(net720));
 sky130_fd_sc_hd__buf_2 fanout721 (.A(net725),
    .X(net721));
 sky130_fd_sc_hd__clkbuf_2 fanout722 (.A(net725),
    .X(net722));
 sky130_fd_sc_hd__clkbuf_2 fanout723 (.A(net724),
    .X(net723));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout724 (.A(net725),
    .X(net724));
 sky130_fd_sc_hd__clkbuf_2 fanout725 (.A(FrameStrobe[14]),
    .X(net725));
 sky130_fd_sc_hd__clkbuf_2 fanout726 (.A(net727),
    .X(net726));
 sky130_fd_sc_hd__clkbuf_2 fanout727 (.A(net729),
    .X(net727));
 sky130_fd_sc_hd__buf_2 fanout728 (.A(FrameStrobe[13]),
    .X(net728));
 sky130_fd_sc_hd__clkbuf_2 fanout729 (.A(FrameStrobe[13]),
    .X(net729));
 sky130_fd_sc_hd__clkbuf_2 fanout730 (.A(net732),
    .X(net730));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout731 (.A(net732),
    .X(net731));
 sky130_fd_sc_hd__clkbuf_2 fanout732 (.A(net734),
    .X(net732));
 sky130_fd_sc_hd__buf_2 fanout733 (.A(net734),
    .X(net733));
 sky130_fd_sc_hd__clkbuf_2 fanout734 (.A(FrameStrobe[12]),
    .X(net734));
 sky130_fd_sc_hd__clkbuf_2 fanout735 (.A(net736),
    .X(net735));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout736 (.A(net737),
    .X(net736));
 sky130_fd_sc_hd__buf_2 fanout737 (.A(net738),
    .X(net737));
 sky130_fd_sc_hd__clkbuf_2 fanout738 (.A(FrameStrobe[11]),
    .X(net738));
 sky130_fd_sc_hd__buf_2 fanout739 (.A(net741),
    .X(net739));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout740 (.A(net741),
    .X(net740));
 sky130_fd_sc_hd__clkbuf_2 fanout741 (.A(net742),
    .X(net741));
 sky130_fd_sc_hd__buf_2 fanout742 (.A(net54),
    .X(net742));
 sky130_fd_sc_hd__buf_2 fanout743 (.A(net745),
    .X(net743));
 sky130_fd_sc_hd__clkbuf_2 fanout744 (.A(net745),
    .X(net744));
 sky130_fd_sc_hd__clkbuf_2 fanout745 (.A(net746),
    .X(net745));
 sky130_fd_sc_hd__clkbuf_2 fanout746 (.A(FrameStrobe[0]),
    .X(net746));
 sky130_fd_sc_hd__clkbuf_4 fanout747 (.A(net748),
    .X(net747));
 sky130_fd_sc_hd__buf_4 fanout748 (.A(net53),
    .X(net748));
 sky130_fd_sc_hd__clkbuf_4 fanout749 (.A(net750),
    .X(net749));
 sky130_fd_sc_hd__buf_4 fanout750 (.A(net52),
    .X(net750));
 sky130_fd_sc_hd__clkbuf_4 fanout751 (.A(net752),
    .X(net751));
 sky130_fd_sc_hd__buf_4 fanout752 (.A(net51),
    .X(net752));
 sky130_fd_sc_hd__clkbuf_4 fanout753 (.A(net754),
    .X(net753));
 sky130_fd_sc_hd__buf_4 fanout754 (.A(net50),
    .X(net754));
 sky130_fd_sc_hd__clkbuf_4 fanout755 (.A(net756),
    .X(net755));
 sky130_fd_sc_hd__clkbuf_4 fanout756 (.A(net49),
    .X(net756));
 sky130_fd_sc_hd__clkbuf_4 fanout757 (.A(FrameData[4]),
    .X(net757));
 sky130_fd_sc_hd__clkbuf_4 fanout758 (.A(FrameData[4]),
    .X(net758));
 sky130_fd_sc_hd__clkbuf_4 fanout759 (.A(net760),
    .X(net759));
 sky130_fd_sc_hd__clkbuf_4 fanout760 (.A(net48),
    .X(net760));
 sky130_fd_sc_hd__clkbuf_4 fanout761 (.A(net762),
    .X(net761));
 sky130_fd_sc_hd__buf_4 fanout762 (.A(net47),
    .X(net762));
 sky130_fd_sc_hd__buf_4 fanout763 (.A(net764),
    .X(net763));
 sky130_fd_sc_hd__buf_4 fanout764 (.A(net46),
    .X(net764));
 sky130_fd_sc_hd__clkbuf_4 fanout765 (.A(net766),
    .X(net765));
 sky130_fd_sc_hd__buf_4 fanout766 (.A(FrameData[2]),
    .X(net766));
 sky130_fd_sc_hd__clkbuf_4 fanout767 (.A(net768),
    .X(net767));
 sky130_fd_sc_hd__buf_4 fanout768 (.A(net45),
    .X(net768));
 sky130_fd_sc_hd__buf_4 fanout769 (.A(net770),
    .X(net769));
 sky130_fd_sc_hd__buf_4 fanout770 (.A(net44),
    .X(net770));
 sky130_fd_sc_hd__clkbuf_4 fanout771 (.A(net773),
    .X(net771));
 sky130_fd_sc_hd__buf_2 fanout772 (.A(net773),
    .X(net772));
 sky130_fd_sc_hd__clkbuf_4 fanout773 (.A(FrameData[27]),
    .X(net773));
 sky130_fd_sc_hd__buf_4 fanout774 (.A(net776),
    .X(net774));
 sky130_fd_sc_hd__buf_2 fanout775 (.A(net776),
    .X(net775));
 sky130_fd_sc_hd__clkbuf_4 fanout776 (.A(FrameData[26]),
    .X(net776));
 sky130_fd_sc_hd__clkbuf_4 fanout777 (.A(net778),
    .X(net777));
 sky130_fd_sc_hd__buf_4 fanout778 (.A(net43),
    .X(net778));
 sky130_fd_sc_hd__buf_4 fanout779 (.A(net780),
    .X(net779));
 sky130_fd_sc_hd__buf_4 fanout780 (.A(net42),
    .X(net780));
 sky130_fd_sc_hd__clkbuf_4 fanout781 (.A(FrameData[23]),
    .X(net781));
 sky130_fd_sc_hd__buf_4 fanout782 (.A(FrameData[23]),
    .X(net782));
 sky130_fd_sc_hd__clkbuf_4 fanout783 (.A(FrameData[22]),
    .X(net783));
 sky130_fd_sc_hd__buf_4 fanout784 (.A(FrameData[22]),
    .X(net784));
 sky130_fd_sc_hd__buf_4 fanout785 (.A(net786),
    .X(net785));
 sky130_fd_sc_hd__buf_4 fanout786 (.A(net41),
    .X(net786));
 sky130_fd_sc_hd__clkbuf_4 fanout787 (.A(net788),
    .X(net787));
 sky130_fd_sc_hd__buf_4 fanout788 (.A(net40),
    .X(net788));
 sky130_fd_sc_hd__buf_4 fanout789 (.A(net790),
    .X(net789));
 sky130_fd_sc_hd__clkbuf_4 fanout790 (.A(net39),
    .X(net790));
 sky130_fd_sc_hd__clkbuf_4 fanout791 (.A(net792),
    .X(net791));
 sky130_fd_sc_hd__buf_4 fanout792 (.A(net38),
    .X(net792));
 sky130_fd_sc_hd__buf_4 fanout793 (.A(net794),
    .X(net793));
 sky130_fd_sc_hd__buf_4 fanout794 (.A(net37),
    .X(net794));
 sky130_fd_sc_hd__clkbuf_4 fanout795 (.A(net796),
    .X(net795));
 sky130_fd_sc_hd__buf_4 fanout796 (.A(net36),
    .X(net796));
 sky130_fd_sc_hd__clkbuf_4 fanout797 (.A(net798),
    .X(net797));
 sky130_fd_sc_hd__buf_4 fanout798 (.A(net35),
    .X(net798));
 sky130_fd_sc_hd__clkbuf_4 fanout799 (.A(net800),
    .X(net799));
 sky130_fd_sc_hd__buf_4 fanout800 (.A(net34),
    .X(net800));
 sky130_fd_sc_hd__clkbuf_4 fanout801 (.A(net802),
    .X(net801));
 sky130_fd_sc_hd__buf_4 fanout802 (.A(net33),
    .X(net802));
 sky130_fd_sc_hd__clkbuf_4 fanout803 (.A(net804),
    .X(net803));
 sky130_fd_sc_hd__buf_4 fanout804 (.A(net32),
    .X(net804));
 sky130_fd_sc_hd__clkbuf_4 fanout805 (.A(net806),
    .X(net805));
 sky130_fd_sc_hd__buf_4 fanout806 (.A(net31),
    .X(net806));
 sky130_fd_sc_hd__clkbuf_4 fanout807 (.A(net808),
    .X(net807));
 sky130_fd_sc_hd__clkbuf_4 fanout808 (.A(net30),
    .X(net808));
 sky130_fd_sc_hd__buf_4 fanout809 (.A(net810),
    .X(net809));
 sky130_fd_sc_hd__clkbuf_4 fanout810 (.A(net29),
    .X(net810));
 sky130_fd_sc_hd__buf_4 fanout811 (.A(net812),
    .X(net811));
 sky130_fd_sc_hd__buf_4 fanout812 (.A(net28),
    .X(net812));
 sky130_fd_sc_hd__buf_2 fanout813 (.A(net23),
    .X(net813));
 sky130_fd_sc_hd__buf_2 fanout814 (.A(net22),
    .X(net814));
 sky130_fd_sc_hd__clkbuf_4 fanout815 (.A(net5),
    .X(net815));
 sky130_fd_sc_hd__clkbuf_4 fanout816 (.A(net4),
    .X(net816));
 sky130_fd_sc_hd__buf_6 input1 (.A(Ci),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_4 input2 (.A(E1END[0]),
    .X(net2));
 sky130_fd_sc_hd__buf_2 input3 (.A(E1END[1]),
    .X(net3));
 sky130_fd_sc_hd__buf_1 input4 (.A(E1END[2]),
    .X(net4));
 sky130_fd_sc_hd__dlymetal6s2s_1 input5 (.A(E1END[3]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_2 input6 (.A(E2END[0]),
    .X(net6));
 sky130_fd_sc_hd__dlymetal6s2s_1 input7 (.A(E2END[1]),
    .X(net7));
 sky130_fd_sc_hd__buf_2 input8 (.A(E2END[2]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_2 input9 (.A(E2END[3]),
    .X(net9));
 sky130_fd_sc_hd__buf_1 input10 (.A(E2END[4]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_2 input11 (.A(E2END[5]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_2 input12 (.A(E2END[6]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_2 input13 (.A(E2END[7]),
    .X(net13));
 sky130_fd_sc_hd__buf_1 input14 (.A(E2MID[0]),
    .X(net14));
 sky130_fd_sc_hd__buf_2 input15 (.A(E2MID[1]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_2 input16 (.A(E2MID[2]),
    .X(net16));
 sky130_fd_sc_hd__buf_2 input17 (.A(E2MID[3]),
    .X(net17));
 sky130_fd_sc_hd__buf_1 input18 (.A(E2MID[4]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_2 input19 (.A(E2MID[5]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_2 input20 (.A(E2MID[6]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_2 input21 (.A(E2MID[7]),
    .X(net21));
 sky130_fd_sc_hd__dlymetal6s2s_1 input22 (.A(E6END[0]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_2 input23 (.A(E6END[1]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_2 input24 (.A(EE4END[0]),
    .X(net24));
 sky130_fd_sc_hd__dlymetal6s2s_1 input25 (.A(EE4END[1]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_2 input26 (.A(EE4END[2]),
    .X(net26));
 sky130_fd_sc_hd__dlymetal6s2s_1 input27 (.A(EE4END[3]),
    .X(net27));
 sky130_fd_sc_hd__dlymetal6s2s_1 input28 (.A(FrameData[0]),
    .X(net28));
 sky130_fd_sc_hd__dlymetal6s2s_1 input29 (.A(FrameData[10]),
    .X(net29));
 sky130_fd_sc_hd__dlymetal6s2s_1 input30 (.A(FrameData[11]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_2 input31 (.A(FrameData[12]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_2 input32 (.A(FrameData[13]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_2 input33 (.A(FrameData[14]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_2 input34 (.A(FrameData[15]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_2 input35 (.A(FrameData[16]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_2 input36 (.A(FrameData[17]),
    .X(net36));
 sky130_fd_sc_hd__buf_1 input37 (.A(FrameData[18]),
    .X(net37));
 sky130_fd_sc_hd__buf_1 input38 (.A(FrameData[19]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_2 input39 (.A(FrameData[1]),
    .X(net39));
 sky130_fd_sc_hd__buf_1 input40 (.A(FrameData[20]),
    .X(net40));
 sky130_fd_sc_hd__buf_1 input41 (.A(FrameData[21]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_2 input42 (.A(FrameData[24]),
    .X(net42));
 sky130_fd_sc_hd__buf_1 input43 (.A(FrameData[25]),
    .X(net43));
 sky130_fd_sc_hd__buf_2 input44 (.A(FrameData[28]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_2 input45 (.A(FrameData[29]),
    .X(net45));
 sky130_fd_sc_hd__buf_2 input46 (.A(FrameData[30]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_2 input47 (.A(FrameData[31]),
    .X(net47));
 sky130_fd_sc_hd__dlymetal6s2s_1 input48 (.A(FrameData[3]),
    .X(net48));
 sky130_fd_sc_hd__dlymetal6s2s_1 input49 (.A(FrameData[5]),
    .X(net49));
 sky130_fd_sc_hd__buf_1 input50 (.A(FrameData[6]),
    .X(net50));
 sky130_fd_sc_hd__buf_1 input51 (.A(FrameData[7]),
    .X(net51));
 sky130_fd_sc_hd__buf_1 input52 (.A(FrameData[8]),
    .X(net52));
 sky130_fd_sc_hd__buf_1 input53 (.A(FrameData[9]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_2 input54 (.A(FrameStrobe[10]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_2 input55 (.A(FrameStrobe[19]),
    .X(net55));
 sky130_fd_sc_hd__buf_2 input56 (.A(FrameStrobe[4]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_4 input57 (.A(N1END[0]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_4 input58 (.A(N1END[1]),
    .X(net58));
 sky130_fd_sc_hd__buf_4 input59 (.A(N1END[2]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_4 input60 (.A(N1END[3]),
    .X(net60));
 sky130_fd_sc_hd__buf_2 input61 (.A(N2END[0]),
    .X(net61));
 sky130_fd_sc_hd__dlymetal6s2s_1 input62 (.A(N2END[1]),
    .X(net62));
 sky130_fd_sc_hd__dlymetal6s2s_1 input63 (.A(N2END[2]),
    .X(net63));
 sky130_fd_sc_hd__buf_2 input64 (.A(N2END[3]),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_2 input65 (.A(N2END[4]),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_2 input66 (.A(N2END[5]),
    .X(net66));
 sky130_fd_sc_hd__buf_2 input67 (.A(N2END[6]),
    .X(net67));
 sky130_fd_sc_hd__buf_2 input68 (.A(N2END[7]),
    .X(net68));
 sky130_fd_sc_hd__dlymetal6s2s_1 input69 (.A(N2MID[0]),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_2 input70 (.A(N2MID[1]),
    .X(net70));
 sky130_fd_sc_hd__buf_2 input71 (.A(N2MID[2]),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_2 input72 (.A(N2MID[3]),
    .X(net72));
 sky130_fd_sc_hd__dlymetal6s2s_1 input73 (.A(N2MID[4]),
    .X(net73));
 sky130_fd_sc_hd__buf_2 input74 (.A(N2MID[5]),
    .X(net74));
 sky130_fd_sc_hd__buf_2 input75 (.A(N2MID[6]),
    .X(net75));
 sky130_fd_sc_hd__buf_2 input76 (.A(N2MID[7]),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_2 input77 (.A(N4END[0]),
    .X(net77));
 sky130_fd_sc_hd__dlymetal6s2s_1 input78 (.A(N4END[1]),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_2 input79 (.A(N4END[2]),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_2 input80 (.A(N4END[3]),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_2 input81 (.A(NN4END[0]),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_2 input82 (.A(NN4END[1]),
    .X(net82));
 sky130_fd_sc_hd__buf_1 input83 (.A(NN4END[2]),
    .X(net83));
 sky130_fd_sc_hd__dlymetal6s2s_1 input84 (.A(NN4END[3]),
    .X(net84));
 sky130_fd_sc_hd__buf_2 input85 (.A(S1END[0]),
    .X(net85));
 sky130_fd_sc_hd__buf_2 input86 (.A(S1END[1]),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_2 input87 (.A(S1END[2]),
    .X(net87));
 sky130_fd_sc_hd__buf_2 input88 (.A(S1END[3]),
    .X(net88));
 sky130_fd_sc_hd__buf_2 input89 (.A(S2END[0]),
    .X(net89));
 sky130_fd_sc_hd__buf_2 input90 (.A(S2END[1]),
    .X(net90));
 sky130_fd_sc_hd__buf_2 input91 (.A(S2END[2]),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_2 input92 (.A(S2END[3]),
    .X(net92));
 sky130_fd_sc_hd__buf_2 input93 (.A(S2END[4]),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_2 input94 (.A(S2END[5]),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_2 input95 (.A(S2END[6]),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_2 input96 (.A(S2END[7]),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_2 input97 (.A(S2MID[0]),
    .X(net97));
 sky130_fd_sc_hd__buf_2 input98 (.A(S2MID[1]),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_2 input99 (.A(S2MID[2]),
    .X(net99));
 sky130_fd_sc_hd__buf_2 input100 (.A(S2MID[3]),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_2 input101 (.A(S2MID[4]),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_2 input102 (.A(S2MID[5]),
    .X(net102));
 sky130_fd_sc_hd__dlymetal6s2s_1 input103 (.A(S2MID[6]),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_2 input104 (.A(S2MID[7]),
    .X(net104));
 sky130_fd_sc_hd__buf_2 input105 (.A(S4END[0]),
    .X(net105));
 sky130_fd_sc_hd__buf_2 input106 (.A(S4END[1]),
    .X(net106));
 sky130_fd_sc_hd__buf_2 input107 (.A(S4END[2]),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_2 input108 (.A(S4END[3]),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_2 input109 (.A(SS4END[0]),
    .X(net109));
 sky130_fd_sc_hd__buf_2 input110 (.A(SS4END[1]),
    .X(net110));
 sky130_fd_sc_hd__buf_2 input111 (.A(SS4END[2]),
    .X(net111));
 sky130_fd_sc_hd__dlymetal6s2s_1 input112 (.A(SS4END[3]),
    .X(net112));
 sky130_fd_sc_hd__buf_4 input113 (.A(W1END[0]),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_4 input114 (.A(W1END[1]),
    .X(net114));
 sky130_fd_sc_hd__buf_2 input115 (.A(W1END[2]),
    .X(net115));
 sky130_fd_sc_hd__clkbuf_2 input116 (.A(W1END[3]),
    .X(net116));
 sky130_fd_sc_hd__clkbuf_2 input117 (.A(W2END[0]),
    .X(net117));
 sky130_fd_sc_hd__buf_2 input118 (.A(W2END[1]),
    .X(net118));
 sky130_fd_sc_hd__buf_2 input119 (.A(W2END[2]),
    .X(net119));
 sky130_fd_sc_hd__buf_2 input120 (.A(W2END[3]),
    .X(net120));
 sky130_fd_sc_hd__buf_2 input121 (.A(W2END[4]),
    .X(net121));
 sky130_fd_sc_hd__clkbuf_2 input122 (.A(W2END[5]),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_2 input123 (.A(W2END[6]),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_2 input124 (.A(W2END[7]),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_2 input125 (.A(W2MID[0]),
    .X(net125));
 sky130_fd_sc_hd__dlymetal6s2s_1 input126 (.A(W2MID[1]),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_2 input127 (.A(W2MID[2]),
    .X(net127));
 sky130_fd_sc_hd__clkbuf_2 input128 (.A(W2MID[3]),
    .X(net128));
 sky130_fd_sc_hd__buf_2 input129 (.A(W2MID[4]),
    .X(net129));
 sky130_fd_sc_hd__clkbuf_2 input130 (.A(W2MID[5]),
    .X(net130));
 sky130_fd_sc_hd__clkbuf_2 input131 (.A(W2MID[6]),
    .X(net131));
 sky130_fd_sc_hd__dlymetal6s2s_1 input132 (.A(W2MID[7]),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_4 input133 (.A(W6END[0]),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_4 input134 (.A(W6END[1]),
    .X(net134));
 sky130_fd_sc_hd__buf_2 input135 (.A(WW4END[0]),
    .X(net135));
 sky130_fd_sc_hd__clkbuf_2 input136 (.A(WW4END[1]),
    .X(net136));
 sky130_fd_sc_hd__buf_2 input137 (.A(WW4END[2]),
    .X(net137));
 sky130_fd_sc_hd__clkbuf_2 input138 (.A(WW4END[3]),
    .X(net138));
 sky130_fd_sc_hd__buf_6 output139 (.A(net139),
    .X(Co));
 sky130_fd_sc_hd__buf_8 output140 (.A(\Inst_LUT4AB_switch_matrix.E1BEG0 ),
    .X(E1BEG[0]));
 sky130_fd_sc_hd__buf_4 output141 (.A(net141),
    .X(E1BEG[1]));
 sky130_fd_sc_hd__buf_6 output142 (.A(\Inst_LUT4AB_switch_matrix.E1BEG2 ),
    .X(E1BEG[2]));
 sky130_fd_sc_hd__buf_8 output143 (.A(\Inst_LUT4AB_switch_matrix.E1BEG3 ),
    .X(E1BEG[3]));
 sky130_fd_sc_hd__buf_6 output144 (.A(net144),
    .X(E2BEG[0]));
 sky130_fd_sc_hd__buf_4 output145 (.A(net145),
    .X(E2BEG[1]));
 sky130_fd_sc_hd__buf_6 output146 (.A(net146),
    .X(E2BEG[2]));
 sky130_fd_sc_hd__buf_4 output147 (.A(net147),
    .X(E2BEG[3]));
 sky130_fd_sc_hd__buf_2 output148 (.A(net148),
    .X(E2BEG[4]));
 sky130_fd_sc_hd__buf_4 output149 (.A(net149),
    .X(E2BEG[5]));
 sky130_fd_sc_hd__buf_8 output150 (.A(net150),
    .X(E2BEG[6]));
 sky130_fd_sc_hd__buf_8 output151 (.A(\Inst_LUT4AB_switch_matrix.E2BEG7 ),
    .X(E2BEG[7]));
 sky130_fd_sc_hd__buf_2 output152 (.A(net152),
    .X(E2BEGb[0]));
 sky130_fd_sc_hd__buf_2 output153 (.A(net153),
    .X(E2BEGb[1]));
 sky130_fd_sc_hd__buf_2 output154 (.A(net154),
    .X(E2BEGb[2]));
 sky130_fd_sc_hd__buf_2 output155 (.A(net155),
    .X(E2BEGb[3]));
 sky130_fd_sc_hd__buf_2 output156 (.A(net156),
    .X(E2BEGb[4]));
 sky130_fd_sc_hd__buf_2 output157 (.A(net157),
    .X(E2BEGb[5]));
 sky130_fd_sc_hd__buf_2 output158 (.A(net158),
    .X(E2BEGb[6]));
 sky130_fd_sc_hd__buf_2 output159 (.A(net159),
    .X(E2BEGb[7]));
 sky130_fd_sc_hd__buf_2 output160 (.A(net160),
    .X(E6BEG[0]));
 sky130_fd_sc_hd__buf_8 output161 (.A(\Inst_LUT4AB_switch_matrix.E6BEG0 ),
    .X(E6BEG[10]));
 sky130_fd_sc_hd__buf_6 output162 (.A(\Inst_LUT4AB_switch_matrix.E6BEG1 ),
    .X(E6BEG[11]));
 sky130_fd_sc_hd__buf_2 output163 (.A(net163),
    .X(E6BEG[1]));
 sky130_fd_sc_hd__buf_2 output164 (.A(net164),
    .X(E6BEG[2]));
 sky130_fd_sc_hd__buf_2 output165 (.A(net165),
    .X(E6BEG[3]));
 sky130_fd_sc_hd__buf_2 output166 (.A(net166),
    .X(E6BEG[4]));
 sky130_fd_sc_hd__buf_2 output167 (.A(net167),
    .X(E6BEG[5]));
 sky130_fd_sc_hd__buf_2 output168 (.A(net168),
    .X(E6BEG[6]));
 sky130_fd_sc_hd__buf_2 output169 (.A(net169),
    .X(E6BEG[7]));
 sky130_fd_sc_hd__buf_2 output170 (.A(net170),
    .X(E6BEG[8]));
 sky130_fd_sc_hd__buf_2 output171 (.A(net171),
    .X(E6BEG[9]));
 sky130_fd_sc_hd__buf_2 output172 (.A(net172),
    .X(EE4BEG[0]));
 sky130_fd_sc_hd__buf_2 output173 (.A(net173),
    .X(EE4BEG[10]));
 sky130_fd_sc_hd__buf_2 output174 (.A(net174),
    .X(EE4BEG[11]));
 sky130_fd_sc_hd__buf_4 output175 (.A(net175),
    .X(EE4BEG[12]));
 sky130_fd_sc_hd__buf_8 output176 (.A(\Inst_LUT4AB_switch_matrix.EE4BEG1 ),
    .X(EE4BEG[13]));
 sky130_fd_sc_hd__buf_4 output177 (.A(net177),
    .X(EE4BEG[14]));
 sky130_fd_sc_hd__buf_6 output178 (.A(\Inst_LUT4AB_switch_matrix.EE4BEG3 ),
    .X(EE4BEG[15]));
 sky130_fd_sc_hd__buf_2 output179 (.A(net179),
    .X(EE4BEG[1]));
 sky130_fd_sc_hd__buf_2 output180 (.A(net180),
    .X(EE4BEG[2]));
 sky130_fd_sc_hd__buf_2 output181 (.A(net181),
    .X(EE4BEG[3]));
 sky130_fd_sc_hd__buf_2 output182 (.A(net182),
    .X(EE4BEG[4]));
 sky130_fd_sc_hd__buf_2 output183 (.A(net183),
    .X(EE4BEG[5]));
 sky130_fd_sc_hd__buf_2 output184 (.A(net184),
    .X(EE4BEG[6]));
 sky130_fd_sc_hd__buf_2 output185 (.A(net185),
    .X(EE4BEG[7]));
 sky130_fd_sc_hd__buf_2 output186 (.A(net186),
    .X(EE4BEG[8]));
 sky130_fd_sc_hd__buf_2 output187 (.A(net187),
    .X(EE4BEG[9]));
 sky130_fd_sc_hd__buf_2 output188 (.A(net188),
    .X(FrameData_O[0]));
 sky130_fd_sc_hd__buf_2 output189 (.A(net189),
    .X(FrameData_O[10]));
 sky130_fd_sc_hd__buf_2 output190 (.A(net190),
    .X(FrameData_O[11]));
 sky130_fd_sc_hd__buf_2 output191 (.A(net191),
    .X(FrameData_O[12]));
 sky130_fd_sc_hd__buf_2 output192 (.A(net192),
    .X(FrameData_O[13]));
 sky130_fd_sc_hd__buf_2 output193 (.A(net193),
    .X(FrameData_O[14]));
 sky130_fd_sc_hd__buf_2 output194 (.A(net194),
    .X(FrameData_O[15]));
 sky130_fd_sc_hd__buf_2 output195 (.A(net195),
    .X(FrameData_O[16]));
 sky130_fd_sc_hd__buf_2 output196 (.A(net196),
    .X(FrameData_O[17]));
 sky130_fd_sc_hd__buf_2 output197 (.A(net197),
    .X(FrameData_O[18]));
 sky130_fd_sc_hd__buf_2 output198 (.A(net198),
    .X(FrameData_O[19]));
 sky130_fd_sc_hd__buf_2 output199 (.A(net199),
    .X(FrameData_O[1]));
 sky130_fd_sc_hd__buf_2 output200 (.A(net200),
    .X(FrameData_O[20]));
 sky130_fd_sc_hd__buf_2 output201 (.A(net201),
    .X(FrameData_O[21]));
 sky130_fd_sc_hd__buf_2 output202 (.A(net202),
    .X(FrameData_O[22]));
 sky130_fd_sc_hd__buf_2 output203 (.A(net203),
    .X(FrameData_O[23]));
 sky130_fd_sc_hd__buf_2 output204 (.A(net204),
    .X(FrameData_O[24]));
 sky130_fd_sc_hd__buf_2 output205 (.A(net205),
    .X(FrameData_O[25]));
 sky130_fd_sc_hd__buf_2 output206 (.A(net206),
    .X(FrameData_O[26]));
 sky130_fd_sc_hd__buf_2 output207 (.A(net207),
    .X(FrameData_O[27]));
 sky130_fd_sc_hd__buf_2 output208 (.A(net208),
    .X(FrameData_O[28]));
 sky130_fd_sc_hd__buf_2 output209 (.A(net209),
    .X(FrameData_O[29]));
 sky130_fd_sc_hd__buf_2 output210 (.A(net210),
    .X(FrameData_O[2]));
 sky130_fd_sc_hd__buf_2 output211 (.A(net211),
    .X(FrameData_O[30]));
 sky130_fd_sc_hd__buf_2 output212 (.A(net212),
    .X(FrameData_O[31]));
 sky130_fd_sc_hd__buf_2 output213 (.A(net213),
    .X(FrameData_O[3]));
 sky130_fd_sc_hd__buf_2 output214 (.A(net214),
    .X(FrameData_O[4]));
 sky130_fd_sc_hd__buf_2 output215 (.A(net215),
    .X(FrameData_O[5]));
 sky130_fd_sc_hd__buf_2 output216 (.A(net216),
    .X(FrameData_O[6]));
 sky130_fd_sc_hd__buf_2 output217 (.A(net217),
    .X(FrameData_O[7]));
 sky130_fd_sc_hd__buf_2 output218 (.A(net218),
    .X(FrameData_O[8]));
 sky130_fd_sc_hd__buf_2 output219 (.A(net219),
    .X(FrameData_O[9]));
 sky130_fd_sc_hd__buf_2 output220 (.A(net220),
    .X(FrameStrobe_O[0]));
 sky130_fd_sc_hd__buf_2 output221 (.A(net221),
    .X(FrameStrobe_O[10]));
 sky130_fd_sc_hd__buf_2 output222 (.A(net222),
    .X(FrameStrobe_O[11]));
 sky130_fd_sc_hd__buf_2 output223 (.A(net223),
    .X(FrameStrobe_O[12]));
 sky130_fd_sc_hd__buf_2 output224 (.A(net224),
    .X(FrameStrobe_O[13]));
 sky130_fd_sc_hd__buf_2 output225 (.A(net225),
    .X(FrameStrobe_O[14]));
 sky130_fd_sc_hd__buf_2 output226 (.A(net226),
    .X(FrameStrobe_O[15]));
 sky130_fd_sc_hd__buf_2 output227 (.A(net227),
    .X(FrameStrobe_O[16]));
 sky130_fd_sc_hd__buf_2 output228 (.A(net228),
    .X(FrameStrobe_O[17]));
 sky130_fd_sc_hd__buf_2 output229 (.A(net229),
    .X(FrameStrobe_O[18]));
 sky130_fd_sc_hd__buf_2 output230 (.A(net230),
    .X(FrameStrobe_O[19]));
 sky130_fd_sc_hd__buf_2 output231 (.A(net231),
    .X(FrameStrobe_O[1]));
 sky130_fd_sc_hd__buf_2 output232 (.A(net232),
    .X(FrameStrobe_O[2]));
 sky130_fd_sc_hd__buf_2 output233 (.A(net233),
    .X(FrameStrobe_O[3]));
 sky130_fd_sc_hd__buf_2 output234 (.A(net234),
    .X(FrameStrobe_O[4]));
 sky130_fd_sc_hd__buf_2 output235 (.A(net235),
    .X(FrameStrobe_O[5]));
 sky130_fd_sc_hd__buf_2 output236 (.A(net236),
    .X(FrameStrobe_O[6]));
 sky130_fd_sc_hd__buf_2 output237 (.A(net237),
    .X(FrameStrobe_O[7]));
 sky130_fd_sc_hd__buf_2 output238 (.A(net238),
    .X(FrameStrobe_O[8]));
 sky130_fd_sc_hd__buf_2 output239 (.A(net239),
    .X(FrameStrobe_O[9]));
 sky130_fd_sc_hd__clkbuf_4 output240 (.A(net240),
    .X(N1BEG[0]));
 sky130_fd_sc_hd__buf_4 output241 (.A(net241),
    .X(N1BEG[1]));
 sky130_fd_sc_hd__buf_4 output242 (.A(net242),
    .X(N1BEG[2]));
 sky130_fd_sc_hd__buf_4 output243 (.A(net243),
    .X(N1BEG[3]));
 sky130_fd_sc_hd__buf_6 output244 (.A(net244),
    .X(N2BEG[0]));
 sky130_fd_sc_hd__buf_8 output245 (.A(net245),
    .X(N2BEG[1]));
 sky130_fd_sc_hd__buf_8 output246 (.A(net246),
    .X(N2BEG[2]));
 sky130_fd_sc_hd__buf_6 output247 (.A(net247),
    .X(N2BEG[3]));
 sky130_fd_sc_hd__buf_6 output248 (.A(net248),
    .X(N2BEG[4]));
 sky130_fd_sc_hd__buf_6 output249 (.A(\Inst_LUT4AB_switch_matrix.JN2BEG5 ),
    .X(N2BEG[5]));
 sky130_fd_sc_hd__buf_6 output250 (.A(net250),
    .X(N2BEG[6]));
 sky130_fd_sc_hd__buf_2 output251 (.A(net251),
    .X(N2BEG[7]));
 sky130_fd_sc_hd__buf_2 output252 (.A(net252),
    .X(N2BEGb[0]));
 sky130_fd_sc_hd__buf_2 output253 (.A(net253),
    .X(N2BEGb[1]));
 sky130_fd_sc_hd__buf_2 output254 (.A(net254),
    .X(N2BEGb[2]));
 sky130_fd_sc_hd__buf_2 output255 (.A(net255),
    .X(N2BEGb[3]));
 sky130_fd_sc_hd__buf_2 output256 (.A(net256),
    .X(N2BEGb[4]));
 sky130_fd_sc_hd__buf_2 output257 (.A(net257),
    .X(N2BEGb[5]));
 sky130_fd_sc_hd__buf_2 output258 (.A(net258),
    .X(N2BEGb[6]));
 sky130_fd_sc_hd__buf_2 output259 (.A(net259),
    .X(N2BEGb[7]));
 sky130_fd_sc_hd__buf_2 output260 (.A(net260),
    .X(N4BEG[0]));
 sky130_fd_sc_hd__buf_2 output261 (.A(net261),
    .X(N4BEG[10]));
 sky130_fd_sc_hd__buf_2 output262 (.A(net262),
    .X(N4BEG[11]));
 sky130_fd_sc_hd__buf_4 output263 (.A(net263),
    .X(N4BEG[12]));
 sky130_fd_sc_hd__buf_6 output264 (.A(\Inst_LUT4AB_switch_matrix.N4BEG1 ),
    .X(N4BEG[13]));
 sky130_fd_sc_hd__buf_4 output265 (.A(\Inst_LUT4AB_switch_matrix.N4BEG2 ),
    .X(N4BEG[14]));
 sky130_fd_sc_hd__buf_4 output266 (.A(net266),
    .X(N4BEG[15]));
 sky130_fd_sc_hd__buf_2 output267 (.A(net267),
    .X(N4BEG[1]));
 sky130_fd_sc_hd__buf_2 output268 (.A(net268),
    .X(N4BEG[2]));
 sky130_fd_sc_hd__buf_2 output269 (.A(net269),
    .X(N4BEG[3]));
 sky130_fd_sc_hd__buf_2 output270 (.A(net270),
    .X(N4BEG[4]));
 sky130_fd_sc_hd__buf_2 output271 (.A(net271),
    .X(N4BEG[5]));
 sky130_fd_sc_hd__buf_2 output272 (.A(net272),
    .X(N4BEG[6]));
 sky130_fd_sc_hd__buf_2 output273 (.A(net273),
    .X(N4BEG[7]));
 sky130_fd_sc_hd__buf_2 output274 (.A(net274),
    .X(N4BEG[8]));
 sky130_fd_sc_hd__buf_2 output275 (.A(net275),
    .X(N4BEG[9]));
 sky130_fd_sc_hd__buf_2 output276 (.A(net276),
    .X(NN4BEG[0]));
 sky130_fd_sc_hd__buf_2 output277 (.A(net277),
    .X(NN4BEG[10]));
 sky130_fd_sc_hd__buf_2 output278 (.A(net278),
    .X(NN4BEG[11]));
 sky130_fd_sc_hd__buf_4 output279 (.A(net279),
    .X(NN4BEG[12]));
 sky130_fd_sc_hd__buf_6 output280 (.A(\Inst_LUT4AB_switch_matrix.NN4BEG1 ),
    .X(NN4BEG[13]));
 sky130_fd_sc_hd__clkbuf_4 output281 (.A(net281),
    .X(NN4BEG[14]));
 sky130_fd_sc_hd__buf_8 output282 (.A(\Inst_LUT4AB_switch_matrix.NN4BEG3 ),
    .X(NN4BEG[15]));
 sky130_fd_sc_hd__buf_2 output283 (.A(net283),
    .X(NN4BEG[1]));
 sky130_fd_sc_hd__buf_2 output284 (.A(net284),
    .X(NN4BEG[2]));
 sky130_fd_sc_hd__buf_2 output285 (.A(net285),
    .X(NN4BEG[3]));
 sky130_fd_sc_hd__buf_2 output286 (.A(net286),
    .X(NN4BEG[4]));
 sky130_fd_sc_hd__buf_2 output287 (.A(net287),
    .X(NN4BEG[5]));
 sky130_fd_sc_hd__buf_2 output288 (.A(net288),
    .X(NN4BEG[6]));
 sky130_fd_sc_hd__buf_2 output289 (.A(net289),
    .X(NN4BEG[7]));
 sky130_fd_sc_hd__buf_2 output290 (.A(net290),
    .X(NN4BEG[8]));
 sky130_fd_sc_hd__buf_2 output291 (.A(net291),
    .X(NN4BEG[9]));
 sky130_fd_sc_hd__buf_8 output292 (.A(\Inst_LUT4AB_switch_matrix.S1BEG0 ),
    .X(S1BEG[0]));
 sky130_fd_sc_hd__buf_6 output293 (.A(\Inst_LUT4AB_switch_matrix.S1BEG1 ),
    .X(S1BEG[1]));
 sky130_fd_sc_hd__buf_6 output294 (.A(\Inst_LUT4AB_switch_matrix.S1BEG2 ),
    .X(S1BEG[2]));
 sky130_fd_sc_hd__buf_6 output295 (.A(\Inst_LUT4AB_switch_matrix.S1BEG3 ),
    .X(S1BEG[3]));
 sky130_fd_sc_hd__buf_8 output296 (.A(net296),
    .X(S2BEG[0]));
 sky130_fd_sc_hd__buf_6 output297 (.A(net297),
    .X(S2BEG[1]));
 sky130_fd_sc_hd__buf_6 output298 (.A(net298),
    .X(S2BEG[2]));
 sky130_fd_sc_hd__buf_4 output299 (.A(net299),
    .X(S2BEG[3]));
 sky130_fd_sc_hd__buf_4 output300 (.A(net300),
    .X(S2BEG[4]));
 sky130_fd_sc_hd__buf_6 output301 (.A(net301),
    .X(S2BEG[5]));
 sky130_fd_sc_hd__buf_4 output302 (.A(net302),
    .X(S2BEG[6]));
 sky130_fd_sc_hd__buf_8 output303 (.A(net303),
    .X(S2BEG[7]));
 sky130_fd_sc_hd__buf_2 output304 (.A(net304),
    .X(S2BEGb[0]));
 sky130_fd_sc_hd__buf_2 output305 (.A(net305),
    .X(S2BEGb[1]));
 sky130_fd_sc_hd__buf_2 output306 (.A(net306),
    .X(S2BEGb[2]));
 sky130_fd_sc_hd__buf_2 output307 (.A(net307),
    .X(S2BEGb[3]));
 sky130_fd_sc_hd__buf_2 output308 (.A(net308),
    .X(S2BEGb[4]));
 sky130_fd_sc_hd__buf_2 output309 (.A(net309),
    .X(S2BEGb[5]));
 sky130_fd_sc_hd__buf_2 output310 (.A(net310),
    .X(S2BEGb[6]));
 sky130_fd_sc_hd__buf_2 output311 (.A(net311),
    .X(S2BEGb[7]));
 sky130_fd_sc_hd__buf_2 output312 (.A(net312),
    .X(S4BEG[0]));
 sky130_fd_sc_hd__buf_2 output313 (.A(net313),
    .X(S4BEG[10]));
 sky130_fd_sc_hd__buf_2 output314 (.A(net314),
    .X(S4BEG[11]));
 sky130_fd_sc_hd__buf_4 output315 (.A(net315),
    .X(S4BEG[12]));
 sky130_fd_sc_hd__buf_4 output316 (.A(\Inst_LUT4AB_switch_matrix.S4BEG1 ),
    .X(S4BEG[13]));
 sky130_fd_sc_hd__buf_2 output317 (.A(net317),
    .X(S4BEG[14]));
 sky130_fd_sc_hd__buf_2 output318 (.A(net318),
    .X(S4BEG[15]));
 sky130_fd_sc_hd__buf_2 output319 (.A(net319),
    .X(S4BEG[1]));
 sky130_fd_sc_hd__buf_2 output320 (.A(net320),
    .X(S4BEG[2]));
 sky130_fd_sc_hd__buf_2 output321 (.A(net321),
    .X(S4BEG[3]));
 sky130_fd_sc_hd__buf_2 output322 (.A(net322),
    .X(S4BEG[4]));
 sky130_fd_sc_hd__buf_2 output323 (.A(net323),
    .X(S4BEG[5]));
 sky130_fd_sc_hd__buf_2 output324 (.A(net324),
    .X(S4BEG[6]));
 sky130_fd_sc_hd__buf_2 output325 (.A(net325),
    .X(S4BEG[7]));
 sky130_fd_sc_hd__buf_2 output326 (.A(net326),
    .X(S4BEG[8]));
 sky130_fd_sc_hd__buf_2 output327 (.A(net327),
    .X(S4BEG[9]));
 sky130_fd_sc_hd__buf_2 output328 (.A(net328),
    .X(SS4BEG[0]));
 sky130_fd_sc_hd__buf_2 output329 (.A(net329),
    .X(SS4BEG[10]));
 sky130_fd_sc_hd__buf_2 output330 (.A(net330),
    .X(SS4BEG[11]));
 sky130_fd_sc_hd__buf_2 output331 (.A(net331),
    .X(SS4BEG[12]));
 sky130_fd_sc_hd__buf_6 output332 (.A(\Inst_LUT4AB_switch_matrix.SS4BEG1 ),
    .X(SS4BEG[13]));
 sky130_fd_sc_hd__buf_8 output333 (.A(\Inst_LUT4AB_switch_matrix.SS4BEG2 ),
    .X(SS4BEG[14]));
 sky130_fd_sc_hd__buf_6 output334 (.A(net334),
    .X(SS4BEG[15]));
 sky130_fd_sc_hd__buf_2 output335 (.A(net335),
    .X(SS4BEG[1]));
 sky130_fd_sc_hd__buf_2 output336 (.A(net336),
    .X(SS4BEG[2]));
 sky130_fd_sc_hd__buf_2 output337 (.A(net337),
    .X(SS4BEG[3]));
 sky130_fd_sc_hd__buf_2 output338 (.A(net338),
    .X(SS4BEG[4]));
 sky130_fd_sc_hd__buf_2 output339 (.A(net339),
    .X(SS4BEG[5]));
 sky130_fd_sc_hd__buf_2 output340 (.A(net340),
    .X(SS4BEG[6]));
 sky130_fd_sc_hd__buf_2 output341 (.A(net341),
    .X(SS4BEG[7]));
 sky130_fd_sc_hd__buf_2 output342 (.A(net342),
    .X(SS4BEG[8]));
 sky130_fd_sc_hd__buf_2 output343 (.A(net343),
    .X(SS4BEG[9]));
 sky130_fd_sc_hd__buf_1 output344 (.A(net344),
    .X(UserCLKo));
 sky130_fd_sc_hd__clkbuf_4 output345 (.A(net345),
    .X(W1BEG[0]));
 sky130_fd_sc_hd__buf_8 output346 (.A(\Inst_LUT4AB_switch_matrix.W1BEG1 ),
    .X(W1BEG[1]));
 sky130_fd_sc_hd__buf_6 output347 (.A(\Inst_LUT4AB_switch_matrix.W1BEG2 ),
    .X(W1BEG[2]));
 sky130_fd_sc_hd__buf_8 output348 (.A(\Inst_LUT4AB_switch_matrix.W1BEG3 ),
    .X(W1BEG[3]));
 sky130_fd_sc_hd__buf_4 output349 (.A(net349),
    .X(W2BEG[0]));
 sky130_fd_sc_hd__buf_6 output350 (.A(net350),
    .X(W2BEG[1]));
 sky130_fd_sc_hd__buf_8 output351 (.A(net351),
    .X(W2BEG[2]));
 sky130_fd_sc_hd__buf_6 output352 (.A(net352),
    .X(W2BEG[3]));
 sky130_fd_sc_hd__buf_8 output353 (.A(net353),
    .X(W2BEG[4]));
 sky130_fd_sc_hd__buf_6 output354 (.A(net429),
    .X(W2BEG[5]));
 sky130_fd_sc_hd__buf_6 output355 (.A(net355),
    .X(W2BEG[6]));
 sky130_fd_sc_hd__buf_6 output356 (.A(\Inst_LUT4AB_switch_matrix.JW2BEG7 ),
    .X(W2BEG[7]));
 sky130_fd_sc_hd__buf_2 output357 (.A(net357),
    .X(W2BEGb[0]));
 sky130_fd_sc_hd__buf_2 output358 (.A(net358),
    .X(W2BEGb[1]));
 sky130_fd_sc_hd__buf_2 output359 (.A(net359),
    .X(W2BEGb[2]));
 sky130_fd_sc_hd__buf_2 output360 (.A(net360),
    .X(W2BEGb[3]));
 sky130_fd_sc_hd__buf_2 output361 (.A(net361),
    .X(W2BEGb[4]));
 sky130_fd_sc_hd__buf_2 output362 (.A(net362),
    .X(W2BEGb[5]));
 sky130_fd_sc_hd__buf_2 output363 (.A(net363),
    .X(W2BEGb[6]));
 sky130_fd_sc_hd__buf_2 output364 (.A(net364),
    .X(W2BEGb[7]));
 sky130_fd_sc_hd__buf_2 output365 (.A(net365),
    .X(W6BEG[0]));
 sky130_fd_sc_hd__buf_8 output366 (.A(\Inst_LUT4AB_switch_matrix.W6BEG0 ),
    .X(W6BEG[10]));
 sky130_fd_sc_hd__buf_6 output367 (.A(\Inst_LUT4AB_switch_matrix.W6BEG1 ),
    .X(W6BEG[11]));
 sky130_fd_sc_hd__buf_2 output368 (.A(net368),
    .X(W6BEG[1]));
 sky130_fd_sc_hd__buf_2 output369 (.A(net369),
    .X(W6BEG[2]));
 sky130_fd_sc_hd__buf_2 output370 (.A(net370),
    .X(W6BEG[3]));
 sky130_fd_sc_hd__buf_2 output371 (.A(net371),
    .X(W6BEG[4]));
 sky130_fd_sc_hd__buf_2 output372 (.A(net372),
    .X(W6BEG[5]));
 sky130_fd_sc_hd__buf_2 output373 (.A(net373),
    .X(W6BEG[6]));
 sky130_fd_sc_hd__buf_2 output374 (.A(net374),
    .X(W6BEG[7]));
 sky130_fd_sc_hd__buf_2 output375 (.A(net375),
    .X(W6BEG[8]));
 sky130_fd_sc_hd__buf_2 output376 (.A(net376),
    .X(W6BEG[9]));
 sky130_fd_sc_hd__buf_2 output377 (.A(net377),
    .X(WW4BEG[0]));
 sky130_fd_sc_hd__buf_2 output378 (.A(net378),
    .X(WW4BEG[10]));
 sky130_fd_sc_hd__buf_2 output379 (.A(net379),
    .X(WW4BEG[11]));
 sky130_fd_sc_hd__buf_4 output380 (.A(net380),
    .X(WW4BEG[12]));
 sky130_fd_sc_hd__buf_8 output381 (.A(\Inst_LUT4AB_switch_matrix.WW4BEG1 ),
    .X(WW4BEG[13]));
 sky130_fd_sc_hd__buf_2 output382 (.A(net382),
    .X(WW4BEG[14]));
 sky130_fd_sc_hd__buf_8 output383 (.A(\Inst_LUT4AB_switch_matrix.WW4BEG3 ),
    .X(WW4BEG[15]));
 sky130_fd_sc_hd__buf_2 output384 (.A(net384),
    .X(WW4BEG[1]));
 sky130_fd_sc_hd__buf_2 output385 (.A(net385),
    .X(WW4BEG[2]));
 sky130_fd_sc_hd__buf_2 output386 (.A(net386),
    .X(WW4BEG[3]));
 sky130_fd_sc_hd__buf_2 output387 (.A(net387),
    .X(WW4BEG[4]));
 sky130_fd_sc_hd__buf_2 output388 (.A(net388),
    .X(WW4BEG[5]));
 sky130_fd_sc_hd__buf_2 output389 (.A(net389),
    .X(WW4BEG[6]));
 sky130_fd_sc_hd__buf_2 output390 (.A(net390),
    .X(WW4BEG[7]));
 sky130_fd_sc_hd__buf_2 output391 (.A(net391),
    .X(WW4BEG[8]));
 sky130_fd_sc_hd__buf_2 output392 (.A(net392),
    .X(WW4BEG[9]));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_regs_0_UserCLK (.A(UserCLK),
    .X(UserCLK_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_UserCLK (.A(UserCLK),
    .X(clknet_0_UserCLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_UserCLK (.A(clknet_0_UserCLK),
    .X(clknet_1_0__leaf_UserCLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_UserCLK_regs (.A(UserCLK_regs),
    .X(clknet_0_UserCLK_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_UserCLK_regs (.A(clknet_0_UserCLK_regs),
    .X(clknet_1_0__leaf_UserCLK_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_UserCLK_regs (.A(clknet_0_UserCLK_regs),
    .X(clknet_1_1__leaf_UserCLK_regs));
 sky130_fd_sc_hd__buf_6 rebuffer4 (.A(_0327_),
    .X(net396));
 sky130_fd_sc_hd__mux2_4 clone5 (.A0(net409),
    .A1(net401),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit16.Q ),
    .X(net397));
 sky130_fd_sc_hd__mux2_4 clone6 (.A0(net417),
    .A1(_0396_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit17.Q ),
    .X(net398));
 sky130_fd_sc_hd__clkbuf_2 rebuffer8 (.A(\Inst_LUT4AB_switch_matrix.JS2BEG7 ),
    .X(net400));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer9 (.A(_0355_),
    .X(net401));
 sky130_fd_sc_hd__buf_6 rebuffer10 (.A(\Inst_LUT4AB_switch_matrix.M_AD ),
    .X(net402));
 sky130_fd_sc_hd__buf_6 rebuffer11 (.A(net402),
    .X(net403));
 sky130_fd_sc_hd__buf_6 rebuffer12 (.A(net425),
    .X(net404));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer13 (.A(net404),
    .X(net405));
 sky130_fd_sc_hd__buf_6 rebuffer14 (.A(net446),
    .X(net406));
 sky130_fd_sc_hd__buf_6 rebuffer15 (.A(_0327_),
    .X(net407));
 sky130_fd_sc_hd__clkbuf_2 rebuffer16 (.A(\Inst_LUT4AB_switch_matrix.JS2BEG5 ),
    .X(net408));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer17 (.A(_0354_),
    .X(net409));
 sky130_fd_sc_hd__buf_6 clone18 (.A(H),
    .X(net410));
 sky130_fd_sc_hd__clkbuf_1 clone19 (.A(D),
    .X(net411));
 sky130_fd_sc_hd__buf_6 rebuffer20 (.A(net428),
    .X(net412));
 sky130_fd_sc_hd__clkbuf_1 clone21 (.A(G),
    .X(net413));
 sky130_fd_sc_hd__buf_6 rebuffer22 (.A(\Inst_LUT4AB_switch_matrix.M_AH ),
    .X(net414));
 sky130_fd_sc_hd__buf_6 rebuffer23 (.A(net414),
    .X(net415));
 sky130_fd_sc_hd__buf_6 rebuffer24 (.A(\Inst_LUT4AB_switch_matrix.M_AH ),
    .X(net416));
 sky130_fd_sc_hd__buf_6 rebuffer25 (.A(_0395_),
    .X(net417));
 sky130_fd_sc_hd__clkbuf_2 rebuffer33 (.A(\Inst_LUT4AB_switch_matrix.M_AD ),
    .X(net425));
 sky130_fd_sc_hd__buf_8 clone34 (.A(net663),
    .X(net426));
 sky130_fd_sc_hd__buf_6 rebuffer35 (.A(net433),
    .X(net427));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer36 (.A(_0352_),
    .X(net428));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer37 (.A(\Inst_LUT4AB_switch_matrix.JW2BEG5 ),
    .X(net429));
 sky130_fd_sc_hd__clkbuf_1 clone38 (.A(net655),
    .X(net430));
 sky130_fd_sc_hd__dlymetal6s2s_1 clone40 (.A(\Inst_LUT4AB_switch_matrix.M_EF ),
    .X(net432));
 sky130_fd_sc_hd__buf_6 rebuffer60 (.A(net453),
    .X(net452));
 sky130_fd_sc_hd__buf_6 rebuffer61 (.A(net454),
    .X(net453));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer62 (.A(net398),
    .X(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(EE4END[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(EE4END[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(EE4END[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(EE4END[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(EE4END[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(EE4END[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(EE4END[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(EE4END[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(EE4END[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(EE4END[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(FrameStrobe[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(FrameStrobe[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(FrameStrobe[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(FrameStrobe[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(\Inst_LUT4AB_switch_matrix.JW2BEG6 ));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(N4END[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(N4END[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(N4END[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(N4END[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_41 (.DIODE(N4END[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_42 (.DIODE(N4END[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_43 (.DIODE(N4END[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_44 (.DIODE(N4END[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_45 (.DIODE(N4END[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_46 (.DIODE(N4END[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_47 (.DIODE(N4END[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_48 (.DIODE(NN4END[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_49 (.DIODE(NN4END[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_50 (.DIODE(NN4END[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_51 (.DIODE(NN4END[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_52 (.DIODE(NN4END[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_53 (.DIODE(NN4END[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_54 (.DIODE(NN4END[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_55 (.DIODE(NN4END[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_56 (.DIODE(NN4END[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_57 (.DIODE(NN4END[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_58 (.DIODE(NN4END[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_59 (.DIODE(NN4END[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_60 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_61 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA_62 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_63 (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA_64 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_65 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_66 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA_67 (.DIODE(S4END[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_68 (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA_69 (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA_70 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA_71 (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA_72 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA_73 (.DIODE(W6END[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_74 (.DIODE(_0053_));
 sky130_fd_sc_hd__diode_2 ANTENNA_75 (.DIODE(_0053_));
 sky130_fd_sc_hd__diode_2 ANTENNA_76 (.DIODE(_0053_));
 sky130_fd_sc_hd__diode_2 ANTENNA_77 (.DIODE(_0053_));
 sky130_fd_sc_hd__diode_2 ANTENNA_78 (.DIODE(_0063_));
 sky130_fd_sc_hd__diode_2 ANTENNA_79 (.DIODE(_0063_));
 sky130_fd_sc_hd__diode_2 ANTENNA_80 (.DIODE(_0063_));
 sky130_fd_sc_hd__diode_2 ANTENNA_81 (.DIODE(_0120_));
 sky130_fd_sc_hd__diode_2 ANTENNA_82 (.DIODE(_0120_));
 sky130_fd_sc_hd__diode_2 ANTENNA_83 (.DIODE(_0120_));
 sky130_fd_sc_hd__diode_2 ANTENNA_84 (.DIODE(_0120_));
 sky130_fd_sc_hd__diode_2 ANTENNA_85 (.DIODE(_0120_));
 sky130_fd_sc_hd__diode_2 ANTENNA_86 (.DIODE(_0662_));
 sky130_fd_sc_hd__diode_2 ANTENNA_87 (.DIODE(_0662_));
 sky130_fd_sc_hd__diode_2 ANTENNA_88 (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA_89 (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA_90 (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_91 (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_92 (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_93 (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_94 (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_95 (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_96 (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_97 (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA_98 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_99 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_100 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_101 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_102 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_103 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_104 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA_105 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_106 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_107 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_108 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_109 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_110 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_111 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_112 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_113 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_114 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_115 (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA_116 (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA_117 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA_118 (.DIODE(EE4END[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_119 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA_120 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_121 (.DIODE(FrameStrobe[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_122 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_123 (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA_124 (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA_125 (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA_126 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA_127 (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_128 (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA_129 (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_130 (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_131 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_132 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_133 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_134 (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_135 (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA_136 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_137 (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_138 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_139 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_140 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_141 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_142 (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA_143 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_144 (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA_145 (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA_146 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA_147 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_148 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_149 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_150 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_151 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_152 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_153 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_154 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_155 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_156 (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_157 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_158 (.DIODE(net147));
 sky130_fd_sc_hd__fill_1 FILLER_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_255 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_107 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_367 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_115 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_20 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_14 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_338 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_198 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_31 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_50 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_28 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_368 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_5 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_385 ();
endmodule
