* NGSPICE file created from S_WARMBOOT.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlxtp_1 abstract view
.subckt sky130_fd_sc_hd__dlxtp_1 D GATE VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_1 abstract view
.subckt sky130_fd_sc_hd__inv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

.subckt S_WARMBOOT BOOT_top Co FrameData[0] FrameData[10] FrameData[11] FrameData[12]
+ FrameData[13] FrameData[14] FrameData[15] FrameData[16] FrameData[17] FrameData[18]
+ FrameData[19] FrameData[1] FrameData[20] FrameData[21] FrameData[22] FrameData[23]
+ FrameData[24] FrameData[25] FrameData[26] FrameData[27] FrameData[28] FrameData[29]
+ FrameData[2] FrameData[30] FrameData[31] FrameData[3] FrameData[4] FrameData[5]
+ FrameData[6] FrameData[7] FrameData[8] FrameData[9] FrameData_O[0] FrameData_O[10]
+ FrameData_O[11] FrameData_O[12] FrameData_O[13] FrameData_O[14] FrameData_O[15]
+ FrameData_O[16] FrameData_O[17] FrameData_O[18] FrameData_O[19] FrameData_O[1] FrameData_O[20]
+ FrameData_O[21] FrameData_O[22] FrameData_O[23] FrameData_O[24] FrameData_O[25]
+ FrameData_O[26] FrameData_O[27] FrameData_O[28] FrameData_O[29] FrameData_O[2] FrameData_O[30]
+ FrameData_O[31] FrameData_O[3] FrameData_O[4] FrameData_O[5] FrameData_O[6] FrameData_O[7]
+ FrameData_O[8] FrameData_O[9] FrameStrobe[0] FrameStrobe[10] FrameStrobe[11] FrameStrobe[12]
+ FrameStrobe[13] FrameStrobe[14] FrameStrobe[15] FrameStrobe[16] FrameStrobe[17]
+ FrameStrobe[18] FrameStrobe[19] FrameStrobe[1] FrameStrobe[2] FrameStrobe[3] FrameStrobe[4]
+ FrameStrobe[5] FrameStrobe[6] FrameStrobe[7] FrameStrobe[8] FrameStrobe[9] FrameStrobe_O[0]
+ FrameStrobe_O[10] FrameStrobe_O[11] FrameStrobe_O[12] FrameStrobe_O[13] FrameStrobe_O[14]
+ FrameStrobe_O[15] FrameStrobe_O[16] FrameStrobe_O[17] FrameStrobe_O[18] FrameStrobe_O[19]
+ FrameStrobe_O[1] FrameStrobe_O[2] FrameStrobe_O[3] FrameStrobe_O[4] FrameStrobe_O[5]
+ FrameStrobe_O[6] FrameStrobe_O[7] FrameStrobe_O[8] FrameStrobe_O[9] N1BEG[0] N1BEG[1]
+ N1BEG[2] N1BEG[3] N2BEG[0] N2BEG[1] N2BEG[2] N2BEG[3] N2BEG[4] N2BEG[5] N2BEG[6]
+ N2BEG[7] N2BEGb[0] N2BEGb[1] N2BEGb[2] N2BEGb[3] N2BEGb[4] N2BEGb[5] N2BEGb[6] N2BEGb[7]
+ N4BEG[0] N4BEG[10] N4BEG[11] N4BEG[12] N4BEG[13] N4BEG[14] N4BEG[15] N4BEG[1] N4BEG[2]
+ N4BEG[3] N4BEG[4] N4BEG[5] N4BEG[6] N4BEG[7] N4BEG[8] N4BEG[9] NN4BEG[0] NN4BEG[10]
+ NN4BEG[11] NN4BEG[12] NN4BEG[13] NN4BEG[14] NN4BEG[15] NN4BEG[1] NN4BEG[2] NN4BEG[3]
+ NN4BEG[4] NN4BEG[5] NN4BEG[6] NN4BEG[7] NN4BEG[8] NN4BEG[9] RESET_top S1END[0] S1END[1]
+ S1END[2] S1END[3] S2END[0] S2END[1] S2END[2] S2END[3] S2END[4] S2END[5] S2END[6]
+ S2END[7] S2MID[0] S2MID[1] S2MID[2] S2MID[3] S2MID[4] S2MID[5] S2MID[6] S2MID[7]
+ S4END[0] S4END[10] S4END[11] S4END[12] S4END[13] S4END[14] S4END[15] S4END[1] S4END[2]
+ S4END[3] S4END[4] S4END[5] S4END[6] S4END[7] S4END[8] S4END[9] SLOT_top0 SLOT_top1
+ SLOT_top2 SLOT_top3 SS4END[0] SS4END[10] SS4END[11] SS4END[12] SS4END[13] SS4END[14]
+ SS4END[15] SS4END[1] SS4END[2] SS4END[3] SS4END[4] SS4END[5] SS4END[6] SS4END[7]
+ SS4END[8] SS4END[9] UserCLK UserCLKo VGND VPWR
XFILLER_9_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_0_Left_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_11_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_131_ FrameStrobe[10] VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__clkbuf_1
X_062_ net31 net35 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit17.Q VGND VGND VPWR VPWR
+ _028_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_045_ _011_ _012_ _013_ Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit27.Q Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit28.Q
+ VGND VGND VPWR VPWR _014_ sky130_fd_sc_hd__a221o_1
XFILLER_7_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_114_ net15 VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_5_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout7 net8 VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_2
XANTENNA_5 FrameData[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_319 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput97 net99 VGND VGND VPWR VPWR FrameStrobe_O[19] sky130_fd_sc_hd__buf_2
Xoutput75 net77 VGND VGND VPWR VPWR FrameData_O[28] sky130_fd_sc_hd__buf_2
Xoutput64 net66 VGND VGND VPWR VPWR FrameData_O[18] sky130_fd_sc_hd__buf_2
XFILLER_8_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput86 net88 VGND VGND VPWR VPWR FrameData_O[9] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_2_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_355 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_130_ FrameStrobe[9] VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__clkbuf_1
XFILLER_9_12 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_061_ net27 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit17.Q Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit18.Q
+ VGND VGND VPWR VPWR _027_ sky130_fd_sc_hd__o21ba_1
X_044_ net30 net34 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit26.Q VGND VGND VPWR VPWR
+ _013_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_5_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_113_ net14 VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__buf_1
XFILLER_6_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout8 net22 VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__buf_2
XANTENNA_6 FrameData[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput98 net100 VGND VGND VPWR VPWR FrameStrobe_O[1] sky130_fd_sc_hd__buf_2
Xoutput87 net89 VGND VGND VPWR VPWR FrameStrobe_O[0] sky130_fd_sc_hd__buf_2
Xoutput76 net78 VGND VGND VPWR VPWR FrameData_O[29] sky130_fd_sc_hd__buf_2
Xoutput65 net67 VGND VGND VPWR VPWR FrameData_O[19] sky130_fd_sc_hd__buf_2
XFILLER_0_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput54 net56 VGND VGND VPWR VPWR BOOT_top sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_2_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_367 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_24 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_060_ net39 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit17.Q VGND VGND VPWR VPWR _026_
+ sky130_fd_sc_hd__nand2b_1
XFILLER_9_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_189_ net51 VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__buf_1
XFILLER_11_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_043_ net26 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit26.Q Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit27.Q
+ VGND VGND VPWR VPWR _012_ sky130_fd_sc_hd__o21ba_1
X_112_ net13 VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_5_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_7 net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput88 net90 VGND VGND VPWR VPWR FrameStrobe_O[10] sky130_fd_sc_hd__buf_2
Xoutput99 net101 VGND VGND VPWR VPWR FrameStrobe_O[2] sky130_fd_sc_hd__buf_2
XFILLER_0_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput77 net79 VGND VGND VPWR VPWR FrameData_O[2] sky130_fd_sc_hd__buf_2
Xoutput66 net68 VGND VGND VPWR VPWR FrameData_O[1] sky130_fd_sc_hd__buf_2
Xoutput55 net57 VGND VGND VPWR VPWR FrameData_O[0] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_2_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_379 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_11_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_4_Left_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_36 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_188_ net52 VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__clkbuf_1
XFILLER_11_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_042_ net38 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit26.Q VGND VGND VPWR VPWR _011_
+ sky130_fd_sc_hd__nand2b_1
X_111_ net12 VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__clkbuf_1
XFILLER_1_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_8 FrameStrobe[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput89 net91 VGND VGND VPWR VPWR FrameStrobe_O[11] sky130_fd_sc_hd__buf_2
Xoutput67 net69 VGND VGND VPWR VPWR FrameData_O[20] sky130_fd_sc_hd__buf_2
Xoutput78 net80 VGND VGND VPWR VPWR FrameData_O[30] sky130_fd_sc_hd__buf_2
XFILLER_0_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput56 net58 VGND VGND VPWR VPWR FrameData_O[10] sky130_fd_sc_hd__buf_2
XFILLER_8_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_187_ net53 VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__buf_1
XFILLER_11_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_041_ net42 net46 net50 net54 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit26.Q Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit27.Q
+ VGND VGND VPWR VPWR _010_ sky130_fd_sc_hd__mux4_1
X_110_ net11 VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__buf_1
XFILLER_1_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_9 FrameStrobe[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput57 net59 VGND VGND VPWR VPWR FrameData_O[11] sky130_fd_sc_hd__buf_2
Xoutput79 net81 VGND VGND VPWR VPWR FrameData_O[31] sky130_fd_sc_hd__buf_2
XFILLER_8_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput68 net70 VGND VGND VPWR VPWR FrameData_O[21] sky130_fd_sc_hd__buf_2
XFILLER_5_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_186_ net54 VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_040_ _000_ _005_ _009_ VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__o21a_1
XFILLER_1_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_169_ net47 VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__clkbuf_1
XFILLER_10_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput69 net71 VGND VGND VPWR VPWR FrameData_O[22] sky130_fd_sc_hd__buf_2
XFILLER_8_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput58 net60 VGND VGND VPWR VPWR FrameData_O[12] sky130_fd_sc_hd__buf_2
XS_WARMBOOT_164 VGND VGND VPWR VPWR S_WARMBOOT_164/HI Co sky130_fd_sc_hd__conb_1
XFILLER_5_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_11_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_185_ net55 VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__buf_1
XFILLER_9_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_099_ FrameData[10] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__clkbuf_2
X_168_ S4END[8] VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__clkbuf_1
XFILLER_6_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput59 net61 VGND VGND VPWR VPWR FrameData_O[13] sky130_fd_sc_hd__buf_2
XFILLER_0_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_342 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_9_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_184_ SS4END[8] VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__buf_1
X_167_ S4END[9] VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__buf_1
X_098_ FrameData[9] VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__buf_1
XFILLER_10_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_11_Left_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_62 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_3_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_340 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_183_ SS4END[9] VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__buf_1
XFILLER_10_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_097_ FrameData[8] VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__buf_1
XFILLER_6_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_166_ S4END[10] VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_6_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_149_ net39 VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_371 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_74 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_182_ SS4END[10] VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_9_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_207 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_165_ S4END[11] VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__buf_1
X_096_ FrameData[7] VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__clkbuf_1
XFILLER_6_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_148_ S2MID[4] VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_6_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_079_ net13 net8 VGND VGND VPWR VPWR Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_7_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_31 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_367 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_181_ SS4END[11] VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_0_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_095_ FrameData[6] VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__clkbuf_2
X_164_ S4END[12] VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__clkbuf_2
XFILLER_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_6_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_147_ S2MID[5] VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__clkbuf_1
X_078_ net12 net8 VGND VGND VPWR VPWR Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_8_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_180_ SS4END[12] VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_9_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_3_Left_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_094_ FrameData[5] VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__clkbuf_2
X_163_ S4END[13] VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__buf_1
XFILLER_10_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_146_ S2MID[6] VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_6_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_077_ net11 net8 VGND VGND VPWR VPWR Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_7_99 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_129_ FrameStrobe[8] VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__clkbuf_1
XFILLER_8_127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_093_ FrameData[4] VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__clkbuf_2
X_162_ S4END[14] VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__clkbuf_2
XFILLER_1_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput1 FrameData[13] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__buf_1
X_145_ S2MID[7] VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_6_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_076_ net10 net8 VGND VGND VPWR VPWR Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_059_ net43 net47 net51 net55 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit17.Q Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit18.Q
+ VGND VGND VPWR VPWR _025_ sky130_fd_sc_hd__mux4_1
X_128_ FrameStrobe[7] VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__clkbuf_1
XFILLER_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_161_ S4END[15] VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__clkbuf_1
X_092_ FrameData[3] VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__clkbuf_1
XFILLER_1_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput2 FrameData[14] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__buf_1
XFILLER_5_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_207 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_075_ net9 net8 VGND VGND VPWR VPWR Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_6_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_144_ Inst_S_WARMBOOT_switch_matrix.N1BEG3 VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__buf_1
XFILLER_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_058_ _003_ _020_ _024_ VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__o21a_1
X_127_ FrameStrobe[6] VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_3_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_091_ FrameData[2] VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_160_ net28 VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__buf_1
XFILLER_1_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_7_Left_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput3 FrameData[15] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__buf_1
XFILLER_5_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_143_ Inst_S_WARMBOOT_switch_matrix.N1BEG2 VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__buf_1
X_074_ net6 net8 VGND VGND VPWR VPWR Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_3_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_057_ _021_ _022_ _023_ Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit21.Q Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit22.Q
+ VGND VGND VPWR VPWR _024_ sky130_fd_sc_hd__a221o_1
X_126_ FrameStrobe[5] VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__clkbuf_1
Xinput50 SS4END[4] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_109_ net10 VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_10_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_122 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_090_ FrameData[1] VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__clkbuf_1
XFILLER_10_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput4 FrameData[16] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__buf_1
XFILLER_5_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_142_ Inst_S_WARMBOOT_switch_matrix.N1BEG1 VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__buf_1
XFILLER_2_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_073_ net5 net8 VGND VGND VPWR VPWR Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
X_056_ net28 net32 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit20.Q VGND VGND VPWR VPWR
+ _023_ sky130_fd_sc_hd__mux2_1
Xoutput160 net162 VGND VGND VPWR VPWR SLOT_top1 sky130_fd_sc_hd__buf_2
X_125_ FrameStrobe[4] VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__clkbuf_1
Xinput51 SS4END[5] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__clkbuf_1
Xinput40 S4END[2] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_10_Left_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_7_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_108_ net9 VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_039_ _006_ _007_ _008_ Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit30.Q Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit31.Q
+ VGND VGND VPWR VPWR _009_ sky130_fd_sc_hd__a221o_1
XFILLER_8_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_10_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput5 FrameData[17] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__buf_1
XFILLER_5_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_072_ net4 net7 VGND VGND VPWR VPWR Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
X_141_ Inst_S_WARMBOOT_switch_matrix.N1BEG0 VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__buf_1
XANTENNA_10 FrameStrobe[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput150 net152 VGND VGND VPWR VPWR NN4BEG[1] sky130_fd_sc_hd__buf_2
XFILLER_7_324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_124_ FrameStrobe[3] VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__clkbuf_1
Xoutput161 net163 VGND VGND VPWR VPWR SLOT_top2 sky130_fd_sc_hd__buf_2
X_055_ net24 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit20.Q Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit21.Q
+ VGND VGND VPWR VPWR _022_ sky130_fd_sc_hd__o21ba_1
Xinput41 S4END[3] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__buf_1
Xinput30 S2END[4] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__buf_1
Xinput52 SS4END[6] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_7_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_316 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_107_ net6 VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__clkbuf_2
X_038_ net31 net35 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit29.Q VGND VGND VPWR VPWR
+ _008_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_10_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput6 FrameData[18] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_1
X_140_ FrameStrobe[19] VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__clkbuf_1
X_071_ net3 net7 VGND VGND VPWR VPWR Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_2_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput151 net153 VGND VGND VPWR VPWR NN4BEG[2] sky130_fd_sc_hd__buf_2
Xoutput140 net142 VGND VGND VPWR VPWR N4BEG[7] sky130_fd_sc_hd__buf_2
Xoutput162 net164 VGND VGND VPWR VPWR SLOT_top3 sky130_fd_sc_hd__buf_2
XANTENNA_11 net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput31 S2END[5] VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__buf_1
X_123_ FrameStrobe[2] VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_7_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_054_ net36 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit20.Q VGND VGND VPWR VPWR _021_
+ sky130_fd_sc_hd__nand2b_1
Xinput20 FrameStrobe[0] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__buf_1
Xinput53 SS4END[7] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__clkbuf_2
Xinput42 S4END[4] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__clkbuf_1
XFILLER_4_328 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_037_ net27 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit29.Q Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit30.Q
+ VGND VGND VPWR VPWR _007_ sky130_fd_sc_hd__o21ba_1
X_106_ net5 VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput7 FrameData[19] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_1_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_070_ net2 net7 VGND VGND VPWR VPWR Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_2_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput163 net165 VGND VGND VPWR VPWR UserCLKo sky130_fd_sc_hd__buf_1
Xoutput152 net154 VGND VGND VPWR VPWR NN4BEG[3] sky130_fd_sc_hd__buf_2
Xoutput130 net132 VGND VGND VPWR VPWR N4BEG[12] sky130_fd_sc_hd__buf_2
Xoutput141 net143 VGND VGND VPWR VPWR N4BEG[8] sky130_fd_sc_hd__buf_2
XANTENNA_12 net51 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_359 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_122_ FrameStrobe[1] VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__clkbuf_1
X_053_ net40 net44 net48 net52 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit20.Q Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit21.Q
+ VGND VGND VPWR VPWR _020_ sky130_fd_sc_hd__mux4_1
Xinput43 S4END[5] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__buf_1
Xinput32 S2END[6] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__clkbuf_1
Xinput10 FrameData[22] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__buf_1
Xinput21 RESET_top VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_11_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_105_ net4 VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__clkbuf_1
XFILLER_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_036_ net39 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit29.Q VGND VGND VPWR VPWR _006_
+ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_10_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput8 FrameData[20] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_1_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_2_Left_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput131 net133 VGND VGND VPWR VPWR N4BEG[13] sky130_fd_sc_hd__buf_2
Xoutput120 net122 VGND VGND VPWR VPWR N2BEGb[1] sky130_fd_sc_hd__buf_2
XANTENNA_13 net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput153 net155 VGND VGND VPWR VPWR NN4BEG[4] sky130_fd_sc_hd__buf_2
Xoutput142 net144 VGND VGND VPWR VPWR N4BEG[9] sky130_fd_sc_hd__buf_2
XFILLER_2_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_52 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_323 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_052_ _002_ _015_ _019_ VGND VGND VPWR VPWR net162 sky130_fd_sc_hd__o21a_1
XFILLER_7_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_121_ net8 VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__buf_1
Xinput44 S4END[6] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__clkbuf_1
Xinput33 S2END[7] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__buf_1
Xinput11 FrameData[23] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__buf_1
Xinput22 S1END[0] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__buf_1
XFILLER_6_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_7_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_104_ net3 VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__buf_1
XFILLER_7_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_035_ net43 net47 net51 net55 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit29.Q Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit30.Q
+ VGND VGND VPWR VPWR _005_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_10_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_274 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput9 FrameData[21] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__buf_1
XFILLER_5_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput143 net145 VGND VGND VPWR VPWR NN4BEG[0] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput132 net134 VGND VGND VPWR VPWR N4BEG[14] sky130_fd_sc_hd__buf_2
Xoutput121 net123 VGND VGND VPWR VPWR N2BEGb[2] sky130_fd_sc_hd__buf_2
Xoutput110 net112 VGND VGND VPWR VPWR N1BEG[3] sky130_fd_sc_hd__buf_2
XFILLER_9_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_64 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput154 net156 VGND VGND VPWR VPWR NN4BEG[5] sky130_fd_sc_hd__buf_2
X_120_ net21 VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__clkbuf_2
X_051_ _016_ _017_ _018_ Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit24.Q Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit25.Q
+ VGND VGND VPWR VPWR _019_ sky130_fd_sc_hd__a221o_1
Xinput45 S4END[7] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__buf_1
Xinput34 S2MID[0] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__buf_1
Xinput12 FrameData[24] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput23 S1END[1] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_7_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_103_ net2 VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__buf_1
XFILLER_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_342 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_034_ Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit19.Q VGND VGND VPWR VPWR _004_ sky130_fd_sc_hd__inv_1
XFILLER_8_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_86 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput100 net102 VGND VGND VPWR VPWR FrameStrobe_O[3] sky130_fd_sc_hd__buf_2
Xoutput133 net135 VGND VGND VPWR VPWR N4BEG[15] sky130_fd_sc_hd__buf_2
Xoutput122 net124 VGND VGND VPWR VPWR N2BEGb[3] sky130_fd_sc_hd__buf_2
Xoutput111 net113 VGND VGND VPWR VPWR N2BEG[0] sky130_fd_sc_hd__buf_2
Xoutput144 net146 VGND VGND VPWR VPWR NN4BEG[10] sky130_fd_sc_hd__buf_2
Xoutput155 net157 VGND VGND VPWR VPWR NN4BEG[6] sky130_fd_sc_hd__buf_2
X_050_ net29 net33 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit23.Q VGND VGND VPWR VPWR
+ _018_ sky130_fd_sc_hd__mux2_1
Xinput46 SS4END[0] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__buf_1
Xinput35 S2MID[1] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__buf_1
Xinput24 S1END[2] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__clkbuf_1
XFILLER_11_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput13 FrameData[25] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__buf_1
XFILLER_10_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_7_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_179_ SS4END[13] VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__buf_1
XFILLER_7_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_033_ Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit22.Q VGND VGND VPWR VPWR _003_ sky130_fd_sc_hd__inv_2
XFILLER_3_354 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_102_ net1 VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__buf_1
XFILLER_8_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_107 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_195 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput101 net103 VGND VGND VPWR VPWR FrameStrobe_O[4] sky130_fd_sc_hd__buf_2
XFILLER_11_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput145 net147 VGND VGND VPWR VPWR NN4BEG[11] sky130_fd_sc_hd__buf_2
Xoutput156 net158 VGND VGND VPWR VPWR NN4BEG[7] sky130_fd_sc_hd__buf_2
Xoutput134 net136 VGND VGND VPWR VPWR N4BEG[1] sky130_fd_sc_hd__buf_2
Xoutput123 net125 VGND VGND VPWR VPWR N2BEGb[4] sky130_fd_sc_hd__buf_2
Xoutput112 net114 VGND VGND VPWR VPWR N2BEG[1] sky130_fd_sc_hd__buf_2
XFILLER_9_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_6_Left_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput36 S2MID[2] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__clkbuf_1
Xinput25 S1END[3] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__buf_1
Xinput14 FrameData[26] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__buf_1
Xinput47 SS4END[1] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__clkbuf_1
X_178_ SS4END[14] VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__buf_1
X_101_ FrameData[12] VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__clkbuf_1
X_032_ Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit25.Q VGND VGND VPWR VPWR _002_ sky130_fd_sc_hd__inv_2
XFILLER_3_366 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_9_Left_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_152 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput102 net104 VGND VGND VPWR VPWR FrameStrobe_O[5] sky130_fd_sc_hd__buf_2
Xoutput146 net148 VGND VGND VPWR VPWR NN4BEG[12] sky130_fd_sc_hd__buf_2
Xoutput157 net159 VGND VGND VPWR VPWR NN4BEG[8] sky130_fd_sc_hd__buf_2
Xoutput124 net126 VGND VGND VPWR VPWR N2BEGb[5] sky130_fd_sc_hd__buf_2
Xoutput113 net115 VGND VGND VPWR VPWR N2BEG[2] sky130_fd_sc_hd__buf_2
Xoutput135 net137 VGND VGND VPWR VPWR N4BEG[2] sky130_fd_sc_hd__buf_2
XFILLER_9_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput48 SS4END[2] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__buf_1
Xinput26 S2END[0] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__buf_1
Xinput37 S2MID[3] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__clkbuf_1
X_177_ SS4END[15] VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__buf_1
Xinput15 FrameData[27] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__clkbuf_1
XFILLER_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_100_ FrameData[11] VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__clkbuf_1
X_031_ Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit28.Q VGND VGND VPWR VPWR _001_ sky130_fd_sc_hd__inv_2
XFILLER_3_378 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_193_ UserCLK VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__buf_2
Xoutput103 net105 VGND VGND VPWR VPWR FrameStrobe_O[6] sky130_fd_sc_hd__buf_2
Xoutput158 net160 VGND VGND VPWR VPWR NN4BEG[9] sky130_fd_sc_hd__buf_2
Xoutput147 net149 VGND VGND VPWR VPWR NN4BEG[13] sky130_fd_sc_hd__buf_2
Xoutput136 net138 VGND VGND VPWR VPWR N4BEG[3] sky130_fd_sc_hd__buf_2
Xoutput125 net127 VGND VGND VPWR VPWR N2BEGb[6] sky130_fd_sc_hd__buf_2
Xoutput114 net116 VGND VGND VPWR VPWR N2BEG[3] sky130_fd_sc_hd__buf_2
XFILLER_9_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput49 SS4END[3] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput38 S4END[0] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__clkbuf_1
Xinput27 S2END[1] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__buf_1
XFILLER_10_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput16 FrameData[28] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__buf_1
XFILLER_6_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_176_ net40 VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__buf_1
XFILLER_9_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_12 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_030_ Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit31.Q VGND VGND VPWR VPWR _000_ sky130_fd_sc_hd__inv_1
X_159_ net29 VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__buf_1
XFILLER_0_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_192_ net48 VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__clkbuf_1
Xoutput148 net150 VGND VGND VPWR VPWR NN4BEG[14] sky130_fd_sc_hd__buf_2
Xoutput126 net128 VGND VGND VPWR VPWR N2BEGb[7] sky130_fd_sc_hd__buf_2
Xoutput115 net117 VGND VGND VPWR VPWR N2BEG[4] sky130_fd_sc_hd__buf_2
Xoutput104 net106 VGND VGND VPWR VPWR FrameStrobe_O[7] sky130_fd_sc_hd__buf_2
Xoutput137 net139 VGND VGND VPWR VPWR N4BEG[4] sky130_fd_sc_hd__buf_2
XFILLER_9_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput159 net161 VGND VGND VPWR VPWR SLOT_top0 sky130_fd_sc_hd__buf_2
XFILLER_2_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput39 S4END[1] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__buf_1
Xinput28 S2END[2] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__clkbuf_1
Xinput17 FrameData[29] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__buf_1
XFILLER_6_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_175_ net41 VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__buf_1
X_158_ net30 VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__buf_1
XFILLER_8_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_089_ FrameData[0] VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__clkbuf_2
XFILLER_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_272 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_191_ net49 VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__buf_1
Xoutput105 net107 VGND VGND VPWR VPWR FrameStrobe_O[8] sky130_fd_sc_hd__buf_2
Xoutput149 net151 VGND VGND VPWR VPWR NN4BEG[15] sky130_fd_sc_hd__buf_2
Xoutput138 net140 VGND VGND VPWR VPWR N4BEG[5] sky130_fd_sc_hd__buf_2
Xoutput116 net118 VGND VGND VPWR VPWR N2BEG[5] sky130_fd_sc_hd__buf_2
XFILLER_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput127 net129 VGND VGND VPWR VPWR N4BEG[0] sky130_fd_sc_hd__buf_2
XFILLER_9_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput29 S2END[3] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__buf_1
XFILLER_10_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput18 FrameData[30] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__buf_1
XFILLER_6_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_312 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_174_ net42 VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__buf_1
XFILLER_3_304 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_157_ net31 VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_8_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_190_ net50 VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__clkbuf_1
XFILLER_1_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput106 net108 VGND VGND VPWR VPWR FrameStrobe_O[9] sky130_fd_sc_hd__buf_2
Xoutput139 net141 VGND VGND VPWR VPWR N4BEG[6] sky130_fd_sc_hd__buf_2
Xoutput128 net130 VGND VGND VPWR VPWR N4BEG[10] sky130_fd_sc_hd__buf_2
Xoutput117 net119 VGND VGND VPWR VPWR N2BEG[6] sky130_fd_sc_hd__buf_2
XFILLER_10_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput19 FrameData[31] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__buf_1
XFILLER_6_324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_173_ net43 VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_1_Left_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_316 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_087_ net21 net7 VGND VGND VPWR VPWR Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_6_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_156_ net32 VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_8_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_139_ FrameStrobe[18] VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_5_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput118 net120 VGND VGND VPWR VPWR N2BEG[7] sky130_fd_sc_hd__buf_2
Xoutput129 net131 VGND VGND VPWR VPWR N4BEG[11] sky130_fd_sc_hd__buf_2
Xoutput107 net109 VGND VGND VPWR VPWR N1BEG[0] sky130_fd_sc_hd__buf_2
XFILLER_10_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_336 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_172_ net44 VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__buf_1
XFILLER_5_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_155_ net33 VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__buf_1
X_086_ net20 net7 VGND VGND VPWR VPWR Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_3_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_8_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_069_ net1 net7 VGND VGND VPWR VPWR Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
X_138_ FrameStrobe[17] VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput90 net92 VGND VGND VPWR VPWR FrameStrobe_O[12] sky130_fd_sc_hd__buf_2
Xoutput108 net110 VGND VGND VPWR VPWR N1BEG[1] sky130_fd_sc_hd__buf_2
Xoutput119 net121 VGND VGND VPWR VPWR N2BEGb[0] sky130_fd_sc_hd__buf_2
XFILLER_1_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_348 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_171_ net45 VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__buf_1
XFILLER_10_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_154_ net34 VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__buf_1
XFILLER_10_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_8_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_085_ net19 net7 VGND VGND VPWR VPWR Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_3_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_137_ FrameStrobe[16] VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__buf_1
X_068_ net27 net23 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit13.Q VGND VGND VPWR VPWR
+ Inst_S_WARMBOOT_switch_matrix.N1BEG0 sky130_fd_sc_hd__mux2_1
XFILLER_0_118 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_18 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput109 net111 VGND VGND VPWR VPWR N1BEG[2] sky130_fd_sc_hd__buf_2
XFILLER_9_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput91 net93 VGND VGND VPWR VPWR FrameStrobe_O[13] sky130_fd_sc_hd__buf_2
Xoutput80 net82 VGND VGND VPWR VPWR FrameData_O[3] sky130_fd_sc_hd__buf_2
XFILLER_10_312 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_170_ net46 VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__buf_1
XFILLER_5_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_5_Left_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_084_ net18 net7 VGND VGND VPWR VPWR Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_8_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_153_ net35 VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__clkbuf_1
XFILLER_7_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_136_ FrameStrobe[15] VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__buf_1
XFILLER_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_067_ net26 net23 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit14.Q VGND VGND VPWR VPWR
+ Inst_S_WARMBOOT_switch_matrix.N1BEG1 sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_8_Left_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_119_ net20 VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__buf_1
XFILLER_1_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput92 net94 VGND VGND VPWR VPWR FrameStrobe_O[14] sky130_fd_sc_hd__buf_2
XFILLER_11_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput70 net72 VGND VGND VPWR VPWR FrameData_O[23] sky130_fd_sc_hd__buf_2
Xoutput81 net83 VGND VGND VPWR VPWR FrameData_O[4] sky130_fd_sc_hd__buf_2
XFILLER_10_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_9_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_30 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_083_ net17 net7 VGND VGND VPWR VPWR Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_6_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_152_ net36 VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__buf_1
XFILLER_9_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_066_ net25 net23 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit15.Q VGND VGND VPWR VPWR
+ Inst_S_WARMBOOT_switch_matrix.N1BEG2 sky130_fd_sc_hd__mux2_1
X_135_ FrameStrobe[14] VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__clkbuf_1
XFILLER_8_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_049_ net25 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit23.Q Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit24.Q
+ VGND VGND VPWR VPWR _017_ sky130_fd_sc_hd__o21ba_1
XFILLER_7_231 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_118_ net19 VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__clkbuf_2
XFILLER_4_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_1 FrameData[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput71 net73 VGND VGND VPWR VPWR FrameData_O[24] sky130_fd_sc_hd__buf_2
Xoutput93 net95 VGND VGND VPWR VPWR FrameStrobe_O[15] sky130_fd_sc_hd__buf_2
XFILLER_9_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput82 net84 VGND VGND VPWR VPWR FrameData_O[5] sky130_fd_sc_hd__buf_2
Xoutput60 net62 VGND VGND VPWR VPWR FrameData_O[14] sky130_fd_sc_hd__buf_2
XFILLER_11_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_082_ net16 net7 VGND VGND VPWR VPWR Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
X_151_ net37 VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__buf_1
XFILLER_2_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_065_ net24 net23 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit16.Q VGND VGND VPWR VPWR
+ Inst_S_WARMBOOT_switch_matrix.N1BEG3 sky130_fd_sc_hd__mux2_1
X_134_ FrameStrobe[13] VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__clkbuf_1
X_117_ net18 VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__buf_1
XFILLER_7_243 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_048_ net37 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit23.Q VGND VGND VPWR VPWR _016_
+ sky130_fd_sc_hd__nand2b_1
XFILLER_4_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_2 FrameData[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_64 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput94 net96 VGND VGND VPWR VPWR FrameStrobe_O[16] sky130_fd_sc_hd__buf_2
Xoutput72 net74 VGND VGND VPWR VPWR FrameData_O[25] sky130_fd_sc_hd__buf_2
XFILLER_9_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput61 net63 VGND VGND VPWR VPWR FrameData_O[15] sky130_fd_sc_hd__buf_2
XFILLER_0_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput83 net85 VGND VGND VPWR VPWR FrameData_O[6] sky130_fd_sc_hd__buf_2
XFILLER_9_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_150_ net38 VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__buf_1
XFILLER_10_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_081_ net15 net22 VGND VGND VPWR VPWR Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_6_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_133_ FrameStrobe[12] VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__clkbuf_1
XFILLER_2_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_064_ _004_ _025_ _029_ VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__o21a_1
XFILLER_9_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_255 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_116_ net17 VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__buf_1
X_047_ net41 net45 net49 net53 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit23.Q Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit24.Q
+ VGND VGND VPWR VPWR _015_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_3 FrameData[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput95 net97 VGND VGND VPWR VPWR FrameStrobe_O[17] sky130_fd_sc_hd__buf_2
Xoutput73 net75 VGND VGND VPWR VPWR FrameData_O[26] sky130_fd_sc_hd__buf_2
Xoutput62 net64 VGND VGND VPWR VPWR FrameData_O[16] sky130_fd_sc_hd__buf_2
Xoutput84 net86 VGND VGND VPWR VPWR FrameData_O[7] sky130_fd_sc_hd__buf_2
XFILLER_10_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_080_ net14 net8 VGND VGND VPWR VPWR Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_8_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_132_ FrameStrobe[11] VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__clkbuf_1
XFILLER_2_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_063_ _026_ _027_ _028_ Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit18.Q Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit19.Q
+ VGND VGND VPWR VPWR _029_ sky130_fd_sc_hd__a221o_1
XFILLER_0_89 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_046_ _001_ _010_ _014_ VGND VGND VPWR VPWR net163 sky130_fd_sc_hd__o21a_1
X_115_ net16 VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__buf_1
XFILLER_7_267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_4 FrameData[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_292 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput96 net98 VGND VGND VPWR VPWR FrameStrobe_O[18] sky130_fd_sc_hd__buf_2
Xoutput74 net76 VGND VGND VPWR VPWR FrameData_O[27] sky130_fd_sc_hd__buf_2
Xoutput63 net65 VGND VGND VPWR VPWR FrameData_O[17] sky130_fd_sc_hd__buf_2
Xoutput85 net87 VGND VGND VPWR VPWR FrameData_O[8] sky130_fd_sc_hd__buf_2
.ends

