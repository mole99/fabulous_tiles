VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO DSP
  CLASS BLOCK ;
  FOREIGN DSP ;
  ORIGIN 0.000 0.000 ;
  SIZE 225.000 BY 450.000 ;
  PIN Tile_X0Y0_E1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 316.160 225.000 316.760 ;
    END
  END Tile_X0Y0_E1BEG[0]
  PIN Tile_X0Y0_E1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 317.520 225.000 318.120 ;
    END
  END Tile_X0Y0_E1BEG[1]
  PIN Tile_X0Y0_E1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 224.400 318.880 225.000 319.480 ;
    END
  END Tile_X0Y0_E1BEG[2]
  PIN Tile_X0Y0_E1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 320.240 225.000 320.840 ;
    END
  END Tile_X0Y0_E1BEG[3]
  PIN Tile_X0Y0_E1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.160 0.600 316.760 ;
    END
  END Tile_X0Y0_E1END[0]
  PIN Tile_X0Y0_E1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 317.520 0.600 318.120 ;
    END
  END Tile_X0Y0_E1END[1]
  PIN Tile_X0Y0_E1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 318.880 0.600 319.480 ;
    END
  END Tile_X0Y0_E1END[2]
  PIN Tile_X0Y0_E1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 320.240 0.600 320.840 ;
    END
  END Tile_X0Y0_E1END[3]
  PIN Tile_X0Y0_E2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 321.600 225.000 322.200 ;
    END
  END Tile_X0Y0_E2BEG[0]
  PIN Tile_X0Y0_E2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 322.960 225.000 323.560 ;
    END
  END Tile_X0Y0_E2BEG[1]
  PIN Tile_X0Y0_E2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 224.400 324.320 225.000 324.920 ;
    END
  END Tile_X0Y0_E2BEG[2]
  PIN Tile_X0Y0_E2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 325.680 225.000 326.280 ;
    END
  END Tile_X0Y0_E2BEG[3]
  PIN Tile_X0Y0_E2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 327.040 225.000 327.640 ;
    END
  END Tile_X0Y0_E2BEG[4]
  PIN Tile_X0Y0_E2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 328.400 225.000 329.000 ;
    END
  END Tile_X0Y0_E2BEG[5]
  PIN Tile_X0Y0_E2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 224.400 329.760 225.000 330.360 ;
    END
  END Tile_X0Y0_E2BEG[6]
  PIN Tile_X0Y0_E2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 331.120 225.000 331.720 ;
    END
  END Tile_X0Y0_E2BEG[7]
  PIN Tile_X0Y0_E2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 332.480 225.000 333.080 ;
    END
  END Tile_X0Y0_E2BEGb[0]
  PIN Tile_X0Y0_E2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 333.840 225.000 334.440 ;
    END
  END Tile_X0Y0_E2BEGb[1]
  PIN Tile_X0Y0_E2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 335.200 225.000 335.800 ;
    END
  END Tile_X0Y0_E2BEGb[2]
  PIN Tile_X0Y0_E2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 336.560 225.000 337.160 ;
    END
  END Tile_X0Y0_E2BEGb[3]
  PIN Tile_X0Y0_E2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 337.920 225.000 338.520 ;
    END
  END Tile_X0Y0_E2BEGb[4]
  PIN Tile_X0Y0_E2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 339.280 225.000 339.880 ;
    END
  END Tile_X0Y0_E2BEGb[5]
  PIN Tile_X0Y0_E2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 340.640 225.000 341.240 ;
    END
  END Tile_X0Y0_E2BEGb[6]
  PIN Tile_X0Y0_E2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 342.000 225.000 342.600 ;
    END
  END Tile_X0Y0_E2BEGb[7]
  PIN Tile_X0Y0_E2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 332.480 0.600 333.080 ;
    END
  END Tile_X0Y0_E2END[0]
  PIN Tile_X0Y0_E2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.840 0.600 334.440 ;
    END
  END Tile_X0Y0_E2END[1]
  PIN Tile_X0Y0_E2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 335.200 0.600 335.800 ;
    END
  END Tile_X0Y0_E2END[2]
  PIN Tile_X0Y0_E2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 336.560 0.600 337.160 ;
    END
  END Tile_X0Y0_E2END[3]
  PIN Tile_X0Y0_E2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 337.920 0.600 338.520 ;
    END
  END Tile_X0Y0_E2END[4]
  PIN Tile_X0Y0_E2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 339.280 0.600 339.880 ;
    END
  END Tile_X0Y0_E2END[5]
  PIN Tile_X0Y0_E2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.640 0.600 341.240 ;
    END
  END Tile_X0Y0_E2END[6]
  PIN Tile_X0Y0_E2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 342.000 0.600 342.600 ;
    END
  END Tile_X0Y0_E2END[7]
  PIN Tile_X0Y0_E2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 321.600 0.600 322.200 ;
    END
  END Tile_X0Y0_E2MID[0]
  PIN Tile_X0Y0_E2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 322.960 0.600 323.560 ;
    END
  END Tile_X0Y0_E2MID[1]
  PIN Tile_X0Y0_E2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 324.320 0.600 324.920 ;
    END
  END Tile_X0Y0_E2MID[2]
  PIN Tile_X0Y0_E2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 325.680 0.600 326.280 ;
    END
  END Tile_X0Y0_E2MID[3]
  PIN Tile_X0Y0_E2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 327.040 0.600 327.640 ;
    END
  END Tile_X0Y0_E2MID[4]
  PIN Tile_X0Y0_E2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 328.400 0.600 329.000 ;
    END
  END Tile_X0Y0_E2MID[5]
  PIN Tile_X0Y0_E2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 329.760 0.600 330.360 ;
    END
  END Tile_X0Y0_E2MID[6]
  PIN Tile_X0Y0_E2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 331.120 0.600 331.720 ;
    END
  END Tile_X0Y0_E2MID[7]
  PIN Tile_X0Y0_E6BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 365.120 225.000 365.720 ;
    END
  END Tile_X0Y0_E6BEG[0]
  PIN Tile_X0Y0_E6BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 224.400 378.720 225.000 379.320 ;
    END
  END Tile_X0Y0_E6BEG[10]
  PIN Tile_X0Y0_E6BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 380.080 225.000 380.680 ;
    END
  END Tile_X0Y0_E6BEG[11]
  PIN Tile_X0Y0_E6BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 366.480 225.000 367.080 ;
    END
  END Tile_X0Y0_E6BEG[1]
  PIN Tile_X0Y0_E6BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 367.840 225.000 368.440 ;
    END
  END Tile_X0Y0_E6BEG[2]
  PIN Tile_X0Y0_E6BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 369.200 225.000 369.800 ;
    END
  END Tile_X0Y0_E6BEG[3]
  PIN Tile_X0Y0_E6BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 370.560 225.000 371.160 ;
    END
  END Tile_X0Y0_E6BEG[4]
  PIN Tile_X0Y0_E6BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 371.920 225.000 372.520 ;
    END
  END Tile_X0Y0_E6BEG[5]
  PIN Tile_X0Y0_E6BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 373.280 225.000 373.880 ;
    END
  END Tile_X0Y0_E6BEG[6]
  PIN Tile_X0Y0_E6BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 374.640 225.000 375.240 ;
    END
  END Tile_X0Y0_E6BEG[7]
  PIN Tile_X0Y0_E6BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 376.000 225.000 376.600 ;
    END
  END Tile_X0Y0_E6BEG[8]
  PIN Tile_X0Y0_E6BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 377.360 225.000 377.960 ;
    END
  END Tile_X0Y0_E6BEG[9]
  PIN Tile_X0Y0_E6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 365.120 0.600 365.720 ;
    END
  END Tile_X0Y0_E6END[0]
  PIN Tile_X0Y0_E6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 378.720 0.600 379.320 ;
    END
  END Tile_X0Y0_E6END[10]
  PIN Tile_X0Y0_E6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.080 0.600 380.680 ;
    END
  END Tile_X0Y0_E6END[11]
  PIN Tile_X0Y0_E6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 366.480 0.600 367.080 ;
    END
  END Tile_X0Y0_E6END[1]
  PIN Tile_X0Y0_E6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 367.840 0.600 368.440 ;
    END
  END Tile_X0Y0_E6END[2]
  PIN Tile_X0Y0_E6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 369.200 0.600 369.800 ;
    END
  END Tile_X0Y0_E6END[3]
  PIN Tile_X0Y0_E6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 370.560 0.600 371.160 ;
    END
  END Tile_X0Y0_E6END[4]
  PIN Tile_X0Y0_E6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 371.920 0.600 372.520 ;
    END
  END Tile_X0Y0_E6END[5]
  PIN Tile_X0Y0_E6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 373.280 0.600 373.880 ;
    END
  END Tile_X0Y0_E6END[6]
  PIN Tile_X0Y0_E6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.640 0.600 375.240 ;
    END
  END Tile_X0Y0_E6END[7]
  PIN Tile_X0Y0_E6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 376.000 0.600 376.600 ;
    END
  END Tile_X0Y0_E6END[8]
  PIN Tile_X0Y0_E6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 377.360 0.600 377.960 ;
    END
  END Tile_X0Y0_E6END[9]
  PIN Tile_X0Y0_EE4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 343.360 225.000 343.960 ;
    END
  END Tile_X0Y0_EE4BEG[0]
  PIN Tile_X0Y0_EE4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 356.960 225.000 357.560 ;
    END
  END Tile_X0Y0_EE4BEG[10]
  PIN Tile_X0Y0_EE4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 358.320 225.000 358.920 ;
    END
  END Tile_X0Y0_EE4BEG[11]
  PIN Tile_X0Y0_EE4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 359.680 225.000 360.280 ;
    END
  END Tile_X0Y0_EE4BEG[12]
  PIN Tile_X0Y0_EE4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 224.400 361.040 225.000 361.640 ;
    END
  END Tile_X0Y0_EE4BEG[13]
  PIN Tile_X0Y0_EE4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 362.400 225.000 363.000 ;
    END
  END Tile_X0Y0_EE4BEG[14]
  PIN Tile_X0Y0_EE4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 224.400 363.760 225.000 364.360 ;
    END
  END Tile_X0Y0_EE4BEG[15]
  PIN Tile_X0Y0_EE4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 344.720 225.000 345.320 ;
    END
  END Tile_X0Y0_EE4BEG[1]
  PIN Tile_X0Y0_EE4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 346.080 225.000 346.680 ;
    END
  END Tile_X0Y0_EE4BEG[2]
  PIN Tile_X0Y0_EE4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 347.440 225.000 348.040 ;
    END
  END Tile_X0Y0_EE4BEG[3]
  PIN Tile_X0Y0_EE4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 348.800 225.000 349.400 ;
    END
  END Tile_X0Y0_EE4BEG[4]
  PIN Tile_X0Y0_EE4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 350.160 225.000 350.760 ;
    END
  END Tile_X0Y0_EE4BEG[5]
  PIN Tile_X0Y0_EE4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 351.520 225.000 352.120 ;
    END
  END Tile_X0Y0_EE4BEG[6]
  PIN Tile_X0Y0_EE4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 352.880 225.000 353.480 ;
    END
  END Tile_X0Y0_EE4BEG[7]
  PIN Tile_X0Y0_EE4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 354.240 225.000 354.840 ;
    END
  END Tile_X0Y0_EE4BEG[8]
  PIN Tile_X0Y0_EE4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 355.600 225.000 356.200 ;
    END
  END Tile_X0Y0_EE4BEG[9]
  PIN Tile_X0Y0_EE4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 343.360 0.600 343.960 ;
    END
  END Tile_X0Y0_EE4END[0]
  PIN Tile_X0Y0_EE4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 356.960 0.600 357.560 ;
    END
  END Tile_X0Y0_EE4END[10]
  PIN Tile_X0Y0_EE4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 358.320 0.600 358.920 ;
    END
  END Tile_X0Y0_EE4END[11]
  PIN Tile_X0Y0_EE4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 359.680 0.600 360.280 ;
    END
  END Tile_X0Y0_EE4END[12]
  PIN Tile_X0Y0_EE4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 361.040 0.600 361.640 ;
    END
  END Tile_X0Y0_EE4END[13]
  PIN Tile_X0Y0_EE4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 362.400 0.600 363.000 ;
    END
  END Tile_X0Y0_EE4END[14]
  PIN Tile_X0Y0_EE4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.760 0.600 364.360 ;
    END
  END Tile_X0Y0_EE4END[15]
  PIN Tile_X0Y0_EE4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 344.720 0.600 345.320 ;
    END
  END Tile_X0Y0_EE4END[1]
  PIN Tile_X0Y0_EE4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.080 0.600 346.680 ;
    END
  END Tile_X0Y0_EE4END[2]
  PIN Tile_X0Y0_EE4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 347.440 0.600 348.040 ;
    END
  END Tile_X0Y0_EE4END[3]
  PIN Tile_X0Y0_EE4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 348.800 0.600 349.400 ;
    END
  END Tile_X0Y0_EE4END[4]
  PIN Tile_X0Y0_EE4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.160 0.600 350.760 ;
    END
  END Tile_X0Y0_EE4END[5]
  PIN Tile_X0Y0_EE4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 351.520 0.600 352.120 ;
    END
  END Tile_X0Y0_EE4END[6]
  PIN Tile_X0Y0_EE4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 352.880 0.600 353.480 ;
    END
  END Tile_X0Y0_EE4END[7]
  PIN Tile_X0Y0_EE4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 354.240 0.600 354.840 ;
    END
  END Tile_X0Y0_EE4END[8]
  PIN Tile_X0Y0_EE4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 355.600 0.600 356.200 ;
    END
  END Tile_X0Y0_EE4END[9]
  PIN Tile_X0Y0_FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 381.440 0.600 382.040 ;
    END
  END Tile_X0Y0_FrameData[0]
  PIN Tile_X0Y0_FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 395.040 0.600 395.640 ;
    END
  END Tile_X0Y0_FrameData[10]
  PIN Tile_X0Y0_FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 396.400 0.600 397.000 ;
    END
  END Tile_X0Y0_FrameData[11]
  PIN Tile_X0Y0_FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 397.760 0.600 398.360 ;
    END
  END Tile_X0Y0_FrameData[12]
  PIN Tile_X0Y0_FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 399.120 0.600 399.720 ;
    END
  END Tile_X0Y0_FrameData[13]
  PIN Tile_X0Y0_FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 400.480 0.600 401.080 ;
    END
  END Tile_X0Y0_FrameData[14]
  PIN Tile_X0Y0_FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 401.840 0.600 402.440 ;
    END
  END Tile_X0Y0_FrameData[15]
  PIN Tile_X0Y0_FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 403.200 0.600 403.800 ;
    END
  END Tile_X0Y0_FrameData[16]
  PIN Tile_X0Y0_FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 404.560 0.600 405.160 ;
    END
  END Tile_X0Y0_FrameData[17]
  PIN Tile_X0Y0_FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 405.920 0.600 406.520 ;
    END
  END Tile_X0Y0_FrameData[18]
  PIN Tile_X0Y0_FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 407.280 0.600 407.880 ;
    END
  END Tile_X0Y0_FrameData[19]
  PIN Tile_X0Y0_FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 382.800 0.600 383.400 ;
    END
  END Tile_X0Y0_FrameData[1]
  PIN Tile_X0Y0_FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 408.640 0.600 409.240 ;
    END
  END Tile_X0Y0_FrameData[20]
  PIN Tile_X0Y0_FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 410.000 0.600 410.600 ;
    END
  END Tile_X0Y0_FrameData[21]
  PIN Tile_X0Y0_FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 411.360 0.600 411.960 ;
    END
  END Tile_X0Y0_FrameData[22]
  PIN Tile_X0Y0_FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 412.720 0.600 413.320 ;
    END
  END Tile_X0Y0_FrameData[23]
  PIN Tile_X0Y0_FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 414.080 0.600 414.680 ;
    END
  END Tile_X0Y0_FrameData[24]
  PIN Tile_X0Y0_FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 415.440 0.600 416.040 ;
    END
  END Tile_X0Y0_FrameData[25]
  PIN Tile_X0Y0_FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 416.800 0.600 417.400 ;
    END
  END Tile_X0Y0_FrameData[26]
  PIN Tile_X0Y0_FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 418.160 0.600 418.760 ;
    END
  END Tile_X0Y0_FrameData[27]
  PIN Tile_X0Y0_FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 419.520 0.600 420.120 ;
    END
  END Tile_X0Y0_FrameData[28]
  PIN Tile_X0Y0_FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 420.880 0.600 421.480 ;
    END
  END Tile_X0Y0_FrameData[29]
  PIN Tile_X0Y0_FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.160 0.600 384.760 ;
    END
  END Tile_X0Y0_FrameData[2]
  PIN Tile_X0Y0_FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 422.240 0.600 422.840 ;
    END
  END Tile_X0Y0_FrameData[30]
  PIN Tile_X0Y0_FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 423.600 0.600 424.200 ;
    END
  END Tile_X0Y0_FrameData[31]
  PIN Tile_X0Y0_FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 385.520 0.600 386.120 ;
    END
  END Tile_X0Y0_FrameData[3]
  PIN Tile_X0Y0_FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 386.880 0.600 387.480 ;
    END
  END Tile_X0Y0_FrameData[4]
  PIN Tile_X0Y0_FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 388.240 0.600 388.840 ;
    END
  END Tile_X0Y0_FrameData[5]
  PIN Tile_X0Y0_FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 389.600 0.600 390.200 ;
    END
  END Tile_X0Y0_FrameData[6]
  PIN Tile_X0Y0_FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 390.960 0.600 391.560 ;
    END
  END Tile_X0Y0_FrameData[7]
  PIN Tile_X0Y0_FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 392.320 0.600 392.920 ;
    END
  END Tile_X0Y0_FrameData[8]
  PIN Tile_X0Y0_FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 393.680 0.600 394.280 ;
    END
  END Tile_X0Y0_FrameData[9]
  PIN Tile_X0Y0_FrameData_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 381.440 225.000 382.040 ;
    END
  END Tile_X0Y0_FrameData_O[0]
  PIN Tile_X0Y0_FrameData_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 395.040 225.000 395.640 ;
    END
  END Tile_X0Y0_FrameData_O[10]
  PIN Tile_X0Y0_FrameData_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 396.400 225.000 397.000 ;
    END
  END Tile_X0Y0_FrameData_O[11]
  PIN Tile_X0Y0_FrameData_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 397.760 225.000 398.360 ;
    END
  END Tile_X0Y0_FrameData_O[12]
  PIN Tile_X0Y0_FrameData_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 399.120 225.000 399.720 ;
    END
  END Tile_X0Y0_FrameData_O[13]
  PIN Tile_X0Y0_FrameData_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 400.480 225.000 401.080 ;
    END
  END Tile_X0Y0_FrameData_O[14]
  PIN Tile_X0Y0_FrameData_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 401.840 225.000 402.440 ;
    END
  END Tile_X0Y0_FrameData_O[15]
  PIN Tile_X0Y0_FrameData_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 403.200 225.000 403.800 ;
    END
  END Tile_X0Y0_FrameData_O[16]
  PIN Tile_X0Y0_FrameData_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 404.560 225.000 405.160 ;
    END
  END Tile_X0Y0_FrameData_O[17]
  PIN Tile_X0Y0_FrameData_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 405.920 225.000 406.520 ;
    END
  END Tile_X0Y0_FrameData_O[18]
  PIN Tile_X0Y0_FrameData_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 407.280 225.000 407.880 ;
    END
  END Tile_X0Y0_FrameData_O[19]
  PIN Tile_X0Y0_FrameData_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 382.800 225.000 383.400 ;
    END
  END Tile_X0Y0_FrameData_O[1]
  PIN Tile_X0Y0_FrameData_O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 408.640 225.000 409.240 ;
    END
  END Tile_X0Y0_FrameData_O[20]
  PIN Tile_X0Y0_FrameData_O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 410.000 225.000 410.600 ;
    END
  END Tile_X0Y0_FrameData_O[21]
  PIN Tile_X0Y0_FrameData_O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 411.360 225.000 411.960 ;
    END
  END Tile_X0Y0_FrameData_O[22]
  PIN Tile_X0Y0_FrameData_O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 412.720 225.000 413.320 ;
    END
  END Tile_X0Y0_FrameData_O[23]
  PIN Tile_X0Y0_FrameData_O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 414.080 225.000 414.680 ;
    END
  END Tile_X0Y0_FrameData_O[24]
  PIN Tile_X0Y0_FrameData_O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 415.440 225.000 416.040 ;
    END
  END Tile_X0Y0_FrameData_O[25]
  PIN Tile_X0Y0_FrameData_O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 416.800 225.000 417.400 ;
    END
  END Tile_X0Y0_FrameData_O[26]
  PIN Tile_X0Y0_FrameData_O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 418.160 225.000 418.760 ;
    END
  END Tile_X0Y0_FrameData_O[27]
  PIN Tile_X0Y0_FrameData_O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 419.520 225.000 420.120 ;
    END
  END Tile_X0Y0_FrameData_O[28]
  PIN Tile_X0Y0_FrameData_O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 420.880 225.000 421.480 ;
    END
  END Tile_X0Y0_FrameData_O[29]
  PIN Tile_X0Y0_FrameData_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 384.160 225.000 384.760 ;
    END
  END Tile_X0Y0_FrameData_O[2]
  PIN Tile_X0Y0_FrameData_O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 422.240 225.000 422.840 ;
    END
  END Tile_X0Y0_FrameData_O[30]
  PIN Tile_X0Y0_FrameData_O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 423.600 225.000 424.200 ;
    END
  END Tile_X0Y0_FrameData_O[31]
  PIN Tile_X0Y0_FrameData_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 385.520 225.000 386.120 ;
    END
  END Tile_X0Y0_FrameData_O[3]
  PIN Tile_X0Y0_FrameData_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 386.880 225.000 387.480 ;
    END
  END Tile_X0Y0_FrameData_O[4]
  PIN Tile_X0Y0_FrameData_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 388.240 225.000 388.840 ;
    END
  END Tile_X0Y0_FrameData_O[5]
  PIN Tile_X0Y0_FrameData_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 389.600 225.000 390.200 ;
    END
  END Tile_X0Y0_FrameData_O[6]
  PIN Tile_X0Y0_FrameData_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 390.960 225.000 391.560 ;
    END
  END Tile_X0Y0_FrameData_O[7]
  PIN Tile_X0Y0_FrameData_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 392.320 225.000 392.920 ;
    END
  END Tile_X0Y0_FrameData_O[8]
  PIN Tile_X0Y0_FrameData_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 393.680 225.000 394.280 ;
    END
  END Tile_X0Y0_FrameData_O[9]
  PIN Tile_X0Y0_FrameStrobe_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 171.670 449.720 171.950 450.000 ;
    END
  END Tile_X0Y0_FrameStrobe_O[0]
  PIN Tile_X0Y0_FrameStrobe_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 185.470 449.720 185.750 450.000 ;
    END
  END Tile_X0Y0_FrameStrobe_O[10]
  PIN Tile_X0Y0_FrameStrobe_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 186.850 449.720 187.130 450.000 ;
    END
  END Tile_X0Y0_FrameStrobe_O[11]
  PIN Tile_X0Y0_FrameStrobe_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 188.230 449.720 188.510 450.000 ;
    END
  END Tile_X0Y0_FrameStrobe_O[12]
  PIN Tile_X0Y0_FrameStrobe_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 189.610 449.720 189.890 450.000 ;
    END
  END Tile_X0Y0_FrameStrobe_O[13]
  PIN Tile_X0Y0_FrameStrobe_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 190.990 449.720 191.270 450.000 ;
    END
  END Tile_X0Y0_FrameStrobe_O[14]
  PIN Tile_X0Y0_FrameStrobe_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 192.370 449.720 192.650 450.000 ;
    END
  END Tile_X0Y0_FrameStrobe_O[15]
  PIN Tile_X0Y0_FrameStrobe_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 193.750 449.720 194.030 450.000 ;
    END
  END Tile_X0Y0_FrameStrobe_O[16]
  PIN Tile_X0Y0_FrameStrobe_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 195.130 449.720 195.410 450.000 ;
    END
  END Tile_X0Y0_FrameStrobe_O[17]
  PIN Tile_X0Y0_FrameStrobe_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 196.510 449.720 196.790 450.000 ;
    END
  END Tile_X0Y0_FrameStrobe_O[18]
  PIN Tile_X0Y0_FrameStrobe_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 197.890 449.720 198.170 450.000 ;
    END
  END Tile_X0Y0_FrameStrobe_O[19]
  PIN Tile_X0Y0_FrameStrobe_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 173.050 449.720 173.330 450.000 ;
    END
  END Tile_X0Y0_FrameStrobe_O[1]
  PIN Tile_X0Y0_FrameStrobe_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 174.430 449.720 174.710 450.000 ;
    END
  END Tile_X0Y0_FrameStrobe_O[2]
  PIN Tile_X0Y0_FrameStrobe_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 175.810 449.720 176.090 450.000 ;
    END
  END Tile_X0Y0_FrameStrobe_O[3]
  PIN Tile_X0Y0_FrameStrobe_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 177.190 449.720 177.470 450.000 ;
    END
  END Tile_X0Y0_FrameStrobe_O[4]
  PIN Tile_X0Y0_FrameStrobe_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 178.570 449.720 178.850 450.000 ;
    END
  END Tile_X0Y0_FrameStrobe_O[5]
  PIN Tile_X0Y0_FrameStrobe_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 179.950 449.720 180.230 450.000 ;
    END
  END Tile_X0Y0_FrameStrobe_O[6]
  PIN Tile_X0Y0_FrameStrobe_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 181.330 449.720 181.610 450.000 ;
    END
  END Tile_X0Y0_FrameStrobe_O[7]
  PIN Tile_X0Y0_FrameStrobe_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 182.710 449.720 182.990 450.000 ;
    END
  END Tile_X0Y0_FrameStrobe_O[8]
  PIN Tile_X0Y0_FrameStrobe_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 184.090 449.720 184.370 450.000 ;
    END
  END Tile_X0Y0_FrameStrobe_O[9]
  PIN Tile_X0Y0_N1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 26.770 449.720 27.050 450.000 ;
    END
  END Tile_X0Y0_N1BEG[0]
  PIN Tile_X0Y0_N1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 28.150 449.720 28.430 450.000 ;
    END
  END Tile_X0Y0_N1BEG[1]
  PIN Tile_X0Y0_N1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 29.530 449.720 29.810 450.000 ;
    END
  END Tile_X0Y0_N1BEG[2]
  PIN Tile_X0Y0_N1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 30.910 449.720 31.190 450.000 ;
    END
  END Tile_X0Y0_N1BEG[3]
  PIN Tile_X0Y0_N2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 32.290 449.720 32.570 450.000 ;
    END
  END Tile_X0Y0_N2BEG[0]
  PIN Tile_X0Y0_N2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 33.670 449.720 33.950 450.000 ;
    END
  END Tile_X0Y0_N2BEG[1]
  PIN Tile_X0Y0_N2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 35.050 449.720 35.330 450.000 ;
    END
  END Tile_X0Y0_N2BEG[2]
  PIN Tile_X0Y0_N2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 36.430 449.720 36.710 450.000 ;
    END
  END Tile_X0Y0_N2BEG[3]
  PIN Tile_X0Y0_N2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 37.810 449.720 38.090 450.000 ;
    END
  END Tile_X0Y0_N2BEG[4]
  PIN Tile_X0Y0_N2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 39.190 449.720 39.470 450.000 ;
    END
  END Tile_X0Y0_N2BEG[5]
  PIN Tile_X0Y0_N2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 40.570 449.720 40.850 450.000 ;
    END
  END Tile_X0Y0_N2BEG[6]
  PIN Tile_X0Y0_N2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 41.950 449.720 42.230 450.000 ;
    END
  END Tile_X0Y0_N2BEG[7]
  PIN Tile_X0Y0_N2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 43.330 449.720 43.610 450.000 ;
    END
  END Tile_X0Y0_N2BEGb[0]
  PIN Tile_X0Y0_N2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 44.710 449.720 44.990 450.000 ;
    END
  END Tile_X0Y0_N2BEGb[1]
  PIN Tile_X0Y0_N2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 46.090 449.720 46.370 450.000 ;
    END
  END Tile_X0Y0_N2BEGb[2]
  PIN Tile_X0Y0_N2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 47.470 449.720 47.750 450.000 ;
    END
  END Tile_X0Y0_N2BEGb[3]
  PIN Tile_X0Y0_N2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 48.850 449.720 49.130 450.000 ;
    END
  END Tile_X0Y0_N2BEGb[4]
  PIN Tile_X0Y0_N2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 50.230 449.720 50.510 450.000 ;
    END
  END Tile_X0Y0_N2BEGb[5]
  PIN Tile_X0Y0_N2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 51.610 449.720 51.890 450.000 ;
    END
  END Tile_X0Y0_N2BEGb[6]
  PIN Tile_X0Y0_N2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 52.990 449.720 53.270 450.000 ;
    END
  END Tile_X0Y0_N2BEGb[7]
  PIN Tile_X0Y0_N4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 54.370 449.720 54.650 450.000 ;
    END
  END Tile_X0Y0_N4BEG[0]
  PIN Tile_X0Y0_N4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 68.170 449.720 68.450 450.000 ;
    END
  END Tile_X0Y0_N4BEG[10]
  PIN Tile_X0Y0_N4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 69.550 449.720 69.830 450.000 ;
    END
  END Tile_X0Y0_N4BEG[11]
  PIN Tile_X0Y0_N4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 70.930 449.720 71.210 450.000 ;
    END
  END Tile_X0Y0_N4BEG[12]
  PIN Tile_X0Y0_N4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 72.310 449.720 72.590 450.000 ;
    END
  END Tile_X0Y0_N4BEG[13]
  PIN Tile_X0Y0_N4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 73.690 449.720 73.970 450.000 ;
    END
  END Tile_X0Y0_N4BEG[14]
  PIN Tile_X0Y0_N4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 75.070 449.720 75.350 450.000 ;
    END
  END Tile_X0Y0_N4BEG[15]
  PIN Tile_X0Y0_N4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 55.750 449.720 56.030 450.000 ;
    END
  END Tile_X0Y0_N4BEG[1]
  PIN Tile_X0Y0_N4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 57.130 449.720 57.410 450.000 ;
    END
  END Tile_X0Y0_N4BEG[2]
  PIN Tile_X0Y0_N4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 58.510 449.720 58.790 450.000 ;
    END
  END Tile_X0Y0_N4BEG[3]
  PIN Tile_X0Y0_N4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 59.890 449.720 60.170 450.000 ;
    END
  END Tile_X0Y0_N4BEG[4]
  PIN Tile_X0Y0_N4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 61.270 449.720 61.550 450.000 ;
    END
  END Tile_X0Y0_N4BEG[5]
  PIN Tile_X0Y0_N4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 62.650 449.720 62.930 450.000 ;
    END
  END Tile_X0Y0_N4BEG[6]
  PIN Tile_X0Y0_N4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 64.030 449.720 64.310 450.000 ;
    END
  END Tile_X0Y0_N4BEG[7]
  PIN Tile_X0Y0_N4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 65.410 449.720 65.690 450.000 ;
    END
  END Tile_X0Y0_N4BEG[8]
  PIN Tile_X0Y0_N4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 66.790 449.720 67.070 450.000 ;
    END
  END Tile_X0Y0_N4BEG[9]
  PIN Tile_X0Y0_NN4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 76.450 449.720 76.730 450.000 ;
    END
  END Tile_X0Y0_NN4BEG[0]
  PIN Tile_X0Y0_NN4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 90.250 449.720 90.530 450.000 ;
    END
  END Tile_X0Y0_NN4BEG[10]
  PIN Tile_X0Y0_NN4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 91.630 449.720 91.910 450.000 ;
    END
  END Tile_X0Y0_NN4BEG[11]
  PIN Tile_X0Y0_NN4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 93.010 449.720 93.290 450.000 ;
    END
  END Tile_X0Y0_NN4BEG[12]
  PIN Tile_X0Y0_NN4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 94.390 449.720 94.670 450.000 ;
    END
  END Tile_X0Y0_NN4BEG[13]
  PIN Tile_X0Y0_NN4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 95.770 449.720 96.050 450.000 ;
    END
  END Tile_X0Y0_NN4BEG[14]
  PIN Tile_X0Y0_NN4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 97.150 449.720 97.430 450.000 ;
    END
  END Tile_X0Y0_NN4BEG[15]
  PIN Tile_X0Y0_NN4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 77.830 449.720 78.110 450.000 ;
    END
  END Tile_X0Y0_NN4BEG[1]
  PIN Tile_X0Y0_NN4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 79.210 449.720 79.490 450.000 ;
    END
  END Tile_X0Y0_NN4BEG[2]
  PIN Tile_X0Y0_NN4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 80.590 449.720 80.870 450.000 ;
    END
  END Tile_X0Y0_NN4BEG[3]
  PIN Tile_X0Y0_NN4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 81.970 449.720 82.250 450.000 ;
    END
  END Tile_X0Y0_NN4BEG[4]
  PIN Tile_X0Y0_NN4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 83.350 449.720 83.630 450.000 ;
    END
  END Tile_X0Y0_NN4BEG[5]
  PIN Tile_X0Y0_NN4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 84.730 449.720 85.010 450.000 ;
    END
  END Tile_X0Y0_NN4BEG[6]
  PIN Tile_X0Y0_NN4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 86.110 449.720 86.390 450.000 ;
    END
  END Tile_X0Y0_NN4BEG[7]
  PIN Tile_X0Y0_NN4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 87.490 449.720 87.770 450.000 ;
    END
  END Tile_X0Y0_NN4BEG[8]
  PIN Tile_X0Y0_NN4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 88.870 449.720 89.150 450.000 ;
    END
  END Tile_X0Y0_NN4BEG[9]
  PIN Tile_X0Y0_S1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 98.530 449.720 98.810 450.000 ;
    END
  END Tile_X0Y0_S1END[0]
  PIN Tile_X0Y0_S1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 99.910 449.720 100.190 450.000 ;
    END
  END Tile_X0Y0_S1END[1]
  PIN Tile_X0Y0_S1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 101.290 449.720 101.570 450.000 ;
    END
  END Tile_X0Y0_S1END[2]
  PIN Tile_X0Y0_S1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 102.670 449.720 102.950 450.000 ;
    END
  END Tile_X0Y0_S1END[3]
  PIN Tile_X0Y0_S2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 115.090 449.720 115.370 450.000 ;
    END
  END Tile_X0Y0_S2END[0]
  PIN Tile_X0Y0_S2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 116.470 449.720 116.750 450.000 ;
    END
  END Tile_X0Y0_S2END[1]
  PIN Tile_X0Y0_S2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 117.850 449.720 118.130 450.000 ;
    END
  END Tile_X0Y0_S2END[2]
  PIN Tile_X0Y0_S2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 119.230 449.720 119.510 450.000 ;
    END
  END Tile_X0Y0_S2END[3]
  PIN Tile_X0Y0_S2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 120.610 449.720 120.890 450.000 ;
    END
  END Tile_X0Y0_S2END[4]
  PIN Tile_X0Y0_S2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 121.990 449.720 122.270 450.000 ;
    END
  END Tile_X0Y0_S2END[5]
  PIN Tile_X0Y0_S2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 123.370 449.720 123.650 450.000 ;
    END
  END Tile_X0Y0_S2END[6]
  PIN Tile_X0Y0_S2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 124.750 449.720 125.030 450.000 ;
    END
  END Tile_X0Y0_S2END[7]
  PIN Tile_X0Y0_S2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 104.050 449.720 104.330 450.000 ;
    END
  END Tile_X0Y0_S2MID[0]
  PIN Tile_X0Y0_S2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 105.430 449.720 105.710 450.000 ;
    END
  END Tile_X0Y0_S2MID[1]
  PIN Tile_X0Y0_S2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 106.810 449.720 107.090 450.000 ;
    END
  END Tile_X0Y0_S2MID[2]
  PIN Tile_X0Y0_S2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 108.190 449.720 108.470 450.000 ;
    END
  END Tile_X0Y0_S2MID[3]
  PIN Tile_X0Y0_S2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 109.570 449.720 109.850 450.000 ;
    END
  END Tile_X0Y0_S2MID[4]
  PIN Tile_X0Y0_S2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 110.950 449.720 111.230 450.000 ;
    END
  END Tile_X0Y0_S2MID[5]
  PIN Tile_X0Y0_S2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 112.330 449.720 112.610 450.000 ;
    END
  END Tile_X0Y0_S2MID[6]
  PIN Tile_X0Y0_S2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 113.710 449.720 113.990 450.000 ;
    END
  END Tile_X0Y0_S2MID[7]
  PIN Tile_X0Y0_S4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 126.130 449.720 126.410 450.000 ;
    END
  END Tile_X0Y0_S4END[0]
  PIN Tile_X0Y0_S4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 139.930 449.720 140.210 450.000 ;
    END
  END Tile_X0Y0_S4END[10]
  PIN Tile_X0Y0_S4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.065900 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 141.310 449.720 141.590 450.000 ;
    END
  END Tile_X0Y0_S4END[11]
  PIN Tile_X0Y0_S4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 142.690 449.720 142.970 450.000 ;
    END
  END Tile_X0Y0_S4END[12]
  PIN Tile_X0Y0_S4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 144.070 449.720 144.350 450.000 ;
    END
  END Tile_X0Y0_S4END[13]
  PIN Tile_X0Y0_S4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 145.450 449.720 145.730 450.000 ;
    END
  END Tile_X0Y0_S4END[14]
  PIN Tile_X0Y0_S4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 146.830 449.720 147.110 450.000 ;
    END
  END Tile_X0Y0_S4END[15]
  PIN Tile_X0Y0_S4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 127.510 449.720 127.790 450.000 ;
    END
  END Tile_X0Y0_S4END[1]
  PIN Tile_X0Y0_S4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 128.890 449.720 129.170 450.000 ;
    END
  END Tile_X0Y0_S4END[2]
  PIN Tile_X0Y0_S4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 130.270 449.720 130.550 450.000 ;
    END
  END Tile_X0Y0_S4END[3]
  PIN Tile_X0Y0_S4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 131.650 449.720 131.930 450.000 ;
    END
  END Tile_X0Y0_S4END[4]
  PIN Tile_X0Y0_S4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 133.030 449.720 133.310 450.000 ;
    END
  END Tile_X0Y0_S4END[5]
  PIN Tile_X0Y0_S4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 134.410 449.720 134.690 450.000 ;
    END
  END Tile_X0Y0_S4END[6]
  PIN Tile_X0Y0_S4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 135.790 449.720 136.070 450.000 ;
    END
  END Tile_X0Y0_S4END[7]
  PIN Tile_X0Y0_S4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.065900 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 137.170 449.720 137.450 450.000 ;
    END
  END Tile_X0Y0_S4END[8]
  PIN Tile_X0Y0_S4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 138.550 449.720 138.830 450.000 ;
    END
  END Tile_X0Y0_S4END[9]
  PIN Tile_X0Y0_SS4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 148.210 449.720 148.490 450.000 ;
    END
  END Tile_X0Y0_SS4END[0]
  PIN Tile_X0Y0_SS4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 162.010 449.720 162.290 450.000 ;
    END
  END Tile_X0Y0_SS4END[10]
  PIN Tile_X0Y0_SS4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 163.390 449.720 163.670 450.000 ;
    END
  END Tile_X0Y0_SS4END[11]
  PIN Tile_X0Y0_SS4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 164.770 449.720 165.050 450.000 ;
    END
  END Tile_X0Y0_SS4END[12]
  PIN Tile_X0Y0_SS4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 166.150 449.720 166.430 450.000 ;
    END
  END Tile_X0Y0_SS4END[13]
  PIN Tile_X0Y0_SS4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 167.530 449.720 167.810 450.000 ;
    END
  END Tile_X0Y0_SS4END[14]
  PIN Tile_X0Y0_SS4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 168.910 449.720 169.190 450.000 ;
    END
  END Tile_X0Y0_SS4END[15]
  PIN Tile_X0Y0_SS4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 149.590 449.720 149.870 450.000 ;
    END
  END Tile_X0Y0_SS4END[1]
  PIN Tile_X0Y0_SS4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 150.970 449.720 151.250 450.000 ;
    END
  END Tile_X0Y0_SS4END[2]
  PIN Tile_X0Y0_SS4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 152.350 449.720 152.630 450.000 ;
    END
  END Tile_X0Y0_SS4END[3]
  PIN Tile_X0Y0_SS4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 153.730 449.720 154.010 450.000 ;
    END
  END Tile_X0Y0_SS4END[4]
  PIN Tile_X0Y0_SS4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 155.110 449.720 155.390 450.000 ;
    END
  END Tile_X0Y0_SS4END[5]
  PIN Tile_X0Y0_SS4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 156.490 449.720 156.770 450.000 ;
    END
  END Tile_X0Y0_SS4END[6]
  PIN Tile_X0Y0_SS4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 157.870 449.720 158.150 450.000 ;
    END
  END Tile_X0Y0_SS4END[7]
  PIN Tile_X0Y0_SS4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 159.250 449.720 159.530 450.000 ;
    END
  END Tile_X0Y0_SS4END[8]
  PIN Tile_X0Y0_SS4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 160.630 449.720 160.910 450.000 ;
    END
  END Tile_X0Y0_SS4END[9]
  PIN Tile_X0Y0_UserCLKo
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 170.290 449.720 170.570 450.000 ;
    END
  END Tile_X0Y0_UserCLKo
  PIN Tile_X0Y0_W1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 250.880 0.600 251.480 ;
    END
  END Tile_X0Y0_W1BEG[0]
  PIN Tile_X0Y0_W1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 252.240 0.600 252.840 ;
    END
  END Tile_X0Y0_W1BEG[1]
  PIN Tile_X0Y0_W1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 253.600 0.600 254.200 ;
    END
  END Tile_X0Y0_W1BEG[2]
  PIN Tile_X0Y0_W1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 254.960 0.600 255.560 ;
    END
  END Tile_X0Y0_W1BEG[3]
  PIN Tile_X0Y0_W1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 224.400 250.880 225.000 251.480 ;
    END
  END Tile_X0Y0_W1END[0]
  PIN Tile_X0Y0_W1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 252.240 225.000 252.840 ;
    END
  END Tile_X0Y0_W1END[1]
  PIN Tile_X0Y0_W1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 224.400 253.600 225.000 254.200 ;
    END
  END Tile_X0Y0_W1END[2]
  PIN Tile_X0Y0_W1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 224.400 254.960 225.000 255.560 ;
    END
  END Tile_X0Y0_W1END[3]
  PIN Tile_X0Y0_W2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 256.320 0.600 256.920 ;
    END
  END Tile_X0Y0_W2BEG[0]
  PIN Tile_X0Y0_W2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 257.680 0.600 258.280 ;
    END
  END Tile_X0Y0_W2BEG[1]
  PIN Tile_X0Y0_W2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 259.040 0.600 259.640 ;
    END
  END Tile_X0Y0_W2BEG[2]
  PIN Tile_X0Y0_W2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 260.400 0.600 261.000 ;
    END
  END Tile_X0Y0_W2BEG[3]
  PIN Tile_X0Y0_W2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.760 0.600 262.360 ;
    END
  END Tile_X0Y0_W2BEG[4]
  PIN Tile_X0Y0_W2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 263.120 0.600 263.720 ;
    END
  END Tile_X0Y0_W2BEG[5]
  PIN Tile_X0Y0_W2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 264.480 0.600 265.080 ;
    END
  END Tile_X0Y0_W2BEG[6]
  PIN Tile_X0Y0_W2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.840 0.600 266.440 ;
    END
  END Tile_X0Y0_W2BEG[7]
  PIN Tile_X0Y0_W2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 267.200 0.600 267.800 ;
    END
  END Tile_X0Y0_W2BEGb[0]
  PIN Tile_X0Y0_W2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 268.560 0.600 269.160 ;
    END
  END Tile_X0Y0_W2BEGb[1]
  PIN Tile_X0Y0_W2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 269.920 0.600 270.520 ;
    END
  END Tile_X0Y0_W2BEGb[2]
  PIN Tile_X0Y0_W2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 271.280 0.600 271.880 ;
    END
  END Tile_X0Y0_W2BEGb[3]
  PIN Tile_X0Y0_W2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.640 0.600 273.240 ;
    END
  END Tile_X0Y0_W2BEGb[4]
  PIN Tile_X0Y0_W2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 274.000 0.600 274.600 ;
    END
  END Tile_X0Y0_W2BEGb[5]
  PIN Tile_X0Y0_W2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 275.360 0.600 275.960 ;
    END
  END Tile_X0Y0_W2BEGb[6]
  PIN Tile_X0Y0_W2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 276.720 0.600 277.320 ;
    END
  END Tile_X0Y0_W2BEGb[7]
  PIN Tile_X0Y0_W2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 224.400 267.200 225.000 267.800 ;
    END
  END Tile_X0Y0_W2END[0]
  PIN Tile_X0Y0_W2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 224.400 268.560 225.000 269.160 ;
    END
  END Tile_X0Y0_W2END[1]
  PIN Tile_X0Y0_W2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 224.400 269.920 225.000 270.520 ;
    END
  END Tile_X0Y0_W2END[2]
  PIN Tile_X0Y0_W2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 224.400 271.280 225.000 271.880 ;
    END
  END Tile_X0Y0_W2END[3]
  PIN Tile_X0Y0_W2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 224.400 272.640 225.000 273.240 ;
    END
  END Tile_X0Y0_W2END[4]
  PIN Tile_X0Y0_W2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 224.400 274.000 225.000 274.600 ;
    END
  END Tile_X0Y0_W2END[5]
  PIN Tile_X0Y0_W2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 224.400 275.360 225.000 275.960 ;
    END
  END Tile_X0Y0_W2END[6]
  PIN Tile_X0Y0_W2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 224.400 276.720 225.000 277.320 ;
    END
  END Tile_X0Y0_W2END[7]
  PIN Tile_X0Y0_W2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 224.400 256.320 225.000 256.920 ;
    END
  END Tile_X0Y0_W2MID[0]
  PIN Tile_X0Y0_W2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 224.400 257.680 225.000 258.280 ;
    END
  END Tile_X0Y0_W2MID[1]
  PIN Tile_X0Y0_W2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 224.400 259.040 225.000 259.640 ;
    END
  END Tile_X0Y0_W2MID[2]
  PIN Tile_X0Y0_W2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 224.400 260.400 225.000 261.000 ;
    END
  END Tile_X0Y0_W2MID[3]
  PIN Tile_X0Y0_W2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 224.400 261.760 225.000 262.360 ;
    END
  END Tile_X0Y0_W2MID[4]
  PIN Tile_X0Y0_W2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 224.400 263.120 225.000 263.720 ;
    END
  END Tile_X0Y0_W2MID[5]
  PIN Tile_X0Y0_W2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 224.400 264.480 225.000 265.080 ;
    END
  END Tile_X0Y0_W2MID[6]
  PIN Tile_X0Y0_W2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 224.400 265.840 225.000 266.440 ;
    END
  END Tile_X0Y0_W2MID[7]
  PIN Tile_X0Y0_W6BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.840 0.600 300.440 ;
    END
  END Tile_X0Y0_W6BEG[0]
  PIN Tile_X0Y0_W6BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 313.440 0.600 314.040 ;
    END
  END Tile_X0Y0_W6BEG[10]
  PIN Tile_X0Y0_W6BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 314.800 0.600 315.400 ;
    END
  END Tile_X0Y0_W6BEG[11]
  PIN Tile_X0Y0_W6BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 301.200 0.600 301.800 ;
    END
  END Tile_X0Y0_W6BEG[1]
  PIN Tile_X0Y0_W6BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 302.560 0.600 303.160 ;
    END
  END Tile_X0Y0_W6BEG[2]
  PIN Tile_X0Y0_W6BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 303.920 0.600 304.520 ;
    END
  END Tile_X0Y0_W6BEG[3]
  PIN Tile_X0Y0_W6BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 305.280 0.600 305.880 ;
    END
  END Tile_X0Y0_W6BEG[4]
  PIN Tile_X0Y0_W6BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 306.640 0.600 307.240 ;
    END
  END Tile_X0Y0_W6BEG[5]
  PIN Tile_X0Y0_W6BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 308.000 0.600 308.600 ;
    END
  END Tile_X0Y0_W6BEG[6]
  PIN Tile_X0Y0_W6BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 309.360 0.600 309.960 ;
    END
  END Tile_X0Y0_W6BEG[7]
  PIN Tile_X0Y0_W6BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 310.720 0.600 311.320 ;
    END
  END Tile_X0Y0_W6BEG[8]
  PIN Tile_X0Y0_W6BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.080 0.600 312.680 ;
    END
  END Tile_X0Y0_W6BEG[9]
  PIN Tile_X0Y0_W6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 224.400 299.840 225.000 300.440 ;
    END
  END Tile_X0Y0_W6END[0]
  PIN Tile_X0Y0_W6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 313.440 225.000 314.040 ;
    END
  END Tile_X0Y0_W6END[10]
  PIN Tile_X0Y0_W6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 314.800 225.000 315.400 ;
    END
  END Tile_X0Y0_W6END[11]
  PIN Tile_X0Y0_W6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 301.200 225.000 301.800 ;
    END
  END Tile_X0Y0_W6END[1]
  PIN Tile_X0Y0_W6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 302.560 225.000 303.160 ;
    END
  END Tile_X0Y0_W6END[2]
  PIN Tile_X0Y0_W6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 224.400 303.920 225.000 304.520 ;
    END
  END Tile_X0Y0_W6END[3]
  PIN Tile_X0Y0_W6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 305.280 225.000 305.880 ;
    END
  END Tile_X0Y0_W6END[4]
  PIN Tile_X0Y0_W6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 306.640 225.000 307.240 ;
    END
  END Tile_X0Y0_W6END[5]
  PIN Tile_X0Y0_W6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 224.400 308.000 225.000 308.600 ;
    END
  END Tile_X0Y0_W6END[6]
  PIN Tile_X0Y0_W6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 309.360 225.000 309.960 ;
    END
  END Tile_X0Y0_W6END[7]
  PIN Tile_X0Y0_W6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 310.720 225.000 311.320 ;
    END
  END Tile_X0Y0_W6END[8]
  PIN Tile_X0Y0_W6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 312.080 225.000 312.680 ;
    END
  END Tile_X0Y0_W6END[9]
  PIN Tile_X0Y0_WW4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.080 0.600 278.680 ;
    END
  END Tile_X0Y0_WW4BEG[0]
  PIN Tile_X0Y0_WW4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 291.680 0.600 292.280 ;
    END
  END Tile_X0Y0_WW4BEG[10]
  PIN Tile_X0Y0_WW4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 293.040 0.600 293.640 ;
    END
  END Tile_X0Y0_WW4BEG[11]
  PIN Tile_X0Y0_WW4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 294.400 0.600 295.000 ;
    END
  END Tile_X0Y0_WW4BEG[12]
  PIN Tile_X0Y0_WW4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.760 0.600 296.360 ;
    END
  END Tile_X0Y0_WW4BEG[13]
  PIN Tile_X0Y0_WW4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 297.120 0.600 297.720 ;
    END
  END Tile_X0Y0_WW4BEG[14]
  PIN Tile_X0Y0_WW4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 298.480 0.600 299.080 ;
    END
  END Tile_X0Y0_WW4BEG[15]
  PIN Tile_X0Y0_WW4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 279.440 0.600 280.040 ;
    END
  END Tile_X0Y0_WW4BEG[1]
  PIN Tile_X0Y0_WW4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 280.800 0.600 281.400 ;
    END
  END Tile_X0Y0_WW4BEG[2]
  PIN Tile_X0Y0_WW4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.160 0.600 282.760 ;
    END
  END Tile_X0Y0_WW4BEG[3]
  PIN Tile_X0Y0_WW4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 283.520 0.600 284.120 ;
    END
  END Tile_X0Y0_WW4BEG[4]
  PIN Tile_X0Y0_WW4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 284.880 0.600 285.480 ;
    END
  END Tile_X0Y0_WW4BEG[5]
  PIN Tile_X0Y0_WW4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 286.240 0.600 286.840 ;
    END
  END Tile_X0Y0_WW4BEG[6]
  PIN Tile_X0Y0_WW4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 287.600 0.600 288.200 ;
    END
  END Tile_X0Y0_WW4BEG[7]
  PIN Tile_X0Y0_WW4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 288.960 0.600 289.560 ;
    END
  END Tile_X0Y0_WW4BEG[8]
  PIN Tile_X0Y0_WW4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 290.320 0.600 290.920 ;
    END
  END Tile_X0Y0_WW4BEG[9]
  PIN Tile_X0Y0_WW4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 224.400 278.080 225.000 278.680 ;
    END
  END Tile_X0Y0_WW4END[0]
  PIN Tile_X0Y0_WW4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 291.680 225.000 292.280 ;
    END
  END Tile_X0Y0_WW4END[10]
  PIN Tile_X0Y0_WW4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 293.040 225.000 293.640 ;
    END
  END Tile_X0Y0_WW4END[11]
  PIN Tile_X0Y0_WW4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 294.400 225.000 295.000 ;
    END
  END Tile_X0Y0_WW4END[12]
  PIN Tile_X0Y0_WW4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 295.760 225.000 296.360 ;
    END
  END Tile_X0Y0_WW4END[13]
  PIN Tile_X0Y0_WW4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 297.120 225.000 297.720 ;
    END
  END Tile_X0Y0_WW4END[14]
  PIN Tile_X0Y0_WW4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 298.480 225.000 299.080 ;
    END
  END Tile_X0Y0_WW4END[15]
  PIN Tile_X0Y0_WW4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 224.400 279.440 225.000 280.040 ;
    END
  END Tile_X0Y0_WW4END[1]
  PIN Tile_X0Y0_WW4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 224.400 280.800 225.000 281.400 ;
    END
  END Tile_X0Y0_WW4END[2]
  PIN Tile_X0Y0_WW4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 224.400 282.160 225.000 282.760 ;
    END
  END Tile_X0Y0_WW4END[3]
  PIN Tile_X0Y0_WW4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 283.520 225.000 284.120 ;
    END
  END Tile_X0Y0_WW4END[4]
  PIN Tile_X0Y0_WW4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 284.880 225.000 285.480 ;
    END
  END Tile_X0Y0_WW4END[5]
  PIN Tile_X0Y0_WW4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 286.240 225.000 286.840 ;
    END
  END Tile_X0Y0_WW4END[6]
  PIN Tile_X0Y0_WW4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 224.400 287.600 225.000 288.200 ;
    END
  END Tile_X0Y0_WW4END[7]
  PIN Tile_X0Y0_WW4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 224.400 288.960 225.000 289.560 ;
    END
  END Tile_X0Y0_WW4END[8]
  PIN Tile_X0Y0_WW4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 290.320 225.000 290.920 ;
    END
  END Tile_X0Y0_WW4END[9]
  PIN Tile_X0Y1_E1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 91.160 225.000 91.760 ;
    END
  END Tile_X0Y1_E1BEG[0]
  PIN Tile_X0Y1_E1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 92.520 225.000 93.120 ;
    END
  END Tile_X0Y1_E1BEG[1]
  PIN Tile_X0Y1_E1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 93.880 225.000 94.480 ;
    END
  END Tile_X0Y1_E1BEG[2]
  PIN Tile_X0Y1_E1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 95.240 225.000 95.840 ;
    END
  END Tile_X0Y1_E1BEG[3]
  PIN Tile_X0Y1_E1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.160 0.600 91.760 ;
    END
  END Tile_X0Y1_E1END[0]
  PIN Tile_X0Y1_E1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.520 0.600 93.120 ;
    END
  END Tile_X0Y1_E1END[1]
  PIN Tile_X0Y1_E1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.880 0.600 94.480 ;
    END
  END Tile_X0Y1_E1END[2]
  PIN Tile_X0Y1_E1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 0.600 95.840 ;
    END
  END Tile_X0Y1_E1END[3]
  PIN Tile_X0Y1_E2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 96.600 225.000 97.200 ;
    END
  END Tile_X0Y1_E2BEG[0]
  PIN Tile_X0Y1_E2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 97.960 225.000 98.560 ;
    END
  END Tile_X0Y1_E2BEG[1]
  PIN Tile_X0Y1_E2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 99.320 225.000 99.920 ;
    END
  END Tile_X0Y1_E2BEG[2]
  PIN Tile_X0Y1_E2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 100.680 225.000 101.280 ;
    END
  END Tile_X0Y1_E2BEG[3]
  PIN Tile_X0Y1_E2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 102.040 225.000 102.640 ;
    END
  END Tile_X0Y1_E2BEG[4]
  PIN Tile_X0Y1_E2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 103.400 225.000 104.000 ;
    END
  END Tile_X0Y1_E2BEG[5]
  PIN Tile_X0Y1_E2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.400 104.760 225.000 105.360 ;
    END
  END Tile_X0Y1_E2BEG[6]
  PIN Tile_X0Y1_E2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 106.120 225.000 106.720 ;
    END
  END Tile_X0Y1_E2BEG[7]
  PIN Tile_X0Y1_E2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 107.480 225.000 108.080 ;
    END
  END Tile_X0Y1_E2BEGb[0]
  PIN Tile_X0Y1_E2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 108.840 225.000 109.440 ;
    END
  END Tile_X0Y1_E2BEGb[1]
  PIN Tile_X0Y1_E2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 110.200 225.000 110.800 ;
    END
  END Tile_X0Y1_E2BEGb[2]
  PIN Tile_X0Y1_E2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 111.560 225.000 112.160 ;
    END
  END Tile_X0Y1_E2BEGb[3]
  PIN Tile_X0Y1_E2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 112.920 225.000 113.520 ;
    END
  END Tile_X0Y1_E2BEGb[4]
  PIN Tile_X0Y1_E2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 114.280 225.000 114.880 ;
    END
  END Tile_X0Y1_E2BEGb[5]
  PIN Tile_X0Y1_E2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 115.640 225.000 116.240 ;
    END
  END Tile_X0Y1_E2BEGb[6]
  PIN Tile_X0Y1_E2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 117.000 225.000 117.600 ;
    END
  END Tile_X0Y1_E2BEGb[7]
  PIN Tile_X0Y1_E2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 107.480 0.600 108.080 ;
    END
  END Tile_X0Y1_E2END[0]
  PIN Tile_X0Y1_E2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 0.600 109.440 ;
    END
  END Tile_X0Y1_E2END[1]
  PIN Tile_X0Y1_E2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.200 0.600 110.800 ;
    END
  END Tile_X0Y1_E2END[2]
  PIN Tile_X0Y1_E2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 111.560 0.600 112.160 ;
    END
  END Tile_X0Y1_E2END[3]
  PIN Tile_X0Y1_E2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.920 0.600 113.520 ;
    END
  END Tile_X0Y1_E2END[4]
  PIN Tile_X0Y1_E2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.280 0.600 114.880 ;
    END
  END Tile_X0Y1_E2END[5]
  PIN Tile_X0Y1_E2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 0.600 116.240 ;
    END
  END Tile_X0Y1_E2END[6]
  PIN Tile_X0Y1_E2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.000 0.600 117.600 ;
    END
  END Tile_X0Y1_E2END[7]
  PIN Tile_X0Y1_E2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 96.600 0.600 97.200 ;
    END
  END Tile_X0Y1_E2MID[0]
  PIN Tile_X0Y1_E2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.960 0.600 98.560 ;
    END
  END Tile_X0Y1_E2MID[1]
  PIN Tile_X0Y1_E2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 99.320 0.600 99.920 ;
    END
  END Tile_X0Y1_E2MID[2]
  PIN Tile_X0Y1_E2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.680 0.600 101.280 ;
    END
  END Tile_X0Y1_E2MID[3]
  PIN Tile_X0Y1_E2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 0.600 102.640 ;
    END
  END Tile_X0Y1_E2MID[4]
  PIN Tile_X0Y1_E2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 103.400 0.600 104.000 ;
    END
  END Tile_X0Y1_E2MID[5]
  PIN Tile_X0Y1_E2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.760 0.600 105.360 ;
    END
  END Tile_X0Y1_E2MID[6]
  PIN Tile_X0Y1_E2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.120 0.600 106.720 ;
    END
  END Tile_X0Y1_E2MID[7]
  PIN Tile_X0Y1_E6BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 140.120 225.000 140.720 ;
    END
  END Tile_X0Y1_E6BEG[0]
  PIN Tile_X0Y1_E6BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 153.720 225.000 154.320 ;
    END
  END Tile_X0Y1_E6BEG[10]
  PIN Tile_X0Y1_E6BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 155.080 225.000 155.680 ;
    END
  END Tile_X0Y1_E6BEG[11]
  PIN Tile_X0Y1_E6BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 141.480 225.000 142.080 ;
    END
  END Tile_X0Y1_E6BEG[1]
  PIN Tile_X0Y1_E6BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 142.840 225.000 143.440 ;
    END
  END Tile_X0Y1_E6BEG[2]
  PIN Tile_X0Y1_E6BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 144.200 225.000 144.800 ;
    END
  END Tile_X0Y1_E6BEG[3]
  PIN Tile_X0Y1_E6BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 145.560 225.000 146.160 ;
    END
  END Tile_X0Y1_E6BEG[4]
  PIN Tile_X0Y1_E6BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 146.920 225.000 147.520 ;
    END
  END Tile_X0Y1_E6BEG[5]
  PIN Tile_X0Y1_E6BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 148.280 225.000 148.880 ;
    END
  END Tile_X0Y1_E6BEG[6]
  PIN Tile_X0Y1_E6BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 149.640 225.000 150.240 ;
    END
  END Tile_X0Y1_E6BEG[7]
  PIN Tile_X0Y1_E6BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 151.000 225.000 151.600 ;
    END
  END Tile_X0Y1_E6BEG[8]
  PIN Tile_X0Y1_E6BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 152.360 225.000 152.960 ;
    END
  END Tile_X0Y1_E6BEG[9]
  PIN Tile_X0Y1_E6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.120 0.600 140.720 ;
    END
  END Tile_X0Y1_E6END[0]
  PIN Tile_X0Y1_E6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.720 0.600 154.320 ;
    END
  END Tile_X0Y1_E6END[10]
  PIN Tile_X0Y1_E6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.080 0.600 155.680 ;
    END
  END Tile_X0Y1_E6END[11]
  PIN Tile_X0Y1_E6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 141.480 0.600 142.080 ;
    END
  END Tile_X0Y1_E6END[1]
  PIN Tile_X0Y1_E6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 0.600 143.440 ;
    END
  END Tile_X0Y1_E6END[2]
  PIN Tile_X0Y1_E6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 144.200 0.600 144.800 ;
    END
  END Tile_X0Y1_E6END[3]
  PIN Tile_X0Y1_E6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 145.560 0.600 146.160 ;
    END
  END Tile_X0Y1_E6END[4]
  PIN Tile_X0Y1_E6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.920 0.600 147.520 ;
    END
  END Tile_X0Y1_E6END[5]
  PIN Tile_X0Y1_E6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.280 0.600 148.880 ;
    END
  END Tile_X0Y1_E6END[6]
  PIN Tile_X0Y1_E6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 0.600 150.240 ;
    END
  END Tile_X0Y1_E6END[7]
  PIN Tile_X0Y1_E6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.000 0.600 151.600 ;
    END
  END Tile_X0Y1_E6END[8]
  PIN Tile_X0Y1_E6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 152.360 0.600 152.960 ;
    END
  END Tile_X0Y1_E6END[9]
  PIN Tile_X0Y1_EE4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 118.360 225.000 118.960 ;
    END
  END Tile_X0Y1_EE4BEG[0]
  PIN Tile_X0Y1_EE4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 131.960 225.000 132.560 ;
    END
  END Tile_X0Y1_EE4BEG[10]
  PIN Tile_X0Y1_EE4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 133.320 225.000 133.920 ;
    END
  END Tile_X0Y1_EE4BEG[11]
  PIN Tile_X0Y1_EE4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 224.400 134.680 225.000 135.280 ;
    END
  END Tile_X0Y1_EE4BEG[12]
  PIN Tile_X0Y1_EE4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 224.400 136.040 225.000 136.640 ;
    END
  END Tile_X0Y1_EE4BEG[13]
  PIN Tile_X0Y1_EE4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 137.400 225.000 138.000 ;
    END
  END Tile_X0Y1_EE4BEG[14]
  PIN Tile_X0Y1_EE4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 224.400 138.760 225.000 139.360 ;
    END
  END Tile_X0Y1_EE4BEG[15]
  PIN Tile_X0Y1_EE4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 119.720 225.000 120.320 ;
    END
  END Tile_X0Y1_EE4BEG[1]
  PIN Tile_X0Y1_EE4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 121.080 225.000 121.680 ;
    END
  END Tile_X0Y1_EE4BEG[2]
  PIN Tile_X0Y1_EE4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 122.440 225.000 123.040 ;
    END
  END Tile_X0Y1_EE4BEG[3]
  PIN Tile_X0Y1_EE4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 123.800 225.000 124.400 ;
    END
  END Tile_X0Y1_EE4BEG[4]
  PIN Tile_X0Y1_EE4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 125.160 225.000 125.760 ;
    END
  END Tile_X0Y1_EE4BEG[5]
  PIN Tile_X0Y1_EE4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 126.520 225.000 127.120 ;
    END
  END Tile_X0Y1_EE4BEG[6]
  PIN Tile_X0Y1_EE4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 127.880 225.000 128.480 ;
    END
  END Tile_X0Y1_EE4BEG[7]
  PIN Tile_X0Y1_EE4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 129.240 225.000 129.840 ;
    END
  END Tile_X0Y1_EE4BEG[8]
  PIN Tile_X0Y1_EE4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 130.600 225.000 131.200 ;
    END
  END Tile_X0Y1_EE4BEG[9]
  PIN Tile_X0Y1_EE4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 118.360 0.600 118.960 ;
    END
  END Tile_X0Y1_EE4END[0]
  PIN Tile_X0Y1_EE4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.960 0.600 132.560 ;
    END
  END Tile_X0Y1_EE4END[10]
  PIN Tile_X0Y1_EE4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 133.320 0.600 133.920 ;
    END
  END Tile_X0Y1_EE4END[11]
  PIN Tile_X0Y1_EE4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.680 0.600 135.280 ;
    END
  END Tile_X0Y1_EE4END[12]
  PIN Tile_X0Y1_EE4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 0.600 136.640 ;
    END
  END Tile_X0Y1_EE4END[13]
  PIN Tile_X0Y1_EE4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 137.400 0.600 138.000 ;
    END
  END Tile_X0Y1_EE4END[14]
  PIN Tile_X0Y1_EE4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.760 0.600 139.360 ;
    END
  END Tile_X0Y1_EE4END[15]
  PIN Tile_X0Y1_EE4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.720 0.600 120.320 ;
    END
  END Tile_X0Y1_EE4END[1]
  PIN Tile_X0Y1_EE4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.080 0.600 121.680 ;
    END
  END Tile_X0Y1_EE4END[2]
  PIN Tile_X0Y1_EE4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 0.600 123.040 ;
    END
  END Tile_X0Y1_EE4END[3]
  PIN Tile_X0Y1_EE4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.800 0.600 124.400 ;
    END
  END Tile_X0Y1_EE4END[4]
  PIN Tile_X0Y1_EE4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.160 0.600 125.760 ;
    END
  END Tile_X0Y1_EE4END[5]
  PIN Tile_X0Y1_EE4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 126.520 0.600 127.120 ;
    END
  END Tile_X0Y1_EE4END[6]
  PIN Tile_X0Y1_EE4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.880 0.600 128.480 ;
    END
  END Tile_X0Y1_EE4END[7]
  PIN Tile_X0Y1_EE4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 0.600 129.840 ;
    END
  END Tile_X0Y1_EE4END[8]
  PIN Tile_X0Y1_EE4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 130.600 0.600 131.200 ;
    END
  END Tile_X0Y1_EE4END[9]
  PIN Tile_X0Y1_FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 0.600 157.040 ;
    END
  END Tile_X0Y1_FrameData[0]
  PIN Tile_X0Y1_FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 0.600 170.640 ;
    END
  END Tile_X0Y1_FrameData[10]
  PIN Tile_X0Y1_FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 171.400 0.600 172.000 ;
    END
  END Tile_X0Y1_FrameData[11]
  PIN Tile_X0Y1_FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.760 0.600 173.360 ;
    END
  END Tile_X0Y1_FrameData[12]
  PIN Tile_X0Y1_FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.120 0.600 174.720 ;
    END
  END Tile_X0Y1_FrameData[13]
  PIN Tile_X0Y1_FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 175.480 0.600 176.080 ;
    END
  END Tile_X0Y1_FrameData[14]
  PIN Tile_X0Y1_FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 0.600 177.440 ;
    END
  END Tile_X0Y1_FrameData[15]
  PIN Tile_X0Y1_FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.200 0.600 178.800 ;
    END
  END Tile_X0Y1_FrameData[16]
  PIN Tile_X0Y1_FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 179.560 0.600 180.160 ;
    END
  END Tile_X0Y1_FrameData[17]
  PIN Tile_X0Y1_FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.920 0.600 181.520 ;
    END
  END Tile_X0Y1_FrameData[18]
  PIN Tile_X0Y1_FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 182.280 0.600 182.880 ;
    END
  END Tile_X0Y1_FrameData[19]
  PIN Tile_X0Y1_FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 157.800 0.600 158.400 ;
    END
  END Tile_X0Y1_FrameData[1]
  PIN Tile_X0Y1_FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 0.600 184.240 ;
    END
  END Tile_X0Y1_FrameData[20]
  PIN Tile_X0Y1_FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.000 0.600 185.600 ;
    END
  END Tile_X0Y1_FrameData[21]
  PIN Tile_X0Y1_FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 186.360 0.600 186.960 ;
    END
  END Tile_X0Y1_FrameData[22]
  PIN Tile_X0Y1_FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.720 0.600 188.320 ;
    END
  END Tile_X0Y1_FrameData[23]
  PIN Tile_X0Y1_FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 189.080 0.600 189.680 ;
    END
  END Tile_X0Y1_FrameData[24]
  PIN Tile_X0Y1_FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.440 0.600 191.040 ;
    END
  END Tile_X0Y1_FrameData[25]
  PIN Tile_X0Y1_FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.800 0.600 192.400 ;
    END
  END Tile_X0Y1_FrameData[26]
  PIN Tile_X0Y1_FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.160 0.600 193.760 ;
    END
  END Tile_X0Y1_FrameData[27]
  PIN Tile_X0Y1_FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 194.520 0.600 195.120 ;
    END
  END Tile_X0Y1_FrameData[28]
  PIN Tile_X0Y1_FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 195.880 0.600 196.480 ;
    END
  END Tile_X0Y1_FrameData[29]
  PIN Tile_X0Y1_FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.160 0.600 159.760 ;
    END
  END Tile_X0Y1_FrameData[2]
  PIN Tile_X0Y1_FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.240 0.600 197.840 ;
    END
  END Tile_X0Y1_FrameData[30]
  PIN Tile_X0Y1_FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 198.600 0.600 199.200 ;
    END
  END Tile_X0Y1_FrameData[31]
  PIN Tile_X0Y1_FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 160.520 0.600 161.120 ;
    END
  END Tile_X0Y1_FrameData[3]
  PIN Tile_X0Y1_FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.880 0.600 162.480 ;
    END
  END Tile_X0Y1_FrameData[4]
  PIN Tile_X0Y1_FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 0.600 163.840 ;
    END
  END Tile_X0Y1_FrameData[5]
  PIN Tile_X0Y1_FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 164.600 0.600 165.200 ;
    END
  END Tile_X0Y1_FrameData[6]
  PIN Tile_X0Y1_FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.960 0.600 166.560 ;
    END
  END Tile_X0Y1_FrameData[7]
  PIN Tile_X0Y1_FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 167.320 0.600 167.920 ;
    END
  END Tile_X0Y1_FrameData[8]
  PIN Tile_X0Y1_FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.680 0.600 169.280 ;
    END
  END Tile_X0Y1_FrameData[9]
  PIN Tile_X0Y1_FrameData_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 156.440 225.000 157.040 ;
    END
  END Tile_X0Y1_FrameData_O[0]
  PIN Tile_X0Y1_FrameData_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 170.040 225.000 170.640 ;
    END
  END Tile_X0Y1_FrameData_O[10]
  PIN Tile_X0Y1_FrameData_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 171.400 225.000 172.000 ;
    END
  END Tile_X0Y1_FrameData_O[11]
  PIN Tile_X0Y1_FrameData_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 172.760 225.000 173.360 ;
    END
  END Tile_X0Y1_FrameData_O[12]
  PIN Tile_X0Y1_FrameData_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 174.120 225.000 174.720 ;
    END
  END Tile_X0Y1_FrameData_O[13]
  PIN Tile_X0Y1_FrameData_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 175.480 225.000 176.080 ;
    END
  END Tile_X0Y1_FrameData_O[14]
  PIN Tile_X0Y1_FrameData_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 176.840 225.000 177.440 ;
    END
  END Tile_X0Y1_FrameData_O[15]
  PIN Tile_X0Y1_FrameData_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 178.200 225.000 178.800 ;
    END
  END Tile_X0Y1_FrameData_O[16]
  PIN Tile_X0Y1_FrameData_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 179.560 225.000 180.160 ;
    END
  END Tile_X0Y1_FrameData_O[17]
  PIN Tile_X0Y1_FrameData_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 180.920 225.000 181.520 ;
    END
  END Tile_X0Y1_FrameData_O[18]
  PIN Tile_X0Y1_FrameData_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 182.280 225.000 182.880 ;
    END
  END Tile_X0Y1_FrameData_O[19]
  PIN Tile_X0Y1_FrameData_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 157.800 225.000 158.400 ;
    END
  END Tile_X0Y1_FrameData_O[1]
  PIN Tile_X0Y1_FrameData_O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 183.640 225.000 184.240 ;
    END
  END Tile_X0Y1_FrameData_O[20]
  PIN Tile_X0Y1_FrameData_O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 185.000 225.000 185.600 ;
    END
  END Tile_X0Y1_FrameData_O[21]
  PIN Tile_X0Y1_FrameData_O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 186.360 225.000 186.960 ;
    END
  END Tile_X0Y1_FrameData_O[22]
  PIN Tile_X0Y1_FrameData_O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 187.720 225.000 188.320 ;
    END
  END Tile_X0Y1_FrameData_O[23]
  PIN Tile_X0Y1_FrameData_O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 189.080 225.000 189.680 ;
    END
  END Tile_X0Y1_FrameData_O[24]
  PIN Tile_X0Y1_FrameData_O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 190.440 225.000 191.040 ;
    END
  END Tile_X0Y1_FrameData_O[25]
  PIN Tile_X0Y1_FrameData_O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 191.800 225.000 192.400 ;
    END
  END Tile_X0Y1_FrameData_O[26]
  PIN Tile_X0Y1_FrameData_O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 193.160 225.000 193.760 ;
    END
  END Tile_X0Y1_FrameData_O[27]
  PIN Tile_X0Y1_FrameData_O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 194.520 225.000 195.120 ;
    END
  END Tile_X0Y1_FrameData_O[28]
  PIN Tile_X0Y1_FrameData_O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 195.880 225.000 196.480 ;
    END
  END Tile_X0Y1_FrameData_O[29]
  PIN Tile_X0Y1_FrameData_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 159.160 225.000 159.760 ;
    END
  END Tile_X0Y1_FrameData_O[2]
  PIN Tile_X0Y1_FrameData_O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 197.240 225.000 197.840 ;
    END
  END Tile_X0Y1_FrameData_O[30]
  PIN Tile_X0Y1_FrameData_O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 198.600 225.000 199.200 ;
    END
  END Tile_X0Y1_FrameData_O[31]
  PIN Tile_X0Y1_FrameData_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 160.520 225.000 161.120 ;
    END
  END Tile_X0Y1_FrameData_O[3]
  PIN Tile_X0Y1_FrameData_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 161.880 225.000 162.480 ;
    END
  END Tile_X0Y1_FrameData_O[4]
  PIN Tile_X0Y1_FrameData_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 163.240 225.000 163.840 ;
    END
  END Tile_X0Y1_FrameData_O[5]
  PIN Tile_X0Y1_FrameData_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 164.600 225.000 165.200 ;
    END
  END Tile_X0Y1_FrameData_O[6]
  PIN Tile_X0Y1_FrameData_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 165.960 225.000 166.560 ;
    END
  END Tile_X0Y1_FrameData_O[7]
  PIN Tile_X0Y1_FrameData_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 167.320 225.000 167.920 ;
    END
  END Tile_X0Y1_FrameData_O[8]
  PIN Tile_X0Y1_FrameData_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 168.680 225.000 169.280 ;
    END
  END Tile_X0Y1_FrameData_O[9]
  PIN Tile_X0Y1_FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.295400 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 171.670 0.000 171.950 0.280 ;
    END
  END Tile_X0Y1_FrameStrobe[0]
  PIN Tile_X0Y1_FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.889100 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met2 ;
        RECT 185.470 0.000 185.750 0.280 ;
    END
  END Tile_X0Y1_FrameStrobe[10]
  PIN Tile_X0Y1_FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.241400 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 186.850 0.000 187.130 0.280 ;
    END
  END Tile_X0Y1_FrameStrobe[11]
  PIN Tile_X0Y1_FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.224900 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 188.230 0.000 188.510 0.280 ;
    END
  END Tile_X0Y1_FrameStrobe[12]
  PIN Tile_X0Y1_FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 189.610 0.000 189.890 0.280 ;
    END
  END Tile_X0Y1_FrameStrobe[13]
  PIN Tile_X0Y1_FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 190.990 0.000 191.270 0.280 ;
    END
  END Tile_X0Y1_FrameStrobe[14]
  PIN Tile_X0Y1_FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 192.370 0.000 192.650 0.280 ;
    END
  END Tile_X0Y1_FrameStrobe[15]
  PIN Tile_X0Y1_FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 193.750 0.000 194.030 0.280 ;
    END
  END Tile_X0Y1_FrameStrobe[16]
  PIN Tile_X0Y1_FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 195.130 0.000 195.410 0.280 ;
    END
  END Tile_X0Y1_FrameStrobe[17]
  PIN Tile_X0Y1_FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 196.510 0.000 196.790 0.280 ;
    END
  END Tile_X0Y1_FrameStrobe[18]
  PIN Tile_X0Y1_FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 197.890 0.000 198.170 0.280 ;
    END
  END Tile_X0Y1_FrameStrobe[19]
  PIN Tile_X0Y1_FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 173.050 0.000 173.330 0.280 ;
    END
  END Tile_X0Y1_FrameStrobe[1]
  PIN Tile_X0Y1_FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.585000 ;
    PORT
      LAYER met2 ;
        RECT 174.430 0.000 174.710 0.280 ;
    END
  END Tile_X0Y1_FrameStrobe[2]
  PIN Tile_X0Y1_FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 175.810 0.000 176.090 0.280 ;
    END
  END Tile_X0Y1_FrameStrobe[3]
  PIN Tile_X0Y1_FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.372000 ;
    PORT
      LAYER met2 ;
        RECT 177.190 0.000 177.470 0.280 ;
    END
  END Tile_X0Y1_FrameStrobe[4]
  PIN Tile_X0Y1_FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.711000 ;
    PORT
      LAYER met2 ;
        RECT 178.570 0.000 178.850 0.280 ;
    END
  END Tile_X0Y1_FrameStrobe[5]
  PIN Tile_X0Y1_FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 179.950 0.000 180.230 0.280 ;
    END
  END Tile_X0Y1_FrameStrobe[6]
  PIN Tile_X0Y1_FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.639000 ;
    PORT
      LAYER met2 ;
        RECT 181.330 0.000 181.610 0.280 ;
    END
  END Tile_X0Y1_FrameStrobe[7]
  PIN Tile_X0Y1_FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.241400 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 182.710 0.000 182.990 0.280 ;
    END
  END Tile_X0Y1_FrameStrobe[8]
  PIN Tile_X0Y1_FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.482800 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met2 ;
        RECT 184.090 0.000 184.370 0.280 ;
    END
  END Tile_X0Y1_FrameStrobe[9]
  PIN Tile_X0Y1_N1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 26.770 0.000 27.050 0.280 ;
    END
  END Tile_X0Y1_N1END[0]
  PIN Tile_X0Y1_N1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 28.150 0.000 28.430 0.280 ;
    END
  END Tile_X0Y1_N1END[1]
  PIN Tile_X0Y1_N1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 29.530 0.000 29.810 0.280 ;
    END
  END Tile_X0Y1_N1END[2]
  PIN Tile_X0Y1_N1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 30.910 0.000 31.190 0.280 ;
    END
  END Tile_X0Y1_N1END[3]
  PIN Tile_X0Y1_N2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 43.330 0.000 43.610 0.280 ;
    END
  END Tile_X0Y1_N2END[0]
  PIN Tile_X0Y1_N2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 44.710 0.000 44.990 0.280 ;
    END
  END Tile_X0Y1_N2END[1]
  PIN Tile_X0Y1_N2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 46.090 0.000 46.370 0.280 ;
    END
  END Tile_X0Y1_N2END[2]
  PIN Tile_X0Y1_N2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 47.470 0.000 47.750 0.280 ;
    END
  END Tile_X0Y1_N2END[3]
  PIN Tile_X0Y1_N2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 48.850 0.000 49.130 0.280 ;
    END
  END Tile_X0Y1_N2END[4]
  PIN Tile_X0Y1_N2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 50.230 0.000 50.510 0.280 ;
    END
  END Tile_X0Y1_N2END[5]
  PIN Tile_X0Y1_N2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 0.280 ;
    END
  END Tile_X0Y1_N2END[6]
  PIN Tile_X0Y1_N2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 52.990 0.000 53.270 0.280 ;
    END
  END Tile_X0Y1_N2END[7]
  PIN Tile_X0Y1_N2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 0.280 ;
    END
  END Tile_X0Y1_N2MID[0]
  PIN Tile_X0Y1_N2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 33.670 0.000 33.950 0.280 ;
    END
  END Tile_X0Y1_N2MID[1]
  PIN Tile_X0Y1_N2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 35.050 0.000 35.330 0.280 ;
    END
  END Tile_X0Y1_N2MID[2]
  PIN Tile_X0Y1_N2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 36.430 0.000 36.710 0.280 ;
    END
  END Tile_X0Y1_N2MID[3]
  PIN Tile_X0Y1_N2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 37.810 0.000 38.090 0.280 ;
    END
  END Tile_X0Y1_N2MID[4]
  PIN Tile_X0Y1_N2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 39.190 0.000 39.470 0.280 ;
    END
  END Tile_X0Y1_N2MID[5]
  PIN Tile_X0Y1_N2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 40.570 0.000 40.850 0.280 ;
    END
  END Tile_X0Y1_N2MID[6]
  PIN Tile_X0Y1_N2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 0.280 ;
    END
  END Tile_X0Y1_N2MID[7]
  PIN Tile_X0Y1_N4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 54.370 0.000 54.650 0.280 ;
    END
  END Tile_X0Y1_N4END[0]
  PIN Tile_X0Y1_N4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 68.170 0.000 68.450 0.280 ;
    END
  END Tile_X0Y1_N4END[10]
  PIN Tile_X0Y1_N4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 69.550 0.000 69.830 0.280 ;
    END
  END Tile_X0Y1_N4END[11]
  PIN Tile_X0Y1_N4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 0.280 ;
    END
  END Tile_X0Y1_N4END[12]
  PIN Tile_X0Y1_N4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 72.310 0.000 72.590 0.280 ;
    END
  END Tile_X0Y1_N4END[13]
  PIN Tile_X0Y1_N4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 73.690 0.000 73.970 0.280 ;
    END
  END Tile_X0Y1_N4END[14]
  PIN Tile_X0Y1_N4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 75.070 0.000 75.350 0.280 ;
    END
  END Tile_X0Y1_N4END[15]
  PIN Tile_X0Y1_N4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 55.750 0.000 56.030 0.280 ;
    END
  END Tile_X0Y1_N4END[1]
  PIN Tile_X0Y1_N4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 57.130 0.000 57.410 0.280 ;
    END
  END Tile_X0Y1_N4END[2]
  PIN Tile_X0Y1_N4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 58.510 0.000 58.790 0.280 ;
    END
  END Tile_X0Y1_N4END[3]
  PIN Tile_X0Y1_N4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 59.890 0.000 60.170 0.280 ;
    END
  END Tile_X0Y1_N4END[4]
  PIN Tile_X0Y1_N4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 0.280 ;
    END
  END Tile_X0Y1_N4END[5]
  PIN Tile_X0Y1_N4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 62.650 0.000 62.930 0.280 ;
    END
  END Tile_X0Y1_N4END[6]
  PIN Tile_X0Y1_N4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 64.030 0.000 64.310 0.280 ;
    END
  END Tile_X0Y1_N4END[7]
  PIN Tile_X0Y1_N4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.674100 ;
    ANTENNADIFFAREA 3.477600 ;
    PORT
      LAYER met2 ;
        RECT 65.410 0.000 65.690 0.280 ;
    END
  END Tile_X0Y1_N4END[8]
  PIN Tile_X0Y1_N4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.239400 ;
    ANTENNADIFFAREA 3.042900 ;
    PORT
      LAYER met2 ;
        RECT 66.790 0.000 67.070 0.280 ;
    END
  END Tile_X0Y1_N4END[9]
  PIN Tile_X0Y1_NN4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 76.450 0.000 76.730 0.280 ;
    END
  END Tile_X0Y1_NN4END[0]
  PIN Tile_X0Y1_NN4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 0.280 ;
    END
  END Tile_X0Y1_NN4END[10]
  PIN Tile_X0Y1_NN4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 91.630 0.000 91.910 0.280 ;
    END
  END Tile_X0Y1_NN4END[11]
  PIN Tile_X0Y1_NN4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 93.010 0.000 93.290 0.280 ;
    END
  END Tile_X0Y1_NN4END[12]
  PIN Tile_X0Y1_NN4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 94.390 0.000 94.670 0.280 ;
    END
  END Tile_X0Y1_NN4END[13]
  PIN Tile_X0Y1_NN4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 95.770 0.000 96.050 0.280 ;
    END
  END Tile_X0Y1_NN4END[14]
  PIN Tile_X0Y1_NN4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 97.150 0.000 97.430 0.280 ;
    END
  END Tile_X0Y1_NN4END[15]
  PIN Tile_X0Y1_NN4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 77.830 0.000 78.110 0.280 ;
    END
  END Tile_X0Y1_NN4END[1]
  PIN Tile_X0Y1_NN4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 79.210 0.000 79.490 0.280 ;
    END
  END Tile_X0Y1_NN4END[2]
  PIN Tile_X0Y1_NN4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 0.280 ;
    END
  END Tile_X0Y1_NN4END[3]
  PIN Tile_X0Y1_NN4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 81.970 0.000 82.250 0.280 ;
    END
  END Tile_X0Y1_NN4END[4]
  PIN Tile_X0Y1_NN4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 83.350 0.000 83.630 0.280 ;
    END
  END Tile_X0Y1_NN4END[5]
  PIN Tile_X0Y1_NN4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 84.730 0.000 85.010 0.280 ;
    END
  END Tile_X0Y1_NN4END[6]
  PIN Tile_X0Y1_NN4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 86.110 0.000 86.390 0.280 ;
    END
  END Tile_X0Y1_NN4END[7]
  PIN Tile_X0Y1_NN4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 87.490 0.000 87.770 0.280 ;
    END
  END Tile_X0Y1_NN4END[8]
  PIN Tile_X0Y1_NN4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 88.870 0.000 89.150 0.280 ;
    END
  END Tile_X0Y1_NN4END[9]
  PIN Tile_X0Y1_S1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 98.530 0.000 98.810 0.280 ;
    END
  END Tile_X0Y1_S1BEG[0]
  PIN Tile_X0Y1_S1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 0.280 ;
    END
  END Tile_X0Y1_S1BEG[1]
  PIN Tile_X0Y1_S1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 101.290 0.000 101.570 0.280 ;
    END
  END Tile_X0Y1_S1BEG[2]
  PIN Tile_X0Y1_S1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 102.670 0.000 102.950 0.280 ;
    END
  END Tile_X0Y1_S1BEG[3]
  PIN Tile_X0Y1_S2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 104.050 0.000 104.330 0.280 ;
    END
  END Tile_X0Y1_S2BEG[0]
  PIN Tile_X0Y1_S2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 105.430 0.000 105.710 0.280 ;
    END
  END Tile_X0Y1_S2BEG[1]
  PIN Tile_X0Y1_S2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 106.810 0.000 107.090 0.280 ;
    END
  END Tile_X0Y1_S2BEG[2]
  PIN Tile_X0Y1_S2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 108.190 0.000 108.470 0.280 ;
    END
  END Tile_X0Y1_S2BEG[3]
  PIN Tile_X0Y1_S2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 0.280 ;
    END
  END Tile_X0Y1_S2BEG[4]
  PIN Tile_X0Y1_S2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 110.950 0.000 111.230 0.280 ;
    END
  END Tile_X0Y1_S2BEG[5]
  PIN Tile_X0Y1_S2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 112.330 0.000 112.610 0.280 ;
    END
  END Tile_X0Y1_S2BEG[6]
  PIN Tile_X0Y1_S2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 113.710 0.000 113.990 0.280 ;
    END
  END Tile_X0Y1_S2BEG[7]
  PIN Tile_X0Y1_S2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 115.090 0.000 115.370 0.280 ;
    END
  END Tile_X0Y1_S2BEGb[0]
  PIN Tile_X0Y1_S2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 116.470 0.000 116.750 0.280 ;
    END
  END Tile_X0Y1_S2BEGb[1]
  PIN Tile_X0Y1_S2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 117.850 0.000 118.130 0.280 ;
    END
  END Tile_X0Y1_S2BEGb[2]
  PIN Tile_X0Y1_S2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 119.230 0.000 119.510 0.280 ;
    END
  END Tile_X0Y1_S2BEGb[3]
  PIN Tile_X0Y1_S2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 120.610 0.000 120.890 0.280 ;
    END
  END Tile_X0Y1_S2BEGb[4]
  PIN Tile_X0Y1_S2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 121.990 0.000 122.270 0.280 ;
    END
  END Tile_X0Y1_S2BEGb[5]
  PIN Tile_X0Y1_S2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 123.370 0.000 123.650 0.280 ;
    END
  END Tile_X0Y1_S2BEGb[6]
  PIN Tile_X0Y1_S2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 124.750 0.000 125.030 0.280 ;
    END
  END Tile_X0Y1_S2BEGb[7]
  PIN Tile_X0Y1_S4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 126.130 0.000 126.410 0.280 ;
    END
  END Tile_X0Y1_S4BEG[0]
  PIN Tile_X0Y1_S4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 139.930 0.000 140.210 0.280 ;
    END
  END Tile_X0Y1_S4BEG[10]
  PIN Tile_X0Y1_S4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 141.310 0.000 141.590 0.280 ;
    END
  END Tile_X0Y1_S4BEG[11]
  PIN Tile_X0Y1_S4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 142.690 0.000 142.970 0.280 ;
    END
  END Tile_X0Y1_S4BEG[12]
  PIN Tile_X0Y1_S4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 144.070 0.000 144.350 0.280 ;
    END
  END Tile_X0Y1_S4BEG[13]
  PIN Tile_X0Y1_S4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 145.450 0.000 145.730 0.280 ;
    END
  END Tile_X0Y1_S4BEG[14]
  PIN Tile_X0Y1_S4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 146.830 0.000 147.110 0.280 ;
    END
  END Tile_X0Y1_S4BEG[15]
  PIN Tile_X0Y1_S4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 127.510 0.000 127.790 0.280 ;
    END
  END Tile_X0Y1_S4BEG[1]
  PIN Tile_X0Y1_S4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 0.280 ;
    END
  END Tile_X0Y1_S4BEG[2]
  PIN Tile_X0Y1_S4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 130.270 0.000 130.550 0.280 ;
    END
  END Tile_X0Y1_S4BEG[3]
  PIN Tile_X0Y1_S4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 131.650 0.000 131.930 0.280 ;
    END
  END Tile_X0Y1_S4BEG[4]
  PIN Tile_X0Y1_S4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 133.030 0.000 133.310 0.280 ;
    END
  END Tile_X0Y1_S4BEG[5]
  PIN Tile_X0Y1_S4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 134.410 0.000 134.690 0.280 ;
    END
  END Tile_X0Y1_S4BEG[6]
  PIN Tile_X0Y1_S4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 135.790 0.000 136.070 0.280 ;
    END
  END Tile_X0Y1_S4BEG[7]
  PIN Tile_X0Y1_S4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 137.170 0.000 137.450 0.280 ;
    END
  END Tile_X0Y1_S4BEG[8]
  PIN Tile_X0Y1_S4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 138.550 0.000 138.830 0.280 ;
    END
  END Tile_X0Y1_S4BEG[9]
  PIN Tile_X0Y1_SS4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 148.210 0.000 148.490 0.280 ;
    END
  END Tile_X0Y1_SS4BEG[0]
  PIN Tile_X0Y1_SS4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 162.010 0.000 162.290 0.280 ;
    END
  END Tile_X0Y1_SS4BEG[10]
  PIN Tile_X0Y1_SS4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 163.390 0.000 163.670 0.280 ;
    END
  END Tile_X0Y1_SS4BEG[11]
  PIN Tile_X0Y1_SS4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 164.770 0.000 165.050 0.280 ;
    END
  END Tile_X0Y1_SS4BEG[12]
  PIN Tile_X0Y1_SS4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 166.150 0.000 166.430 0.280 ;
    END
  END Tile_X0Y1_SS4BEG[13]
  PIN Tile_X0Y1_SS4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 167.530 0.000 167.810 0.280 ;
    END
  END Tile_X0Y1_SS4BEG[14]
  PIN Tile_X0Y1_SS4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 168.910 0.000 169.190 0.280 ;
    END
  END Tile_X0Y1_SS4BEG[15]
  PIN Tile_X0Y1_SS4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 149.590 0.000 149.870 0.280 ;
    END
  END Tile_X0Y1_SS4BEG[1]
  PIN Tile_X0Y1_SS4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 150.970 0.000 151.250 0.280 ;
    END
  END Tile_X0Y1_SS4BEG[2]
  PIN Tile_X0Y1_SS4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 152.350 0.000 152.630 0.280 ;
    END
  END Tile_X0Y1_SS4BEG[3]
  PIN Tile_X0Y1_SS4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 153.730 0.000 154.010 0.280 ;
    END
  END Tile_X0Y1_SS4BEG[4]
  PIN Tile_X0Y1_SS4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 155.110 0.000 155.390 0.280 ;
    END
  END Tile_X0Y1_SS4BEG[5]
  PIN Tile_X0Y1_SS4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 156.490 0.000 156.770 0.280 ;
    END
  END Tile_X0Y1_SS4BEG[6]
  PIN Tile_X0Y1_SS4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 157.870 0.000 158.150 0.280 ;
    END
  END Tile_X0Y1_SS4BEG[7]
  PIN Tile_X0Y1_SS4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 159.250 0.000 159.530 0.280 ;
    END
  END Tile_X0Y1_SS4BEG[8]
  PIN Tile_X0Y1_SS4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 160.630 0.000 160.910 0.280 ;
    END
  END Tile_X0Y1_SS4BEG[9]
  PIN Tile_X0Y1_UserCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.704000 ;
    PORT
      LAYER met2 ;
        RECT 170.290 0.000 170.570 0.280 ;
    END
  END Tile_X0Y1_UserCLK
  PIN Tile_X0Y1_W1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.880 0.600 26.480 ;
    END
  END Tile_X0Y1_W1BEG[0]
  PIN Tile_X0Y1_W1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 0.600 27.840 ;
    END
  END Tile_X0Y1_W1BEG[1]
  PIN Tile_X0Y1_W1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 28.600 0.600 29.200 ;
    END
  END Tile_X0Y1_W1BEG[2]
  PIN Tile_X0Y1_W1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.960 0.600 30.560 ;
    END
  END Tile_X0Y1_W1BEG[3]
  PIN Tile_X0Y1_W1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 224.400 25.880 225.000 26.480 ;
    END
  END Tile_X0Y1_W1END[0]
  PIN Tile_X0Y1_W1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 27.240 225.000 27.840 ;
    END
  END Tile_X0Y1_W1END[1]
  PIN Tile_X0Y1_W1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 28.600 225.000 29.200 ;
    END
  END Tile_X0Y1_W1END[2]
  PIN Tile_X0Y1_W1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 29.960 225.000 30.560 ;
    END
  END Tile_X0Y1_W1END[3]
  PIN Tile_X0Y1_W2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 31.320 0.600 31.920 ;
    END
  END Tile_X0Y1_W2BEG[0]
  PIN Tile_X0Y1_W2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.680 0.600 33.280 ;
    END
  END Tile_X0Y1_W2BEG[1]
  PIN Tile_X0Y1_W2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 0.600 34.640 ;
    END
  END Tile_X0Y1_W2BEG[2]
  PIN Tile_X0Y1_W2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.400 0.600 36.000 ;
    END
  END Tile_X0Y1_W2BEG[3]
  PIN Tile_X0Y1_W2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.760 0.600 37.360 ;
    END
  END Tile_X0Y1_W2BEG[4]
  PIN Tile_X0Y1_W2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.120 0.600 38.720 ;
    END
  END Tile_X0Y1_W2BEG[5]
  PIN Tile_X0Y1_W2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.480 0.600 40.080 ;
    END
  END Tile_X0Y1_W2BEG[6]
  PIN Tile_X0Y1_W2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 0.600 41.440 ;
    END
  END Tile_X0Y1_W2BEG[7]
  PIN Tile_X0Y1_W2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.200 0.600 42.800 ;
    END
  END Tile_X0Y1_W2BEGb[0]
  PIN Tile_X0Y1_W2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.560 0.600 44.160 ;
    END
  END Tile_X0Y1_W2BEGb[1]
  PIN Tile_X0Y1_W2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.920 0.600 45.520 ;
    END
  END Tile_X0Y1_W2BEGb[2]
  PIN Tile_X0Y1_W2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.280 0.600 46.880 ;
    END
  END Tile_X0Y1_W2BEGb[3]
  PIN Tile_X0Y1_W2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 0.600 48.240 ;
    END
  END Tile_X0Y1_W2BEGb[4]
  PIN Tile_X0Y1_W2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.000 0.600 49.600 ;
    END
  END Tile_X0Y1_W2BEGb[5]
  PIN Tile_X0Y1_W2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 50.360 0.600 50.960 ;
    END
  END Tile_X0Y1_W2BEGb[6]
  PIN Tile_X0Y1_W2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.720 0.600 52.320 ;
    END
  END Tile_X0Y1_W2BEGb[7]
  PIN Tile_X0Y1_W2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 224.400 42.200 225.000 42.800 ;
    END
  END Tile_X0Y1_W2END[0]
  PIN Tile_X0Y1_W2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 224.400 43.560 225.000 44.160 ;
    END
  END Tile_X0Y1_W2END[1]
  PIN Tile_X0Y1_W2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 224.400 44.920 225.000 45.520 ;
    END
  END Tile_X0Y1_W2END[2]
  PIN Tile_X0Y1_W2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 224.400 46.280 225.000 46.880 ;
    END
  END Tile_X0Y1_W2END[3]
  PIN Tile_X0Y1_W2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 224.400 47.640 225.000 48.240 ;
    END
  END Tile_X0Y1_W2END[4]
  PIN Tile_X0Y1_W2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 224.400 49.000 225.000 49.600 ;
    END
  END Tile_X0Y1_W2END[5]
  PIN Tile_X0Y1_W2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 224.400 50.360 225.000 50.960 ;
    END
  END Tile_X0Y1_W2END[6]
  PIN Tile_X0Y1_W2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 224.400 51.720 225.000 52.320 ;
    END
  END Tile_X0Y1_W2END[7]
  PIN Tile_X0Y1_W2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 224.400 31.320 225.000 31.920 ;
    END
  END Tile_X0Y1_W2MID[0]
  PIN Tile_X0Y1_W2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 224.400 32.680 225.000 33.280 ;
    END
  END Tile_X0Y1_W2MID[1]
  PIN Tile_X0Y1_W2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 224.400 34.040 225.000 34.640 ;
    END
  END Tile_X0Y1_W2MID[2]
  PIN Tile_X0Y1_W2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 224.400 35.400 225.000 36.000 ;
    END
  END Tile_X0Y1_W2MID[3]
  PIN Tile_X0Y1_W2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 224.400 36.760 225.000 37.360 ;
    END
  END Tile_X0Y1_W2MID[4]
  PIN Tile_X0Y1_W2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 224.400 38.120 225.000 38.720 ;
    END
  END Tile_X0Y1_W2MID[5]
  PIN Tile_X0Y1_W2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 224.400 39.480 225.000 40.080 ;
    END
  END Tile_X0Y1_W2MID[6]
  PIN Tile_X0Y1_W2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 224.400 40.840 225.000 41.440 ;
    END
  END Tile_X0Y1_W2MID[7]
  PIN Tile_X0Y1_W6BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 0.600 75.440 ;
    END
  END Tile_X0Y1_W6BEG[0]
  PIN Tile_X0Y1_W6BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 0.600 89.040 ;
    END
  END Tile_X0Y1_W6BEG[10]
  PIN Tile_X0Y1_W6BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.800 0.600 90.400 ;
    END
  END Tile_X0Y1_W6BEG[11]
  PIN Tile_X0Y1_W6BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.200 0.600 76.800 ;
    END
  END Tile_X0Y1_W6BEG[1]
  PIN Tile_X0Y1_W6BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 77.560 0.600 78.160 ;
    END
  END Tile_X0Y1_W6BEG[2]
  PIN Tile_X0Y1_W6BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.920 0.600 79.520 ;
    END
  END Tile_X0Y1_W6BEG[3]
  PIN Tile_X0Y1_W6BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.280 0.600 80.880 ;
    END
  END Tile_X0Y1_W6BEG[4]
  PIN Tile_X0Y1_W6BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 0.600 82.240 ;
    END
  END Tile_X0Y1_W6BEG[5]
  PIN Tile_X0Y1_W6BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.000 0.600 83.600 ;
    END
  END Tile_X0Y1_W6BEG[6]
  PIN Tile_X0Y1_W6BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.360 0.600 84.960 ;
    END
  END Tile_X0Y1_W6BEG[7]
  PIN Tile_X0Y1_W6BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.720 0.600 86.320 ;
    END
  END Tile_X0Y1_W6BEG[8]
  PIN Tile_X0Y1_W6BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.080 0.600 87.680 ;
    END
  END Tile_X0Y1_W6BEG[9]
  PIN Tile_X0Y1_W6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 224.400 74.840 225.000 75.440 ;
    END
  END Tile_X0Y1_W6END[0]
  PIN Tile_X0Y1_W6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 88.440 225.000 89.040 ;
    END
  END Tile_X0Y1_W6END[10]
  PIN Tile_X0Y1_W6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 89.800 225.000 90.400 ;
    END
  END Tile_X0Y1_W6END[11]
  PIN Tile_X0Y1_W6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 224.400 76.200 225.000 76.800 ;
    END
  END Tile_X0Y1_W6END[1]
  PIN Tile_X0Y1_W6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 224.400 77.560 225.000 78.160 ;
    END
  END Tile_X0Y1_W6END[2]
  PIN Tile_X0Y1_W6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 224.400 78.920 225.000 79.520 ;
    END
  END Tile_X0Y1_W6END[3]
  PIN Tile_X0Y1_W6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 224.400 80.280 225.000 80.880 ;
    END
  END Tile_X0Y1_W6END[4]
  PIN Tile_X0Y1_W6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 224.400 81.640 225.000 82.240 ;
    END
  END Tile_X0Y1_W6END[5]
  PIN Tile_X0Y1_W6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 224.400 83.000 225.000 83.600 ;
    END
  END Tile_X0Y1_W6END[6]
  PIN Tile_X0Y1_W6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 224.400 84.360 225.000 84.960 ;
    END
  END Tile_X0Y1_W6END[7]
  PIN Tile_X0Y1_W6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 224.400 85.720 225.000 86.320 ;
    END
  END Tile_X0Y1_W6END[8]
  PIN Tile_X0Y1_W6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 224.400 87.080 225.000 87.680 ;
    END
  END Tile_X0Y1_W6END[9]
  PIN Tile_X0Y1_WW4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.080 0.600 53.680 ;
    END
  END Tile_X0Y1_WW4BEG[0]
  PIN Tile_X0Y1_WW4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.680 0.600 67.280 ;
    END
  END Tile_X0Y1_WW4BEG[10]
  PIN Tile_X0Y1_WW4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 0.600 68.640 ;
    END
  END Tile_X0Y1_WW4BEG[11]
  PIN Tile_X0Y1_WW4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.400 0.600 70.000 ;
    END
  END Tile_X0Y1_WW4BEG[12]
  PIN Tile_X0Y1_WW4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.760 0.600 71.360 ;
    END
  END Tile_X0Y1_WW4BEG[13]
  PIN Tile_X0Y1_WW4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.120 0.600 72.720 ;
    END
  END Tile_X0Y1_WW4BEG[14]
  PIN Tile_X0Y1_WW4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 73.480 0.600 74.080 ;
    END
  END Tile_X0Y1_WW4BEG[15]
  PIN Tile_X0Y1_WW4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 0.600 55.040 ;
    END
  END Tile_X0Y1_WW4BEG[1]
  PIN Tile_X0Y1_WW4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.800 0.600 56.400 ;
    END
  END Tile_X0Y1_WW4BEG[2]
  PIN Tile_X0Y1_WW4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.160 0.600 57.760 ;
    END
  END Tile_X0Y1_WW4BEG[3]
  PIN Tile_X0Y1_WW4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 58.520 0.600 59.120 ;
    END
  END Tile_X0Y1_WW4BEG[4]
  PIN Tile_X0Y1_WW4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.880 0.600 60.480 ;
    END
  END Tile_X0Y1_WW4BEG[5]
  PIN Tile_X0Y1_WW4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 0.600 61.840 ;
    END
  END Tile_X0Y1_WW4BEG[6]
  PIN Tile_X0Y1_WW4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.600 0.600 63.200 ;
    END
  END Tile_X0Y1_WW4BEG[7]
  PIN Tile_X0Y1_WW4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.960 0.600 64.560 ;
    END
  END Tile_X0Y1_WW4BEG[8]
  PIN Tile_X0Y1_WW4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 65.320 0.600 65.920 ;
    END
  END Tile_X0Y1_WW4BEG[9]
  PIN Tile_X0Y1_WW4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 224.400 53.080 225.000 53.680 ;
    END
  END Tile_X0Y1_WW4END[0]
  PIN Tile_X0Y1_WW4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 66.680 225.000 67.280 ;
    END
  END Tile_X0Y1_WW4END[10]
  PIN Tile_X0Y1_WW4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 68.040 225.000 68.640 ;
    END
  END Tile_X0Y1_WW4END[11]
  PIN Tile_X0Y1_WW4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 224.400 69.400 225.000 70.000 ;
    END
  END Tile_X0Y1_WW4END[12]
  PIN Tile_X0Y1_WW4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 224.400 70.760 225.000 71.360 ;
    END
  END Tile_X0Y1_WW4END[13]
  PIN Tile_X0Y1_WW4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 224.400 72.120 225.000 72.720 ;
    END
  END Tile_X0Y1_WW4END[14]
  PIN Tile_X0Y1_WW4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 224.400 73.480 225.000 74.080 ;
    END
  END Tile_X0Y1_WW4END[15]
  PIN Tile_X0Y1_WW4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 224.400 54.440 225.000 55.040 ;
    END
  END Tile_X0Y1_WW4END[1]
  PIN Tile_X0Y1_WW4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 224.400 55.800 225.000 56.400 ;
    END
  END Tile_X0Y1_WW4END[2]
  PIN Tile_X0Y1_WW4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 224.400 57.160 225.000 57.760 ;
    END
  END Tile_X0Y1_WW4END[3]
  PIN Tile_X0Y1_WW4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 58.520 225.000 59.120 ;
    END
  END Tile_X0Y1_WW4END[4]
  PIN Tile_X0Y1_WW4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 59.880 225.000 60.480 ;
    END
  END Tile_X0Y1_WW4END[5]
  PIN Tile_X0Y1_WW4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 61.240 225.000 61.840 ;
    END
  END Tile_X0Y1_WW4END[6]
  PIN Tile_X0Y1_WW4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 224.400 62.600 225.000 63.200 ;
    END
  END Tile_X0Y1_WW4END[7]
  PIN Tile_X0Y1_WW4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 224.400 63.960 225.000 64.560 ;
    END
  END Tile_X0Y1_WW4END[8]
  PIN Tile_X0Y1_WW4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 224.400 65.320 225.000 65.920 ;
    END
  END Tile_X0Y1_WW4END[9]
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 15.020 0.000 16.620 450.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 45.020 0.000 46.620 450.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 75.020 0.000 76.620 450.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 105.020 0.000 106.620 450.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 135.020 0.000 136.620 450.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 165.020 0.000 166.620 450.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 195.020 0.000 196.620 450.000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 9.720 0.000 11.320 450.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 39.720 0.000 41.320 450.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 69.720 0.000 71.320 450.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 99.720 0.000 101.320 450.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 129.720 0.000 131.320 450.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 159.720 0.000 161.320 450.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 189.720 0.000 191.320 450.000 ;
    END
  END VPWR
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 219.610 438.110 ;
      LAYER li1 ;
        RECT 5.520 10.795 219.420 438.005 ;
      LAYER met1 ;
        RECT 0.070 0.040 224.870 449.780 ;
      LAYER met2 ;
        RECT 0.090 449.440 26.490 449.890 ;
        RECT 27.330 449.440 27.870 449.890 ;
        RECT 28.710 449.440 29.250 449.890 ;
        RECT 30.090 449.440 30.630 449.890 ;
        RECT 31.470 449.440 32.010 449.890 ;
        RECT 32.850 449.440 33.390 449.890 ;
        RECT 34.230 449.440 34.770 449.890 ;
        RECT 35.610 449.440 36.150 449.890 ;
        RECT 36.990 449.440 37.530 449.890 ;
        RECT 38.370 449.440 38.910 449.890 ;
        RECT 39.750 449.440 40.290 449.890 ;
        RECT 41.130 449.440 41.670 449.890 ;
        RECT 42.510 449.440 43.050 449.890 ;
        RECT 43.890 449.440 44.430 449.890 ;
        RECT 45.270 449.440 45.810 449.890 ;
        RECT 46.650 449.440 47.190 449.890 ;
        RECT 48.030 449.440 48.570 449.890 ;
        RECT 49.410 449.440 49.950 449.890 ;
        RECT 50.790 449.440 51.330 449.890 ;
        RECT 52.170 449.440 52.710 449.890 ;
        RECT 53.550 449.440 54.090 449.890 ;
        RECT 54.930 449.440 55.470 449.890 ;
        RECT 56.310 449.440 56.850 449.890 ;
        RECT 57.690 449.440 58.230 449.890 ;
        RECT 59.070 449.440 59.610 449.890 ;
        RECT 60.450 449.440 60.990 449.890 ;
        RECT 61.830 449.440 62.370 449.890 ;
        RECT 63.210 449.440 63.750 449.890 ;
        RECT 64.590 449.440 65.130 449.890 ;
        RECT 65.970 449.440 66.510 449.890 ;
        RECT 67.350 449.440 67.890 449.890 ;
        RECT 68.730 449.440 69.270 449.890 ;
        RECT 70.110 449.440 70.650 449.890 ;
        RECT 71.490 449.440 72.030 449.890 ;
        RECT 72.870 449.440 73.410 449.890 ;
        RECT 74.250 449.440 74.790 449.890 ;
        RECT 75.630 449.440 76.170 449.890 ;
        RECT 77.010 449.440 77.550 449.890 ;
        RECT 78.390 449.440 78.930 449.890 ;
        RECT 79.770 449.440 80.310 449.890 ;
        RECT 81.150 449.440 81.690 449.890 ;
        RECT 82.530 449.440 83.070 449.890 ;
        RECT 83.910 449.440 84.450 449.890 ;
        RECT 85.290 449.440 85.830 449.890 ;
        RECT 86.670 449.440 87.210 449.890 ;
        RECT 88.050 449.440 88.590 449.890 ;
        RECT 89.430 449.440 89.970 449.890 ;
        RECT 90.810 449.440 91.350 449.890 ;
        RECT 92.190 449.440 92.730 449.890 ;
        RECT 93.570 449.440 94.110 449.890 ;
        RECT 94.950 449.440 95.490 449.890 ;
        RECT 96.330 449.440 96.870 449.890 ;
        RECT 97.710 449.440 98.250 449.890 ;
        RECT 99.090 449.440 99.630 449.890 ;
        RECT 100.470 449.440 101.010 449.890 ;
        RECT 101.850 449.440 102.390 449.890 ;
        RECT 103.230 449.440 103.770 449.890 ;
        RECT 104.610 449.440 105.150 449.890 ;
        RECT 105.990 449.440 106.530 449.890 ;
        RECT 107.370 449.440 107.910 449.890 ;
        RECT 108.750 449.440 109.290 449.890 ;
        RECT 110.130 449.440 110.670 449.890 ;
        RECT 111.510 449.440 112.050 449.890 ;
        RECT 112.890 449.440 113.430 449.890 ;
        RECT 114.270 449.440 114.810 449.890 ;
        RECT 115.650 449.440 116.190 449.890 ;
        RECT 117.030 449.440 117.570 449.890 ;
        RECT 118.410 449.440 118.950 449.890 ;
        RECT 119.790 449.440 120.330 449.890 ;
        RECT 121.170 449.440 121.710 449.890 ;
        RECT 122.550 449.440 123.090 449.890 ;
        RECT 123.930 449.440 124.470 449.890 ;
        RECT 125.310 449.440 125.850 449.890 ;
        RECT 126.690 449.440 127.230 449.890 ;
        RECT 128.070 449.440 128.610 449.890 ;
        RECT 129.450 449.440 129.990 449.890 ;
        RECT 130.830 449.440 131.370 449.890 ;
        RECT 132.210 449.440 132.750 449.890 ;
        RECT 133.590 449.440 134.130 449.890 ;
        RECT 134.970 449.440 135.510 449.890 ;
        RECT 136.350 449.440 136.890 449.890 ;
        RECT 137.730 449.440 138.270 449.890 ;
        RECT 139.110 449.440 139.650 449.890 ;
        RECT 140.490 449.440 141.030 449.890 ;
        RECT 141.870 449.440 142.410 449.890 ;
        RECT 143.250 449.440 143.790 449.890 ;
        RECT 144.630 449.440 145.170 449.890 ;
        RECT 146.010 449.440 146.550 449.890 ;
        RECT 147.390 449.440 147.930 449.890 ;
        RECT 148.770 449.440 149.310 449.890 ;
        RECT 150.150 449.440 150.690 449.890 ;
        RECT 151.530 449.440 152.070 449.890 ;
        RECT 152.910 449.440 153.450 449.890 ;
        RECT 154.290 449.440 154.830 449.890 ;
        RECT 155.670 449.440 156.210 449.890 ;
        RECT 157.050 449.440 157.590 449.890 ;
        RECT 158.430 449.440 158.970 449.890 ;
        RECT 159.810 449.440 160.350 449.890 ;
        RECT 161.190 449.440 161.730 449.890 ;
        RECT 162.570 449.440 163.110 449.890 ;
        RECT 163.950 449.440 164.490 449.890 ;
        RECT 165.330 449.440 165.870 449.890 ;
        RECT 166.710 449.440 167.250 449.890 ;
        RECT 168.090 449.440 168.630 449.890 ;
        RECT 169.470 449.440 170.010 449.890 ;
        RECT 170.850 449.440 171.390 449.890 ;
        RECT 172.230 449.440 172.770 449.890 ;
        RECT 173.610 449.440 174.150 449.890 ;
        RECT 174.990 449.440 175.530 449.890 ;
        RECT 176.370 449.440 176.910 449.890 ;
        RECT 177.750 449.440 178.290 449.890 ;
        RECT 179.130 449.440 179.670 449.890 ;
        RECT 180.510 449.440 181.050 449.890 ;
        RECT 181.890 449.440 182.430 449.890 ;
        RECT 183.270 449.440 183.810 449.890 ;
        RECT 184.650 449.440 185.190 449.890 ;
        RECT 186.030 449.440 186.570 449.890 ;
        RECT 187.410 449.440 187.950 449.890 ;
        RECT 188.790 449.440 189.330 449.890 ;
        RECT 190.170 449.440 190.710 449.890 ;
        RECT 191.550 449.440 192.090 449.890 ;
        RECT 192.930 449.440 193.470 449.890 ;
        RECT 194.310 449.440 194.850 449.890 ;
        RECT 195.690 449.440 196.230 449.890 ;
        RECT 197.070 449.440 197.610 449.890 ;
        RECT 198.450 449.440 224.840 449.890 ;
        RECT 0.090 0.560 224.840 449.440 ;
        RECT 0.090 0.010 26.490 0.560 ;
        RECT 27.330 0.010 27.870 0.560 ;
        RECT 28.710 0.010 29.250 0.560 ;
        RECT 30.090 0.010 30.630 0.560 ;
        RECT 31.470 0.010 32.010 0.560 ;
        RECT 32.850 0.010 33.390 0.560 ;
        RECT 34.230 0.010 34.770 0.560 ;
        RECT 35.610 0.010 36.150 0.560 ;
        RECT 36.990 0.010 37.530 0.560 ;
        RECT 38.370 0.010 38.910 0.560 ;
        RECT 39.750 0.010 40.290 0.560 ;
        RECT 41.130 0.010 41.670 0.560 ;
        RECT 42.510 0.010 43.050 0.560 ;
        RECT 43.890 0.010 44.430 0.560 ;
        RECT 45.270 0.010 45.810 0.560 ;
        RECT 46.650 0.010 47.190 0.560 ;
        RECT 48.030 0.010 48.570 0.560 ;
        RECT 49.410 0.010 49.950 0.560 ;
        RECT 50.790 0.010 51.330 0.560 ;
        RECT 52.170 0.010 52.710 0.560 ;
        RECT 53.550 0.010 54.090 0.560 ;
        RECT 54.930 0.010 55.470 0.560 ;
        RECT 56.310 0.010 56.850 0.560 ;
        RECT 57.690 0.010 58.230 0.560 ;
        RECT 59.070 0.010 59.610 0.560 ;
        RECT 60.450 0.010 60.990 0.560 ;
        RECT 61.830 0.010 62.370 0.560 ;
        RECT 63.210 0.010 63.750 0.560 ;
        RECT 64.590 0.010 65.130 0.560 ;
        RECT 65.970 0.010 66.510 0.560 ;
        RECT 67.350 0.010 67.890 0.560 ;
        RECT 68.730 0.010 69.270 0.560 ;
        RECT 70.110 0.010 70.650 0.560 ;
        RECT 71.490 0.010 72.030 0.560 ;
        RECT 72.870 0.010 73.410 0.560 ;
        RECT 74.250 0.010 74.790 0.560 ;
        RECT 75.630 0.010 76.170 0.560 ;
        RECT 77.010 0.010 77.550 0.560 ;
        RECT 78.390 0.010 78.930 0.560 ;
        RECT 79.770 0.010 80.310 0.560 ;
        RECT 81.150 0.010 81.690 0.560 ;
        RECT 82.530 0.010 83.070 0.560 ;
        RECT 83.910 0.010 84.450 0.560 ;
        RECT 85.290 0.010 85.830 0.560 ;
        RECT 86.670 0.010 87.210 0.560 ;
        RECT 88.050 0.010 88.590 0.560 ;
        RECT 89.430 0.010 89.970 0.560 ;
        RECT 90.810 0.010 91.350 0.560 ;
        RECT 92.190 0.010 92.730 0.560 ;
        RECT 93.570 0.010 94.110 0.560 ;
        RECT 94.950 0.010 95.490 0.560 ;
        RECT 96.330 0.010 96.870 0.560 ;
        RECT 97.710 0.010 98.250 0.560 ;
        RECT 99.090 0.010 99.630 0.560 ;
        RECT 100.470 0.010 101.010 0.560 ;
        RECT 101.850 0.010 102.390 0.560 ;
        RECT 103.230 0.010 103.770 0.560 ;
        RECT 104.610 0.010 105.150 0.560 ;
        RECT 105.990 0.010 106.530 0.560 ;
        RECT 107.370 0.010 107.910 0.560 ;
        RECT 108.750 0.010 109.290 0.560 ;
        RECT 110.130 0.010 110.670 0.560 ;
        RECT 111.510 0.010 112.050 0.560 ;
        RECT 112.890 0.010 113.430 0.560 ;
        RECT 114.270 0.010 114.810 0.560 ;
        RECT 115.650 0.010 116.190 0.560 ;
        RECT 117.030 0.010 117.570 0.560 ;
        RECT 118.410 0.010 118.950 0.560 ;
        RECT 119.790 0.010 120.330 0.560 ;
        RECT 121.170 0.010 121.710 0.560 ;
        RECT 122.550 0.010 123.090 0.560 ;
        RECT 123.930 0.010 124.470 0.560 ;
        RECT 125.310 0.010 125.850 0.560 ;
        RECT 126.690 0.010 127.230 0.560 ;
        RECT 128.070 0.010 128.610 0.560 ;
        RECT 129.450 0.010 129.990 0.560 ;
        RECT 130.830 0.010 131.370 0.560 ;
        RECT 132.210 0.010 132.750 0.560 ;
        RECT 133.590 0.010 134.130 0.560 ;
        RECT 134.970 0.010 135.510 0.560 ;
        RECT 136.350 0.010 136.890 0.560 ;
        RECT 137.730 0.010 138.270 0.560 ;
        RECT 139.110 0.010 139.650 0.560 ;
        RECT 140.490 0.010 141.030 0.560 ;
        RECT 141.870 0.010 142.410 0.560 ;
        RECT 143.250 0.010 143.790 0.560 ;
        RECT 144.630 0.010 145.170 0.560 ;
        RECT 146.010 0.010 146.550 0.560 ;
        RECT 147.390 0.010 147.930 0.560 ;
        RECT 148.770 0.010 149.310 0.560 ;
        RECT 150.150 0.010 150.690 0.560 ;
        RECT 151.530 0.010 152.070 0.560 ;
        RECT 152.910 0.010 153.450 0.560 ;
        RECT 154.290 0.010 154.830 0.560 ;
        RECT 155.670 0.010 156.210 0.560 ;
        RECT 157.050 0.010 157.590 0.560 ;
        RECT 158.430 0.010 158.970 0.560 ;
        RECT 159.810 0.010 160.350 0.560 ;
        RECT 161.190 0.010 161.730 0.560 ;
        RECT 162.570 0.010 163.110 0.560 ;
        RECT 163.950 0.010 164.490 0.560 ;
        RECT 165.330 0.010 165.870 0.560 ;
        RECT 166.710 0.010 167.250 0.560 ;
        RECT 168.090 0.010 168.630 0.560 ;
        RECT 169.470 0.010 170.010 0.560 ;
        RECT 170.850 0.010 171.390 0.560 ;
        RECT 172.230 0.010 172.770 0.560 ;
        RECT 173.610 0.010 174.150 0.560 ;
        RECT 174.990 0.010 175.530 0.560 ;
        RECT 176.370 0.010 176.910 0.560 ;
        RECT 177.750 0.010 178.290 0.560 ;
        RECT 179.130 0.010 179.670 0.560 ;
        RECT 180.510 0.010 181.050 0.560 ;
        RECT 181.890 0.010 182.430 0.560 ;
        RECT 183.270 0.010 183.810 0.560 ;
        RECT 184.650 0.010 185.190 0.560 ;
        RECT 186.030 0.010 186.570 0.560 ;
        RECT 187.410 0.010 187.950 0.560 ;
        RECT 188.790 0.010 189.330 0.560 ;
        RECT 190.170 0.010 190.710 0.560 ;
        RECT 191.550 0.010 192.090 0.560 ;
        RECT 192.930 0.010 193.470 0.560 ;
        RECT 194.310 0.010 194.850 0.560 ;
        RECT 195.690 0.010 196.230 0.560 ;
        RECT 197.070 0.010 197.610 0.560 ;
        RECT 198.450 0.010 224.840 0.560 ;
      LAYER met3 ;
        RECT 0.065 424.600 224.400 443.865 ;
        RECT 1.000 250.480 224.000 424.600 ;
        RECT 0.065 199.600 224.400 250.480 ;
        RECT 1.000 25.480 224.000 199.600 ;
        RECT 0.065 0.175 224.400 25.480 ;
      LAYER met4 ;
        RECT 1.215 0.175 9.320 443.865 ;
        RECT 11.720 0.175 14.620 443.865 ;
        RECT 17.020 0.175 39.320 443.865 ;
        RECT 41.720 0.175 44.620 443.865 ;
        RECT 47.020 0.175 69.320 443.865 ;
        RECT 71.720 0.175 74.620 443.865 ;
        RECT 77.020 0.175 99.320 443.865 ;
        RECT 101.720 0.175 104.620 443.865 ;
        RECT 107.020 0.175 129.320 443.865 ;
        RECT 131.720 0.175 134.620 443.865 ;
        RECT 137.020 0.175 159.320 443.865 ;
        RECT 161.720 0.175 164.620 443.865 ;
        RECT 167.020 0.175 189.320 443.865 ;
        RECT 191.720 0.175 194.620 443.865 ;
        RECT 197.020 0.175 224.170 443.865 ;
  END
END DSP
END LIBRARY

