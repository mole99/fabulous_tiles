* NGSPICE file created from IHP_SRAM.ext - technology: ihp-sg13g2

* Black-box entry subcircuit for sg13g2_mux4_1 abstract view
.subckt sg13g2_mux4_1 S0 A0 A1 A2 A3 S1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_1 abstract view
.subckt sg13g2_inv_1 VDD Y A VSS
.ends

* Black-box entry subcircuit for sg13g2_decap_8 abstract view
.subckt sg13g2_decap_8 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_1 abstract view
.subckt sg13g2_fill_1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dlhq_1 abstract view
.subckt sg13g2_dlhq_1 D GATE Q VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_1 abstract view
.subckt sg13g2_buf_1 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21oi_1 abstract view
.subckt sg13g2_a21oi_1 VSS VDD A1 A2 Y B1
.ends

* Black-box entry subcircuit for sg13g2_fill_2 abstract view
.subckt sg13g2_fill_2 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_decap_4 abstract view
.subckt sg13g2_decap_4 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2b_1 abstract view
.subckt sg13g2_nand2b_1 Y B A_N VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_o21ai_1 abstract view
.subckt sg13g2_o21ai_1 B1 VDD Y VSS A1 A2
.ends

* Black-box entry subcircuit for sg13g2_mux2_1 abstract view
.subckt sg13g2_mux2_1 A0 A1 S X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2b_1 abstract view
.subckt sg13g2_nor2b_1 A B_N Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2_1 abstract view
.subckt sg13g2_nor2_1 A B Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor3_1 abstract view
.subckt sg13g2_nor3_1 A B C Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2_1 abstract view
.subckt sg13g2_nand2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_tielo abstract view
.subckt sg13g2_tielo VDD VSS L_LO
.ends

* Black-box entry subcircuit for sg13g2_a221oi_1 abstract view
.subckt sg13g2_a221oi_1 VSS VDD B2 C1 B1 A1 Y A2
.ends

* Black-box entry subcircuit for sg13g2_nand3_1 abstract view
.subckt sg13g2_nand3_1 B C A Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand3b_1 abstract view
.subckt sg13g2_nand3b_1 B C Y VDD VSS A_N
.ends

* Black-box entry subcircuit for sg13g2_tiehi abstract view
.subckt sg13g2_tiehi VDD VSS L_HI
.ends

* Black-box entry subcircuit for sg13g2_a22oi_1 abstract view
.subckt sg13g2_a22oi_1 Y B1 B2 A2 A1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand4_1 abstract view
.subckt sg13g2_nand4_1 B C A Y VDD VSS D
.ends

* Black-box entry subcircuit for sg13g2_or2_1 abstract view
.subckt sg13g2_or2_1 VSS VDD X B A
.ends

* Black-box entry subcircuit for sg13g2_or3_1 abstract view
.subckt sg13g2_or3_1 A B C X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and2_1 abstract view
.subckt sg13g2_and2_1 A B X VDD VSS
.ends

.subckt IHP_SRAM ADDR_SRAM0 ADDR_SRAM1 ADDR_SRAM2 ADDR_SRAM3 ADDR_SRAM4 ADDR_SRAM5
+ ADDR_SRAM6 ADDR_SRAM7 ADDR_SRAM8 ADDR_SRAM9 BM_SRAM0 BM_SRAM1 BM_SRAM10 BM_SRAM11
+ BM_SRAM12 BM_SRAM13 BM_SRAM14 BM_SRAM15 BM_SRAM16 BM_SRAM17 BM_SRAM18 BM_SRAM19
+ BM_SRAM2 BM_SRAM20 BM_SRAM21 BM_SRAM22 BM_SRAM23 BM_SRAM24 BM_SRAM25 BM_SRAM26 BM_SRAM27
+ BM_SRAM28 BM_SRAM29 BM_SRAM3 BM_SRAM30 BM_SRAM31 BM_SRAM4 BM_SRAM5 BM_SRAM6 BM_SRAM7
+ BM_SRAM8 BM_SRAM9 CLK_SRAM CONFIGURED_top DIN_SRAM0 DIN_SRAM1 DIN_SRAM10 DIN_SRAM11
+ DIN_SRAM12 DIN_SRAM13 DIN_SRAM14 DIN_SRAM15 DIN_SRAM16 DIN_SRAM17 DIN_SRAM18 DIN_SRAM19
+ DIN_SRAM2 DIN_SRAM20 DIN_SRAM21 DIN_SRAM22 DIN_SRAM23 DIN_SRAM24 DIN_SRAM25 DIN_SRAM26
+ DIN_SRAM27 DIN_SRAM28 DIN_SRAM29 DIN_SRAM3 DIN_SRAM30 DIN_SRAM31 DIN_SRAM4 DIN_SRAM5
+ DIN_SRAM6 DIN_SRAM7 DIN_SRAM8 DIN_SRAM9 DOUT_SRAM0 DOUT_SRAM1 DOUT_SRAM10 DOUT_SRAM11
+ DOUT_SRAM12 DOUT_SRAM13 DOUT_SRAM14 DOUT_SRAM15 DOUT_SRAM16 DOUT_SRAM17 DOUT_SRAM18
+ DOUT_SRAM19 DOUT_SRAM2 DOUT_SRAM20 DOUT_SRAM21 DOUT_SRAM22 DOUT_SRAM23 DOUT_SRAM24
+ DOUT_SRAM25 DOUT_SRAM26 DOUT_SRAM27 DOUT_SRAM28 DOUT_SRAM29 DOUT_SRAM3 DOUT_SRAM30
+ DOUT_SRAM31 DOUT_SRAM4 DOUT_SRAM5 DOUT_SRAM6 DOUT_SRAM7 DOUT_SRAM8 DOUT_SRAM9 MEN_SRAM
+ REN_SRAM TIE_HIGH_SRAM TIE_LOW_SRAM Tile_X0Y0_E1END[0] Tile_X0Y0_E1END[1] Tile_X0Y0_E1END[2]
+ Tile_X0Y0_E1END[3] Tile_X0Y0_E2END[0] Tile_X0Y0_E2END[1] Tile_X0Y0_E2END[2] Tile_X0Y0_E2END[3]
+ Tile_X0Y0_E2END[4] Tile_X0Y0_E2END[5] Tile_X0Y0_E2END[6] Tile_X0Y0_E2END[7] Tile_X0Y0_E2MID[0]
+ Tile_X0Y0_E2MID[1] Tile_X0Y0_E2MID[2] Tile_X0Y0_E2MID[3] Tile_X0Y0_E2MID[4] Tile_X0Y0_E2MID[5]
+ Tile_X0Y0_E2MID[6] Tile_X0Y0_E2MID[7] Tile_X0Y0_E6END[0] Tile_X0Y0_E6END[10] Tile_X0Y0_E6END[11]
+ Tile_X0Y0_E6END[1] Tile_X0Y0_E6END[2] Tile_X0Y0_E6END[3] Tile_X0Y0_E6END[4] Tile_X0Y0_E6END[5]
+ Tile_X0Y0_E6END[6] Tile_X0Y0_E6END[7] Tile_X0Y0_E6END[8] Tile_X0Y0_E6END[9] Tile_X0Y0_EE4END[0]
+ Tile_X0Y0_EE4END[10] Tile_X0Y0_EE4END[11] Tile_X0Y0_EE4END[12] Tile_X0Y0_EE4END[13]
+ Tile_X0Y0_EE4END[14] Tile_X0Y0_EE4END[15] Tile_X0Y0_EE4END[1] Tile_X0Y0_EE4END[2]
+ Tile_X0Y0_EE4END[3] Tile_X0Y0_EE4END[4] Tile_X0Y0_EE4END[5] Tile_X0Y0_EE4END[6]
+ Tile_X0Y0_EE4END[7] Tile_X0Y0_EE4END[8] Tile_X0Y0_EE4END[9] Tile_X0Y0_FrameData[0]
+ Tile_X0Y0_FrameData[10] Tile_X0Y0_FrameData[11] Tile_X0Y0_FrameData[12] Tile_X0Y0_FrameData[13]
+ Tile_X0Y0_FrameData[14] Tile_X0Y0_FrameData[15] Tile_X0Y0_FrameData[16] Tile_X0Y0_FrameData[17]
+ Tile_X0Y0_FrameData[18] Tile_X0Y0_FrameData[19] Tile_X0Y0_FrameData[1] Tile_X0Y0_FrameData[20]
+ Tile_X0Y0_FrameData[21] Tile_X0Y0_FrameData[22] Tile_X0Y0_FrameData[23] Tile_X0Y0_FrameData[24]
+ Tile_X0Y0_FrameData[25] Tile_X0Y0_FrameData[26] Tile_X0Y0_FrameData[27] Tile_X0Y0_FrameData[28]
+ Tile_X0Y0_FrameData[29] Tile_X0Y0_FrameData[2] Tile_X0Y0_FrameData[30] Tile_X0Y0_FrameData[31]
+ Tile_X0Y0_FrameData[3] Tile_X0Y0_FrameData[4] Tile_X0Y0_FrameData[5] Tile_X0Y0_FrameData[6]
+ Tile_X0Y0_FrameData[7] Tile_X0Y0_FrameData[8] Tile_X0Y0_FrameData[9] Tile_X0Y0_FrameData_O[0]
+ Tile_X0Y0_FrameData_O[10] Tile_X0Y0_FrameData_O[11] Tile_X0Y0_FrameData_O[12] Tile_X0Y0_FrameData_O[13]
+ Tile_X0Y0_FrameData_O[14] Tile_X0Y0_FrameData_O[15] Tile_X0Y0_FrameData_O[16] Tile_X0Y0_FrameData_O[17]
+ Tile_X0Y0_FrameData_O[18] Tile_X0Y0_FrameData_O[19] Tile_X0Y0_FrameData_O[1] Tile_X0Y0_FrameData_O[20]
+ Tile_X0Y0_FrameData_O[21] Tile_X0Y0_FrameData_O[22] Tile_X0Y0_FrameData_O[23] Tile_X0Y0_FrameData_O[24]
+ Tile_X0Y0_FrameData_O[25] Tile_X0Y0_FrameData_O[26] Tile_X0Y0_FrameData_O[27] Tile_X0Y0_FrameData_O[28]
+ Tile_X0Y0_FrameData_O[29] Tile_X0Y0_FrameData_O[2] Tile_X0Y0_FrameData_O[30] Tile_X0Y0_FrameData_O[31]
+ Tile_X0Y0_FrameData_O[3] Tile_X0Y0_FrameData_O[4] Tile_X0Y0_FrameData_O[5] Tile_X0Y0_FrameData_O[6]
+ Tile_X0Y0_FrameData_O[7] Tile_X0Y0_FrameData_O[8] Tile_X0Y0_FrameData_O[9] Tile_X0Y0_FrameStrobe_O[0]
+ Tile_X0Y0_FrameStrobe_O[10] Tile_X0Y0_FrameStrobe_O[11] Tile_X0Y0_FrameStrobe_O[12]
+ Tile_X0Y0_FrameStrobe_O[13] Tile_X0Y0_FrameStrobe_O[14] Tile_X0Y0_FrameStrobe_O[15]
+ Tile_X0Y0_FrameStrobe_O[16] Tile_X0Y0_FrameStrobe_O[17] Tile_X0Y0_FrameStrobe_O[18]
+ Tile_X0Y0_FrameStrobe_O[19] Tile_X0Y0_FrameStrobe_O[1] Tile_X0Y0_FrameStrobe_O[2]
+ Tile_X0Y0_FrameStrobe_O[3] Tile_X0Y0_FrameStrobe_O[4] Tile_X0Y0_FrameStrobe_O[5]
+ Tile_X0Y0_FrameStrobe_O[6] Tile_X0Y0_FrameStrobe_O[7] Tile_X0Y0_FrameStrobe_O[8]
+ Tile_X0Y0_FrameStrobe_O[9] Tile_X0Y0_N1BEG[0] Tile_X0Y0_N1BEG[1] Tile_X0Y0_N1BEG[2]
+ Tile_X0Y0_N1BEG[3] Tile_X0Y0_N2BEG[0] Tile_X0Y0_N2BEG[1] Tile_X0Y0_N2BEG[2] Tile_X0Y0_N2BEG[3]
+ Tile_X0Y0_N2BEG[4] Tile_X0Y0_N2BEG[5] Tile_X0Y0_N2BEG[6] Tile_X0Y0_N2BEG[7] Tile_X0Y0_N2BEGb[0]
+ Tile_X0Y0_N2BEGb[1] Tile_X0Y0_N2BEGb[2] Tile_X0Y0_N2BEGb[3] Tile_X0Y0_N2BEGb[4]
+ Tile_X0Y0_N2BEGb[5] Tile_X0Y0_N2BEGb[6] Tile_X0Y0_N2BEGb[7] Tile_X0Y0_N4BEG[0] Tile_X0Y0_N4BEG[10]
+ Tile_X0Y0_N4BEG[11] Tile_X0Y0_N4BEG[12] Tile_X0Y0_N4BEG[13] Tile_X0Y0_N4BEG[14]
+ Tile_X0Y0_N4BEG[15] Tile_X0Y0_N4BEG[1] Tile_X0Y0_N4BEG[2] Tile_X0Y0_N4BEG[3] Tile_X0Y0_N4BEG[4]
+ Tile_X0Y0_N4BEG[5] Tile_X0Y0_N4BEG[6] Tile_X0Y0_N4BEG[7] Tile_X0Y0_N4BEG[8] Tile_X0Y0_N4BEG[9]
+ Tile_X0Y0_S1END[0] Tile_X0Y0_S1END[1] Tile_X0Y0_S1END[2] Tile_X0Y0_S1END[3] Tile_X0Y0_S2END[0]
+ Tile_X0Y0_S2END[1] Tile_X0Y0_S2END[2] Tile_X0Y0_S2END[3] Tile_X0Y0_S2END[4] Tile_X0Y0_S2END[5]
+ Tile_X0Y0_S2END[6] Tile_X0Y0_S2END[7] Tile_X0Y0_S2MID[0] Tile_X0Y0_S2MID[1] Tile_X0Y0_S2MID[2]
+ Tile_X0Y0_S2MID[3] Tile_X0Y0_S2MID[4] Tile_X0Y0_S2MID[5] Tile_X0Y0_S2MID[6] Tile_X0Y0_S2MID[7]
+ Tile_X0Y0_S4END[0] Tile_X0Y0_S4END[10] Tile_X0Y0_S4END[11] Tile_X0Y0_S4END[12] Tile_X0Y0_S4END[13]
+ Tile_X0Y0_S4END[14] Tile_X0Y0_S4END[15] Tile_X0Y0_S4END[1] Tile_X0Y0_S4END[2] Tile_X0Y0_S4END[3]
+ Tile_X0Y0_S4END[4] Tile_X0Y0_S4END[5] Tile_X0Y0_S4END[6] Tile_X0Y0_S4END[7] Tile_X0Y0_S4END[8]
+ Tile_X0Y0_S4END[9] Tile_X0Y0_UserCLKo Tile_X0Y0_W1BEG[0] Tile_X0Y0_W1BEG[1] Tile_X0Y0_W1BEG[2]
+ Tile_X0Y0_W1BEG[3] Tile_X0Y0_W2BEG[0] Tile_X0Y0_W2BEG[1] Tile_X0Y0_W2BEG[2] Tile_X0Y0_W2BEG[3]
+ Tile_X0Y0_W2BEG[4] Tile_X0Y0_W2BEG[5] Tile_X0Y0_W2BEG[6] Tile_X0Y0_W2BEG[7] Tile_X0Y0_W2BEGb[0]
+ Tile_X0Y0_W2BEGb[1] Tile_X0Y0_W2BEGb[2] Tile_X0Y0_W2BEGb[3] Tile_X0Y0_W2BEGb[4]
+ Tile_X0Y0_W2BEGb[5] Tile_X0Y0_W2BEGb[6] Tile_X0Y0_W2BEGb[7] Tile_X0Y0_W6BEG[0] Tile_X0Y0_W6BEG[10]
+ Tile_X0Y0_W6BEG[11] Tile_X0Y0_W6BEG[1] Tile_X0Y0_W6BEG[2] Tile_X0Y0_W6BEG[3] Tile_X0Y0_W6BEG[4]
+ Tile_X0Y0_W6BEG[5] Tile_X0Y0_W6BEG[6] Tile_X0Y0_W6BEG[7] Tile_X0Y0_W6BEG[8] Tile_X0Y0_W6BEG[9]
+ Tile_X0Y0_WW4BEG[0] Tile_X0Y0_WW4BEG[10] Tile_X0Y0_WW4BEG[11] Tile_X0Y0_WW4BEG[12]
+ Tile_X0Y0_WW4BEG[13] Tile_X0Y0_WW4BEG[14] Tile_X0Y0_WW4BEG[15] Tile_X0Y0_WW4BEG[1]
+ Tile_X0Y0_WW4BEG[2] Tile_X0Y0_WW4BEG[3] Tile_X0Y0_WW4BEG[4] Tile_X0Y0_WW4BEG[5]
+ Tile_X0Y0_WW4BEG[6] Tile_X0Y0_WW4BEG[7] Tile_X0Y0_WW4BEG[8] Tile_X0Y0_WW4BEG[9]
+ Tile_X0Y1_E1END[0] Tile_X0Y1_E1END[1] Tile_X0Y1_E1END[2] Tile_X0Y1_E1END[3] Tile_X0Y1_E2END[0]
+ Tile_X0Y1_E2END[1] Tile_X0Y1_E2END[2] Tile_X0Y1_E2END[3] Tile_X0Y1_E2END[4] Tile_X0Y1_E2END[5]
+ Tile_X0Y1_E2END[6] Tile_X0Y1_E2END[7] Tile_X0Y1_E2MID[0] Tile_X0Y1_E2MID[1] Tile_X0Y1_E2MID[2]
+ Tile_X0Y1_E2MID[3] Tile_X0Y1_E2MID[4] Tile_X0Y1_E2MID[5] Tile_X0Y1_E2MID[6] Tile_X0Y1_E2MID[7]
+ Tile_X0Y1_E6END[0] Tile_X0Y1_E6END[10] Tile_X0Y1_E6END[11] Tile_X0Y1_E6END[1] Tile_X0Y1_E6END[2]
+ Tile_X0Y1_E6END[3] Tile_X0Y1_E6END[4] Tile_X0Y1_E6END[5] Tile_X0Y1_E6END[6] Tile_X0Y1_E6END[7]
+ Tile_X0Y1_E6END[8] Tile_X0Y1_E6END[9] Tile_X0Y1_EE4END[0] Tile_X0Y1_EE4END[10] Tile_X0Y1_EE4END[11]
+ Tile_X0Y1_EE4END[12] Tile_X0Y1_EE4END[13] Tile_X0Y1_EE4END[14] Tile_X0Y1_EE4END[15]
+ Tile_X0Y1_EE4END[1] Tile_X0Y1_EE4END[2] Tile_X0Y1_EE4END[3] Tile_X0Y1_EE4END[4]
+ Tile_X0Y1_EE4END[5] Tile_X0Y1_EE4END[6] Tile_X0Y1_EE4END[7] Tile_X0Y1_EE4END[8]
+ Tile_X0Y1_EE4END[9] Tile_X0Y1_FrameData[0] Tile_X0Y1_FrameData[10] Tile_X0Y1_FrameData[11]
+ Tile_X0Y1_FrameData[12] Tile_X0Y1_FrameData[13] Tile_X0Y1_FrameData[14] Tile_X0Y1_FrameData[15]
+ Tile_X0Y1_FrameData[16] Tile_X0Y1_FrameData[17] Tile_X0Y1_FrameData[18] Tile_X0Y1_FrameData[19]
+ Tile_X0Y1_FrameData[1] Tile_X0Y1_FrameData[20] Tile_X0Y1_FrameData[21] Tile_X0Y1_FrameData[22]
+ Tile_X0Y1_FrameData[23] Tile_X0Y1_FrameData[24] Tile_X0Y1_FrameData[25] Tile_X0Y1_FrameData[26]
+ Tile_X0Y1_FrameData[27] Tile_X0Y1_FrameData[28] Tile_X0Y1_FrameData[29] Tile_X0Y1_FrameData[2]
+ Tile_X0Y1_FrameData[30] Tile_X0Y1_FrameData[31] Tile_X0Y1_FrameData[3] Tile_X0Y1_FrameData[4]
+ Tile_X0Y1_FrameData[5] Tile_X0Y1_FrameData[6] Tile_X0Y1_FrameData[7] Tile_X0Y1_FrameData[8]
+ Tile_X0Y1_FrameData[9] Tile_X0Y1_FrameData_O[0] Tile_X0Y1_FrameData_O[10] Tile_X0Y1_FrameData_O[11]
+ Tile_X0Y1_FrameData_O[12] Tile_X0Y1_FrameData_O[13] Tile_X0Y1_FrameData_O[14] Tile_X0Y1_FrameData_O[15]
+ Tile_X0Y1_FrameData_O[16] Tile_X0Y1_FrameData_O[17] Tile_X0Y1_FrameData_O[18] Tile_X0Y1_FrameData_O[19]
+ Tile_X0Y1_FrameData_O[1] Tile_X0Y1_FrameData_O[20] Tile_X0Y1_FrameData_O[21] Tile_X0Y1_FrameData_O[22]
+ Tile_X0Y1_FrameData_O[23] Tile_X0Y1_FrameData_O[24] Tile_X0Y1_FrameData_O[25] Tile_X0Y1_FrameData_O[26]
+ Tile_X0Y1_FrameData_O[27] Tile_X0Y1_FrameData_O[28] Tile_X0Y1_FrameData_O[29] Tile_X0Y1_FrameData_O[2]
+ Tile_X0Y1_FrameData_O[30] Tile_X0Y1_FrameData_O[31] Tile_X0Y1_FrameData_O[3] Tile_X0Y1_FrameData_O[4]
+ Tile_X0Y1_FrameData_O[5] Tile_X0Y1_FrameData_O[6] Tile_X0Y1_FrameData_O[7] Tile_X0Y1_FrameData_O[8]
+ Tile_X0Y1_FrameData_O[9] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_FrameStrobe[10] Tile_X0Y1_FrameStrobe[11]
+ Tile_X0Y1_FrameStrobe[12] Tile_X0Y1_FrameStrobe[13] Tile_X0Y1_FrameStrobe[14] Tile_X0Y1_FrameStrobe[15]
+ Tile_X0Y1_FrameStrobe[16] Tile_X0Y1_FrameStrobe[17] Tile_X0Y1_FrameStrobe[18] Tile_X0Y1_FrameStrobe[19]
+ Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_FrameStrobe[4]
+ Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_FrameStrobe[8]
+ Tile_X0Y1_FrameStrobe[9] Tile_X0Y1_N1END[0] Tile_X0Y1_N1END[1] Tile_X0Y1_N1END[2]
+ Tile_X0Y1_N1END[3] Tile_X0Y1_N2END[0] Tile_X0Y1_N2END[1] Tile_X0Y1_N2END[2] Tile_X0Y1_N2END[3]
+ Tile_X0Y1_N2END[4] Tile_X0Y1_N2END[5] Tile_X0Y1_N2END[6] Tile_X0Y1_N2END[7] Tile_X0Y1_N2MID[0]
+ Tile_X0Y1_N2MID[1] Tile_X0Y1_N2MID[2] Tile_X0Y1_N2MID[3] Tile_X0Y1_N2MID[4] Tile_X0Y1_N2MID[5]
+ Tile_X0Y1_N2MID[6] Tile_X0Y1_N2MID[7] Tile_X0Y1_N4END[0] Tile_X0Y1_N4END[10] Tile_X0Y1_N4END[11]
+ Tile_X0Y1_N4END[12] Tile_X0Y1_N4END[13] Tile_X0Y1_N4END[14] Tile_X0Y1_N4END[15]
+ Tile_X0Y1_N4END[1] Tile_X0Y1_N4END[2] Tile_X0Y1_N4END[3] Tile_X0Y1_N4END[4] Tile_X0Y1_N4END[5]
+ Tile_X0Y1_N4END[6] Tile_X0Y1_N4END[7] Tile_X0Y1_N4END[8] Tile_X0Y1_N4END[9] Tile_X0Y1_S1BEG[0]
+ Tile_X0Y1_S1BEG[1] Tile_X0Y1_S1BEG[2] Tile_X0Y1_S1BEG[3] Tile_X0Y1_S2BEG[0] Tile_X0Y1_S2BEG[1]
+ Tile_X0Y1_S2BEG[2] Tile_X0Y1_S2BEG[3] Tile_X0Y1_S2BEG[4] Tile_X0Y1_S2BEG[5] Tile_X0Y1_S2BEG[6]
+ Tile_X0Y1_S2BEG[7] Tile_X0Y1_S2BEGb[0] Tile_X0Y1_S2BEGb[1] Tile_X0Y1_S2BEGb[2] Tile_X0Y1_S2BEGb[3]
+ Tile_X0Y1_S2BEGb[4] Tile_X0Y1_S2BEGb[5] Tile_X0Y1_S2BEGb[6] Tile_X0Y1_S2BEGb[7]
+ Tile_X0Y1_S4BEG[0] Tile_X0Y1_S4BEG[10] Tile_X0Y1_S4BEG[11] Tile_X0Y1_S4BEG[12] Tile_X0Y1_S4BEG[13]
+ Tile_X0Y1_S4BEG[14] Tile_X0Y1_S4BEG[15] Tile_X0Y1_S4BEG[1] Tile_X0Y1_S4BEG[2] Tile_X0Y1_S4BEG[3]
+ Tile_X0Y1_S4BEG[4] Tile_X0Y1_S4BEG[5] Tile_X0Y1_S4BEG[6] Tile_X0Y1_S4BEG[7] Tile_X0Y1_S4BEG[8]
+ Tile_X0Y1_S4BEG[9] Tile_X0Y1_UserCLK Tile_X0Y1_W1BEG[0] Tile_X0Y1_W1BEG[1] Tile_X0Y1_W1BEG[2]
+ Tile_X0Y1_W1BEG[3] Tile_X0Y1_W2BEG[0] Tile_X0Y1_W2BEG[1] Tile_X0Y1_W2BEG[2] Tile_X0Y1_W2BEG[3]
+ Tile_X0Y1_W2BEG[4] Tile_X0Y1_W2BEG[5] Tile_X0Y1_W2BEG[6] Tile_X0Y1_W2BEG[7] Tile_X0Y1_W2BEGb[0]
+ Tile_X0Y1_W2BEGb[1] Tile_X0Y1_W2BEGb[2] Tile_X0Y1_W2BEGb[3] Tile_X0Y1_W2BEGb[4]
+ Tile_X0Y1_W2BEGb[5] Tile_X0Y1_W2BEGb[6] Tile_X0Y1_W2BEGb[7] Tile_X0Y1_W6BEG[0] Tile_X0Y1_W6BEG[10]
+ Tile_X0Y1_W6BEG[11] Tile_X0Y1_W6BEG[1] Tile_X0Y1_W6BEG[2] Tile_X0Y1_W6BEG[3] Tile_X0Y1_W6BEG[4]
+ Tile_X0Y1_W6BEG[5] Tile_X0Y1_W6BEG[6] Tile_X0Y1_W6BEG[7] Tile_X0Y1_W6BEG[8] Tile_X0Y1_W6BEG[9]
+ Tile_X0Y1_WW4BEG[0] Tile_X0Y1_WW4BEG[10] Tile_X0Y1_WW4BEG[11] Tile_X0Y1_WW4BEG[12]
+ Tile_X0Y1_WW4BEG[13] Tile_X0Y1_WW4BEG[14] Tile_X0Y1_WW4BEG[15] Tile_X0Y1_WW4BEG[1]
+ Tile_X0Y1_WW4BEG[2] Tile_X0Y1_WW4BEG[3] Tile_X0Y1_WW4BEG[4] Tile_X0Y1_WW4BEG[5]
+ Tile_X0Y1_WW4BEG[6] Tile_X0Y1_WW4BEG[7] Tile_X0Y1_WW4BEG[8] Tile_X0Y1_WW4BEG[9]
+ VGND VPWR WEN_SRAM
X_0367_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit24.Q net35
+ net61 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG13 _0059_
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit25.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1BEG1
+ VPWR VGND sg13g2_mux4_1
X_0298_ VPWR _0001_ net151 VGND sg13g2_inv_1
XFILLER_89_100 VPWR VGND sg13g2_decap_8
XFILLER_117_88 VPWR VGND sg13g2_decap_8
XFILLER_26_63 VPWR VGND sg13g2_fill_1
XFILLER_3_34 VPWR VGND sg13g2_decap_8
XFILLER_67_70 VPWR VGND sg13g2_fill_1
X_1270_ net199 net706 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
Xoutput412 net412 Tile_X0Y0_N4BEG[6] VPWR VGND sg13g2_buf_1
Xoutput401 net401 Tile_X0Y0_N4BEG[10] VPWR VGND sg13g2_buf_1
X_0985_ net786 net710 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
X_1606_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG11 net451 VPWR
+ VGND sg13g2_buf_1
Xoutput434 net434 Tile_X0Y0_W2BEGb[5] VPWR VGND sg13g2_buf_1
Xoutput423 net423 Tile_X0Y0_W2BEG[2] VPWR VGND sg13g2_buf_1
Xoutput489 net489 Tile_X0Y1_FrameData_O[31] VPWR VGND sg13g2_buf_1
Xoutput478 net478 Tile_X0Y1_FrameData_O[21] VPWR VGND sg13g2_buf_1
Xoutput467 net467 Tile_X0Y1_FrameData_O[11] VPWR VGND sg13g2_buf_1
X_0419_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit16.Q net37
+ net46 net38 net623 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit17.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG7 VPWR VGND sg13g2_mux4_1
X_1537_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG7 net391 VPWR
+ VGND sg13g2_buf_1
Xoutput445 net445 Tile_X0Y0_W6BEG[6] VPWR VGND sg13g2_buf_1
Xoutput456 net456 Tile_X0Y0_WW4BEG[1] VPWR VGND sg13g2_buf_1
X_1468_ net778 net643 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
X_1399_ net773 net662 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_88_25 VPWR VGND sg13g2_fill_1
Xfanout672 net673 net672 VPWR VGND sg13g2_buf_1
Xfanout683 net684 net683 VPWR VGND sg13g2_buf_1
Xfanout661 net668 net661 VPWR VGND sg13g2_buf_1
Xfanout694 net695 net694 VPWR VGND sg13g2_buf_1
Xfanout650 net651 net650 VPWR VGND sg13g2_buf_1
X_0770_ VGND VPWR _0026_ _0210_ _0211_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit13.Q
+ sg13g2_a21oi_1
XFILLER_78_91 VPWR VGND sg13g2_fill_1
X_1253_ net215 net717 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
X_1322_ net758 net682 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_91_172 VPWR VGND sg13g2_fill_2
XFILLER_91_150 VPWR VGND sg13g2_fill_1
X_1184_ net220 net742 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
X_0968_ net799 net709 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
X_0899_ net794 net733 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
Xoutput253 net253 ADDR_SRAM2 VPWR VGND sg13g2_buf_1
Xoutput275 net275 BM_SRAM21 VPWR VGND sg13g2_buf_1
Xoutput264 net264 BM_SRAM11 VPWR VGND sg13g2_buf_1
Xoutput286 net286 BM_SRAM31 VPWR VGND sg13g2_buf_1
Xoutput297 net297 DIN_SRAM11 VPWR VGND sg13g2_buf_1
XFILLER_2_154 VPWR VGND sg13g2_decap_8
XFILLER_64_60 VPWR VGND sg13g2_decap_4
XFILLER_48_72 VPWR VGND sg13g2_fill_1
XFILLER_119_108 VPWR VGND sg13g2_decap_8
X_0822_ _0258_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit2.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit1.Q VPWR VGND
+ sg13g2_nand2b_1
X_0753_ VGND VPWR _0022_ _0194_ _0196_ _0195_ sg13g2_a21oi_1
X_0684_ _0162_ VPWR net251 VGND Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit19.Q
+ _0164_ sg13g2_o21ai_1
X_1305_ net775 net693 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_29_0 VPWR VGND sg13g2_fill_1
X_1236_ net202 net715 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
X_1098_ net801 net663 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
X_1167_ net207 net742 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_118_174 VPWR VGND sg13g2_decap_8
XFILLER_109_12 VPWR VGND sg13g2_fill_2
XFILLER_109_78 VPWR VGND sg13g2_fill_2
XFILLER_70_164 VPWR VGND sg13g2_fill_1
XFILLER_34_85 VPWR VGND sg13g2_fill_2
X_1021_ net802 net699 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
X_0805_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit13.Q VPWR
+ _0243_ VGND Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit12.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG14 sg13g2_o21ai_1
X_0598_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit28.Q VPWR
+ _0153_ VGND Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit27.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG15 sg13g2_o21ai_1
X_0667_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit8.Q net223
+ net243 _0088_ net138 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit9.Q
+ _0161_ VPWR VGND sg13g2_mux4_1
X_0736_ net142 net174 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit2.Q
+ _0180_ VPWR VGND sg13g2_mux2_1
X_1219_ net217 net728 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_52_120 VPWR VGND sg13g2_decap_8
XFILLER_121_136 VPWR VGND sg13g2_decap_8
XFILLER_106_199 VPWR VGND sg13g2_fill_2
XFILLER_106_177 VPWR VGND sg13g2_fill_1
XFILLER_29_96 VPWR VGND sg13g2_fill_1
XFILLER_77_8 VPWR VGND sg13g2_fill_1
XFILLER_61_94 VPWR VGND sg13g2_fill_1
X_0452_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit6.Q net10
+ net23 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG15 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG7
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit7.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG0
+ VPWR VGND sg13g2_mux4_1
X_1570_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG3 net424 VPWR
+ VGND sg13g2_buf_1
X_0521_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit22.Q net34
+ net76 net69 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG12 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit23.Q
+ net282 VPWR VGND sg13g2_mux4_1
XFILLER_6_45 VPWR VGND sg13g2_decap_8
X_0383_ _0076_ _0074_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit30.Q
+ VPWR VGND sg13g2_nand2b_1
X_1004_ net804 net698 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_103_158 VPWR VGND sg13g2_fill_2
X_1699_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG0 net553 VPWR
+ VGND sg13g2_buf_1
X_0719_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit0.Q net182
+ net175 net166 _0159_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit1.Q
+ net306 VPWR VGND sg13g2_mux4_1
XFILLER_15_65 VPWR VGND sg13g2_fill_2
XFILLER_31_64 VPWR VGND sg13g2_fill_2
Xinput120 Tile_X0Y0_S2END[2] net120 VPWR VGND sg13g2_buf_1
Xinput131 Tile_X0Y0_S2MID[5] net131 VPWR VGND sg13g2_buf_1
Xinput153 Tile_X0Y1_E2END[7] net153 VPWR VGND sg13g2_buf_1
Xinput142 Tile_X0Y1_E1END[0] net142 VPWR VGND sg13g2_buf_1
Xinput186 Tile_X0Y1_EE4END[6] net186 VPWR VGND sg13g2_buf_1
Xinput175 Tile_X0Y1_EE4END[10] net175 VPWR VGND sg13g2_buf_1
Xinput164 Tile_X0Y1_E6END[11] net164 VPWR VGND sg13g2_buf_1
Xinput197 Tile_X0Y1_FrameData[16] net197 VPWR VGND sg13g2_buf_1
XFILLER_31_123 VPWR VGND sg13g2_decap_4
XFILLER_68_4 VPWR VGND sg13g2_fill_2
X_1622_ net779 net467 VPWR VGND sg13g2_buf_1
X_1553_ Tile_X0Y1_N4END[15] net413 VPWR VGND sg13g2_buf_1
X_1484_ net812 net329 VPWR VGND sg13g2_buf_1
X_0504_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit20.Q net75
+ net68 net56 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG11 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit21.Q
+ net314 VPWR VGND sg13g2_mux4_1
X_0435_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit5.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END3
+ net11 net117 net15 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit4.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W1BEG3 VPWR VGND sg13g2_mux4_1
X_0366_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit2.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END1
+ net248 net115 net135 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit3.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG13 VPWR VGND sg13g2_mux4_1
X_0297_ VPWR _0000_ net157 VGND sg13g2_inv_1
XFILLER_117_67 VPWR VGND sg13g2_decap_8
Xfanout810 net85 net810 VPWR VGND sg13g2_buf_1
X_0984_ net785 net709 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
Xoutput402 net402 Tile_X0Y0_N4BEG[11] VPWR VGND sg13g2_buf_1
Xoutput413 net413 Tile_X0Y0_N4BEG[7] VPWR VGND sg13g2_buf_1
Xoutput468 net468 Tile_X0Y1_FrameData_O[12] VPWR VGND sg13g2_buf_1
X_1536_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG6 net390 VPWR
+ VGND sg13g2_buf_1
Xoutput446 net446 Tile_X0Y0_W6BEG[7] VPWR VGND sg13g2_buf_1
X_1605_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG10 net450 VPWR
+ VGND sg13g2_buf_1
Xoutput457 net457 Tile_X0Y0_WW4BEG[2] VPWR VGND sg13g2_buf_1
Xoutput435 net435 Tile_X0Y0_W2BEGb[6] VPWR VGND sg13g2_buf_1
Xoutput424 net424 Tile_X0Y0_W2BEG[3] VPWR VGND sg13g2_buf_1
XFILLER_59_0 VPWR VGND sg13g2_fill_1
Xoutput479 net479 Tile_X0Y1_FrameData_O[22] VPWR VGND sg13g2_buf_1
X_0418_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit10.Q net47
+ net39 net57 net624 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit11.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG6 VPWR VGND sg13g2_mux4_1
X_0349_ _0048_ VPWR _0049_ VGND Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit30.Q
+ net149 sg13g2_o21ai_1
X_1398_ net772 net659 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
X_1467_ net777 net643 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_12_88 VPWR VGND sg13g2_fill_1
XFILLER_10_115 VPWR VGND sg13g2_fill_1
Xfanout640 _0043_ net640 VPWR VGND sg13g2_buf_1
Xfanout651 net222 net651 VPWR VGND sg13g2_buf_1
XFILLER_85_170 VPWR VGND sg13g2_fill_2
Xfanout673 net674 net673 VPWR VGND sg13g2_buf_1
Xfanout684 net691 net684 VPWR VGND sg13g2_buf_1
Xfanout695 net696 net695 VPWR VGND sg13g2_buf_1
XFILLER_37_85 VPWR VGND sg13g2_fill_2
Xfanout662 net668 net662 VPWR VGND sg13g2_buf_1
XFILLER_53_62 VPWR VGND sg13g2_decap_4
XFILLER_83_107 VPWR VGND sg13g2_decap_8
X_1321_ net757 net682 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
X_1252_ net216 net715 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
X_1183_ net221 net742 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
X_0967_ net798 net709 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
X_1519_ Tile_X0Y1_FrameStrobe[13] net364 VPWR VGND sg13g2_buf_1
X_0898_ net102 net735 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
Xoutput298 net298 DIN_SRAM12 VPWR VGND sg13g2_buf_1
Xoutput254 net254 ADDR_SRAM3 VPWR VGND sg13g2_buf_1
Xoutput287 net287 BM_SRAM4 VPWR VGND sg13g2_buf_1
Xoutput265 net265 BM_SRAM12 VPWR VGND sg13g2_buf_1
Xoutput276 net276 BM_SRAM22 VPWR VGND sg13g2_buf_1
XFILLER_23_43 VPWR VGND sg13g2_fill_2
XFILLER_23_98 VPWR VGND sg13g2_fill_2
XFILLER_65_118 VPWR VGND sg13g2_decap_8
XFILLER_2_133 VPWR VGND sg13g2_decap_8
XFILLER_0_69 VPWR VGND sg13g2_decap_4
X_0752_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit7.Q VPWR
+ _0195_ VGND _0192_ _0193_ sg13g2_o21ai_1
X_0821_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit2.Q Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit1.Q
+ _0257_ VPWR VGND sg13g2_nor2b_1
X_0683_ VGND VPWR net146 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit18.Q
+ _0164_ _0163_ sg13g2_a21oi_1
X_1166_ net763 net739 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
X_1304_ net774 net694 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
X_1235_ net203 net714 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_49_181 VPWR VGND sg13g2_fill_1
X_1097_ net800 net663 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_64_173 VPWR VGND sg13g2_decap_8
XFILLER_118_153 VPWR VGND sg13g2_decap_8
XFILLER_47_118 VPWR VGND sg13g2_fill_1
XFILLER_55_195 VPWR VGND sg13g2_fill_2
X_1020_ net791 net702 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_61_121 VPWR VGND sg13g2_fill_1
XFILLER_61_110 VPWR VGND sg13g2_decap_8
X_0735_ _0178_ VPWR _0179_ VGND _0019_ _0161_ sg13g2_o21ai_1
X_0804_ _0031_ net633 _0242_ VPWR VGND sg13g2_nor2_1
X_0597_ net623 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit27.Q
+ _0152_ VPWR VGND sg13g2_nor2b_1
X_0666_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit22.Q net14
+ net8 _0160_ net639 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit23.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG14 VPWR VGND sg13g2_mux4_1
X_1149_ net93 net654 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
X_1218_ net753 net728 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_121_115 VPWR VGND sg13g2_decap_8
XFILLER_106_101 VPWR VGND sg13g2_fill_2
XFILLER_28_151 VPWR VGND sg13g2_fill_1
XFILLER_61_51 VPWR VGND sg13g2_decap_8
X_0520_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit20.Q net75
+ net68 net56 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG11 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit21.Q
+ net281 VPWR VGND sg13g2_mux4_1
X_0451_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit4.Q net18
+ net27 net631 net623 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit5.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb7 VPWR VGND sg13g2_mux4_1
X_0382_ net226 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit30.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit31.Q _0075_ VPWR
+ VGND sg13g2_nor3_1
X_1003_ net803 net698 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_34_121 VPWR VGND sg13g2_fill_2
XFILLER_89_0 VPWR VGND sg13g2_fill_2
XFILLER_34_143 VPWR VGND sg13g2_fill_1
X_1698_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb7 net552 VPWR
+ VGND sg13g2_buf_1
X_0718_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit30.Q net181
+ net189 net165 _0160_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit31.Q
+ net295 VPWR VGND sg13g2_mux4_1
X_0649_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit26.Q net224
+ net244 _0060_ net139 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit27.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG9 VPWR VGND sg13g2_mux4_1
XFILLER_122_24 VPWR VGND sg13g2_fill_1
XFILLER_31_32 VPWR VGND sg13g2_fill_1
Xinput110 Tile_X0Y0_FrameData[6] net110 VPWR VGND sg13g2_buf_1
XFILLER_103_2 VPWR VGND sg13g2_fill_1
Xinput121 Tile_X0Y0_S2END[3] net121 VPWR VGND sg13g2_buf_1
Xinput132 Tile_X0Y0_S2MID[6] net132 VPWR VGND sg13g2_buf_1
Xinput143 Tile_X0Y1_E1END[1] net143 VPWR VGND sg13g2_buf_1
Xinput154 Tile_X0Y1_E2MID[0] net154 VPWR VGND sg13g2_buf_1
Xinput187 Tile_X0Y1_EE4END[7] net187 VPWR VGND sg13g2_buf_1
Xinput165 Tile_X0Y1_E6END[1] net165 VPWR VGND sg13g2_buf_1
Xinput176 Tile_X0Y1_EE4END[11] net176 VPWR VGND sg13g2_buf_1
Xinput198 Tile_X0Y1_FrameData[17] net198 VPWR VGND sg13g2_buf_1
X_1552_ Tile_X0Y1_N4END[14] net412 VPWR VGND sg13g2_buf_1
X_1621_ net780 net466 VPWR VGND sg13g2_buf_1
X_0503_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit18.Q net74
+ net67 net55 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG10 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit19.Q
+ net313 VPWR VGND sg13g2_mux4_1
X_1483_ net113 net359 VPWR VGND sg13g2_buf_1
X_0434_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit3.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END2
+ net10 net116 net16 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit2.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W1BEG2 VPWR VGND sg13g2_mux4_1
X_0365_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit13.Q net143
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG13 net169 _0063_
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit12.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END1
+ VPWR VGND sg13g2_mux4_1
XFILLER_117_46 VPWR VGND sg13g2_decap_8
Xfanout800 net95 net800 VPWR VGND sg13g2_buf_1
Xfanout811 net84 net811 VPWR VGND sg13g2_buf_1
XFILLER_89_124 VPWR VGND sg13g2_fill_2
XFILLER_93_49 VPWR VGND sg13g2_fill_2
XFILLER_13_102 VPWR VGND sg13g2_decap_8
XFILLER_3_69 VPWR VGND sg13g2_decap_8
X_0983_ net784 net709 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_8_150 VPWR VGND sg13g2_fill_2
Xoutput414 net414 Tile_X0Y0_N4BEG[8] VPWR VGND sg13g2_buf_1
Xoutput403 net403 Tile_X0Y0_N4BEG[12] VPWR VGND sg13g2_buf_1
Xoutput469 net469 Tile_X0Y1_FrameData_O[13] VPWR VGND sg13g2_buf_1
X_1535_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG5 net389 VPWR
+ VGND sg13g2_buf_1
Xoutput447 net447 Tile_X0Y0_W6BEG[8] VPWR VGND sg13g2_buf_1
X_1604_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG9 net464 VPWR
+ VGND sg13g2_buf_1
Xoutput458 net458 Tile_X0Y0_WW4BEG[3] VPWR VGND sg13g2_buf_1
Xoutput436 net436 Tile_X0Y0_W2BEGb[7] VPWR VGND sg13g2_buf_1
Xoutput425 net425 Tile_X0Y0_W2BEG[4] VPWR VGND sg13g2_buf_1
X_0417_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit21.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb6
+ net132 net241 net124 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit20.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG6 VPWR VGND sg13g2_mux4_1
X_0348_ _0048_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit30.Q
+ _0002_ VPWR VGND sg13g2_nand2_1
X_1397_ net771 net659 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
X_1466_ net776 net642 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
Xfanout652 net656 net652 VPWR VGND sg13g2_buf_1
Xfanout685 net689 net685 VPWR VGND sg13g2_buf_1
Xfanout663 net667 net663 VPWR VGND sg13g2_buf_1
Xfanout630 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG1 net630
+ VPWR VGND sg13g2_buf_1
Xfanout674 Tile_X0Y1_FrameStrobe[6] net674 VPWR VGND sg13g2_buf_1
Xfanout641 net643 net641 VPWR VGND sg13g2_buf_1
Xfanout696 Tile_X0Y1_FrameStrobe[4] net696 VPWR VGND sg13g2_buf_1
X_1320_ net190 net696 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
X_1182_ net780 net738 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
X_1251_ net754 net714 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_91_174 VPWR VGND sg13g2_fill_1
X_0897_ net103 net735 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
X_0966_ net797 net709 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_71_0 VPWR VGND sg13g2_fill_2
X_1518_ Tile_X0Y1_FrameStrobe[12] net363 VPWR VGND sg13g2_buf_1
Xoutput299 net299 DIN_SRAM13 VPWR VGND sg13g2_buf_1
Xoutput255 net255 ADDR_SRAM4 VPWR VGND sg13g2_buf_1
Xoutput288 net288 BM_SRAM5 VPWR VGND sg13g2_buf_1
X_1449_ net757 net641 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
Xoutput266 net266 BM_SRAM13 VPWR VGND sg13g2_buf_1
Xoutput277 net277 BM_SRAM23 VPWR VGND sg13g2_buf_1
XFILLER_99_48 VPWR VGND sg13g2_fill_2
XFILLER_2_112 VPWR VGND sg13g2_decap_8
XFILLER_2_189 VPWR VGND sg13g2_decap_8
XFILLER_48_85 VPWR VGND sg13g2_fill_1
XFILLER_120_90 VPWR VGND sg13g2_decap_8
X_0751_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG5 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG9
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit5.Q _0194_ VPWR
+ VGND sg13g2_mux2_1
X_0820_ VGND VPWR _0249_ _0251_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S4BEG3
+ _0256_ sg13g2_a21oi_1
X_0682_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit18.Q net154
+ _0163_ VPWR VGND sg13g2_nor2b_1
X_1303_ net773 net694 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
X_1096_ net799 net663 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
X_1234_ net767 net716 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
X_1165_ net762 net739 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_118_132 VPWR VGND sg13g2_decap_8
XFILLER_109_14 VPWR VGND sg13g2_fill_1
X_0949_ net782 net719 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_87_200 VPWR VGND sg13g2_fill_1
XFILLER_70_111 VPWR VGND sg13g2_fill_1
XFILLER_18_66 VPWR VGND sg13g2_fill_1
XFILLER_50_64 VPWR VGND sg13g2_fill_2
XFILLER_78_200 VPWR VGND sg13g2_fill_1
XFILLER_61_188 VPWR VGND sg13g2_decap_4
X_0665_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit10.Q net224
+ net244 _0060_ net139 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit11.Q
+ _0160_ VPWR VGND sg13g2_mux4_1
X_0734_ VPWR _0178_ _0177_ VGND sg13g2_inv_1
X_0803_ VGND VPWR _0032_ _0240_ _0241_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit14.Q
+ sg13g2_a21oi_1
X_0596_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG7 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG11
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit27.Q _0151_ VPWR
+ VGND sg13g2_mux2_1
XFILLER_69_200 VPWR VGND sg13g2_fill_1
XFILLER_111_59 VPWR VGND sg13g2_fill_2
X_1148_ net791 net654 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
X_1079_ net784 net676 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_37_163 VPWR VGND sg13g2_fill_2
X_1217_ net752 net729 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_106_124 VPWR VGND sg13g2_fill_2
XFILLER_20_78 VPWR VGND sg13g2_fill_2
XFILLER_45_31 VPWR VGND sg13g2_fill_2
XFILLER_43_188 VPWR VGND sg13g2_fill_1
XFILLER_61_74 VPWR VGND sg13g2_decap_8
XFILLER_6_25 VPWR VGND sg13g2_fill_2
XFILLER_120_160 VPWR VGND sg13g2_decap_8
X_0381_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit0.Q net37
+ net56 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG15 _0073_
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit1.Q _0074_ VPWR
+ VGND sg13g2_mux4_1
X_0450_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit2.Q net17
+ net26 net630 net624 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit3.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb6 VPWR VGND sg13g2_mux4_1
XIHP_SRAM_582 VPWR VGND TIE_LOW_SRAM sg13g2_tielo
X_1002_ net801 net697 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_19_163 VPWR VGND sg13g2_fill_2
X_1697_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb6 net551 VPWR
+ VGND sg13g2_buf_1
X_0648_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit4.Q net29
+ net33 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG10 net638
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit5.Q Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG5
+ VPWR VGND sg13g2_mux4_1
X_0717_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit28.Q net174
+ net188 net162 _0161_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit29.Q
+ net294 VPWR VGND sg13g2_mux4_1
X_0579_ _0134_ _0136_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S4BEG0
+ VPWR VGND sg13g2_nor2_1
XFILLER_15_67 VPWR VGND sg13g2_fill_1
XFILLER_40_125 VPWR VGND sg13g2_decap_4
XFILLER_31_66 VPWR VGND sg13g2_fill_1
Xinput122 Tile_X0Y0_S2END[4] net122 VPWR VGND sg13g2_buf_1
Xinput133 Tile_X0Y0_S2MID[7] net133 VPWR VGND sg13g2_buf_1
Xinput100 Tile_X0Y0_FrameData[26] net100 VPWR VGND sg13g2_buf_1
Xinput111 Tile_X0Y0_FrameData[7] net111 VPWR VGND sg13g2_buf_1
Xinput144 Tile_X0Y1_E1END[2] net144 VPWR VGND sg13g2_buf_1
XFILLER_16_122 VPWR VGND sg13g2_fill_1
Xinput155 Tile_X0Y1_E2MID[1] net155 VPWR VGND sg13g2_buf_1
Xinput188 Tile_X0Y1_EE4END[8] net188 VPWR VGND sg13g2_buf_1
Xinput177 Tile_X0Y1_EE4END[12] net177 VPWR VGND sg13g2_buf_1
Xinput166 Tile_X0Y1_E6END[2] net166 VPWR VGND sg13g2_buf_1
Xinput199 Tile_X0Y1_FrameData[18] net199 VPWR VGND sg13g2_buf_1
XFILLER_112_91 VPWR VGND sg13g2_fill_1
XFILLER_72_73 VPWR VGND sg13g2_fill_2
X_1551_ Tile_X0Y1_N4END[13] net411 VPWR VGND sg13g2_buf_1
X_0502_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit16.Q net73
+ net81 net65 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG9 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit17.Q
+ net312 VPWR VGND sg13g2_mux4_1
X_1482_ net783 net358 VPWR VGND sg13g2_buf_1
XFILLER_68_6 VPWR VGND sg13g2_fill_1
X_1620_ net750 net496 VPWR VGND sg13g2_buf_1
X_0433_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit1.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END1
+ net13 net115 net17 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit0.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W1BEG1 VPWR VGND sg13g2_mux4_1
X_0364_ VGND VPWR _0061_ _0062_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit27.Q
+ _0009_ _0063_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit26.Q
+ sg13g2_a221oi_1
Xfanout801 net94 net801 VPWR VGND sg13g2_buf_1
Xfanout812 net83 net812 VPWR VGND sg13g2_buf_1
XFILLER_122_200 VPWR VGND sg13g2_fill_1
XFILLER_3_48 VPWR VGND sg13g2_decap_8
X_0982_ net783 net708 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_12_191 VPWR VGND sg13g2_fill_2
Xoutput404 net404 Tile_X0Y0_N4BEG[13] VPWR VGND sg13g2_buf_1
Xoutput415 net415 Tile_X0Y0_N4BEG[9] VPWR VGND sg13g2_buf_1
X_1603_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG8 net463 VPWR
+ VGND sg13g2_buf_1
Xoutput448 net448 Tile_X0Y0_W6BEG[9] VPWR VGND sg13g2_buf_1
Xoutput437 net437 Tile_X0Y0_W6BEG[0] VPWR VGND sg13g2_buf_1
XFILLER_86_128 VPWR VGND sg13g2_fill_1
Xoutput459 net459 Tile_X0Y0_WW4BEG[4] VPWR VGND sg13g2_buf_1
Xoutput426 net426 Tile_X0Y0_W2BEG[5] VPWR VGND sg13g2_buf_1
X_1534_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG4 net388 VPWR
+ VGND sg13g2_buf_1
X_1465_ net775 net643 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
X_0347_ _0044_ _0046_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit28.Q
+ _0047_ VPWR VGND sg13g2_nand3_1
X_1396_ net769 net658 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
X_0416_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit31.Q net155
+ net165 net147 _0083_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit30.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb6 VPWR VGND sg13g2_mux4_1
XFILLER_104_200 VPWR VGND sg13g2_fill_1
Xfanout664 net665 net664 VPWR VGND sg13g2_buf_1
Xfanout653 net656 net653 VPWR VGND sg13g2_buf_1
Xfanout675 net677 net675 VPWR VGND sg13g2_buf_1
Xfanout631 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG0 net631
+ VPWR VGND sg13g2_buf_1
Xfanout697 net699 net697 VPWR VGND sg13g2_buf_1
Xfanout686 net689 net686 VPWR VGND sg13g2_buf_1
XFILLER_77_139 VPWR VGND sg13g2_fill_1
Xfanout642 net643 net642 VPWR VGND sg13g2_buf_1
XFILLER_118_90 VPWR VGND sg13g2_decap_8
XFILLER_5_176 VPWR VGND sg13g2_decap_8
XFILLER_45_8 VPWR VGND sg13g2_fill_2
XFILLER_94_82 VPWR VGND sg13g2_fill_2
X_1181_ net779 net738 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
X_1250_ net753 net716 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
X_0896_ net105 net734 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
X_0965_ net796 net709 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_64_0 VPWR VGND sg13g2_decap_8
X_1517_ Tile_X0Y1_FrameStrobe[11] net362 VPWR VGND sg13g2_buf_1
XFILLER_114_15 VPWR VGND sg13g2_fill_1
XFILLER_4_80 VPWR VGND sg13g2_fill_2
Xoutput256 net256 ADDR_SRAM5 VPWR VGND sg13g2_buf_1
Xoutput289 net289 BM_SRAM6 VPWR VGND sg13g2_buf_1
Xoutput267 net267 BM_SRAM14 VPWR VGND sg13g2_buf_1
X_1448_ net781 net647 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
Xoutput278 net278 BM_SRAM24 VPWR VGND sg13g2_buf_1
XFILLER_82_153 VPWR VGND sg13g2_fill_1
XFILLER_67_194 VPWR VGND sg13g2_fill_2
X_1379_ net754 net669 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_2_168 VPWR VGND sg13g2_decap_8
XFILLER_48_97 VPWR VGND sg13g2_fill_1
XFILLER_9_25 VPWR VGND sg13g2_fill_2
X_0750_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit6.Q VPWR
+ _0193_ VGND Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit5.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG13 sg13g2_o21ai_1
X_0681_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit19.Q net640
+ _0162_ VPWR VGND Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit18.Q
+ sg13g2_nand3b_1
X_1302_ net772 net692 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
X_1233_ net766 net716 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
X_1095_ net798 net663 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
X_1164_ net210 net741 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_118_111 VPWR VGND sg13g2_decap_8
X_0948_ net83 net722 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_118_188 VPWR VGND sg13g2_decap_4
X_0879_ net88 net744 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_91_61 VPWR VGND sg13g2_fill_1
X_0802_ net144 net179 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit12.Q
+ _0240_ VPWR VGND sg13g2_mux2_1
X_0664_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit20.Q net3
+ net7 _0159_ net638 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit21.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG13 VPWR VGND sg13g2_mux4_1
X_0733_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit3.Q VPWR
+ _0177_ VGND net172 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit2.Q
+ sg13g2_o21ai_1
X_0595_ _0148_ _0150_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S4BEG2
+ VPWR VGND sg13g2_nor2_1
X_1216_ net220 net730 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
X_1147_ net788 net654 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
X_1078_ net783 net679 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_43_112 VPWR VGND sg13g2_fill_1
XFILLER_43_134 VPWR VGND sg13g2_fill_1
XFILLER_61_86 VPWR VGND sg13g2_fill_2
XFILLER_43_156 VPWR VGND sg13g2_fill_2
X_0380_ VGND VPWR _0071_ _0072_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit31.Q
+ _0005_ _0073_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit30.Q
+ sg13g2_a221oi_1
XIHP_SRAM_583 VPWR VGND TIE_HIGH_SRAM sg13g2_tiehi
X_1001_ net800 net697 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_34_123 VPWR VGND sg13g2_fill_1
X_0578_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit20.Q _0135_
+ _0136_ VPWR VGND sg13g2_nor2_1
X_0716_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit26.Q net145
+ net187 net180 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG15
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit27.Q net268 VPWR
+ VGND sg13g2_mux4_1
X_0647_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit28.Q net225
+ net245 _0067_ net140 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit29.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG10 VPWR VGND sg13g2_mux4_1
X_1696_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb5 net550 VPWR
+ VGND sg13g2_buf_1
XFILLER_25_178 VPWR VGND sg13g2_fill_2
Xinput123 Tile_X0Y0_S2END[5] net123 VPWR VGND sg13g2_buf_1
Xinput134 Tile_X0Y0_S4END[0] net134 VPWR VGND sg13g2_buf_1
Xinput101 Tile_X0Y0_FrameData[27] net101 VPWR VGND sg13g2_buf_1
Xinput112 Tile_X0Y0_FrameData[8] net112 VPWR VGND sg13g2_buf_1
Xinput145 Tile_X0Y1_E1END[3] net145 VPWR VGND sg13g2_buf_1
Xinput156 Tile_X0Y1_E2MID[2] net156 VPWR VGND sg13g2_buf_1
Xinput178 Tile_X0Y1_EE4END[13] net178 VPWR VGND sg13g2_buf_1
Xinput167 Tile_X0Y1_E6END[3] net167 VPWR VGND sg13g2_buf_1
Xinput189 Tile_X0Y1_EE4END[9] net189 VPWR VGND sg13g2_buf_1
XFILLER_75_8 VPWR VGND sg13g2_fill_2
X_0501_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit14.Q net66
+ net80 net64 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG8 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit15.Q
+ net311 VPWR VGND sg13g2_mux4_1
X_0432_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit31.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END0
+ net12 net114 net18 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit30.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W1BEG0 VPWR VGND sg13g2_mux4_1
X_1481_ net784 net357 VPWR VGND sg13g2_buf_1
X_1550_ Tile_X0Y1_N4END[12] net410 VPWR VGND sg13g2_buf_1
X_0363_ net224 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit26.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit27.Q _0062_ VPWR
+ VGND sg13g2_nor3_1
XFILLER_94_0 VPWR VGND sg13g2_fill_1
Xfanout813 net82 net813 VPWR VGND sg13g2_buf_1
Xfanout802 net93 net802 VPWR VGND sg13g2_buf_1
X_1679_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W1BEG0 net533 VPWR
+ VGND sg13g2_buf_1
XFILLER_3_27 VPWR VGND sg13g2_decap_8
XFILLER_67_63 VPWR VGND sg13g2_decap_8
XFILLER_83_84 VPWR VGND sg13g2_fill_2
X_0981_ net782 net708 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
Xoutput416 net416 Tile_X0Y0_UserCLKo VPWR VGND sg13g2_buf_1
Xoutput405 net405 Tile_X0Y0_N4BEG[14] VPWR VGND sg13g2_buf_1
X_1602_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG7 net462 VPWR
+ VGND sg13g2_buf_1
XFILLER_8_152 VPWR VGND sg13g2_fill_1
Xoutput438 net438 Tile_X0Y0_W6BEG[10] VPWR VGND sg13g2_buf_1
X_1533_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG3 net387 VPWR
+ VGND sg13g2_buf_1
Xoutput449 net449 Tile_X0Y0_WW4BEG[0] VPWR VGND sg13g2_buf_1
Xoutput427 net427 Tile_X0Y0_W2BEG[6] VPWR VGND sg13g2_buf_1
X_0415_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit20.Q net241
+ net233 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG6 net132 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit21.Q
+ _0083_ VPWR VGND sg13g2_mux4_1
X_1464_ net774 net646 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
X_1395_ net768 net658 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
X_0346_ _0046_ _0045_ net150 net129 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit30.Q
+ VPWR VGND sg13g2_a22oi_1
Xfanout654 net656 net654 VPWR VGND sg13g2_buf_1
Xfanout665 net667 net665 VPWR VGND sg13g2_buf_1
XFILLER_85_140 VPWR VGND sg13g2_fill_1
Xfanout698 net699 net698 VPWR VGND sg13g2_buf_1
Xfanout676 net677 net676 VPWR VGND sg13g2_buf_1
Xfanout687 net689 net687 VPWR VGND sg13g2_buf_1
XFILLER_77_129 VPWR VGND sg13g2_fill_2
Xfanout643 net646 net643 VPWR VGND sg13g2_buf_1
Xfanout632 _0084_ net632 VPWR VGND sg13g2_buf_1
XFILLER_68_129 VPWR VGND sg13g2_fill_2
X_1180_ net778 net740 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
X_0964_ net100 net712 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
X_0895_ net106 net734 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
X_1516_ Tile_X0Y1_FrameStrobe[10] net361 VPWR VGND sg13g2_buf_1
Xoutput257 net257 ADDR_SRAM6 VPWR VGND sg13g2_buf_1
Xoutput268 net268 BM_SRAM15 VPWR VGND sg13g2_buf_1
X_1378_ net753 net671 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
X_0329_ VPWR _0032_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit13.Q
+ VGND sg13g2_inv_1
Xoutput279 net279 BM_SRAM25 VPWR VGND sg13g2_buf_1
X_1447_ net770 net647 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_2_147 VPWR VGND sg13g2_decap_8
XFILLER_64_64 VPWR VGND sg13g2_fill_1
XFILLER_64_53 VPWR VGND sg13g2_decap_8
XFILLER_58_162 VPWR VGND sg13g2_decap_4
XFILLER_48_65 VPWR VGND sg13g2_decap_8
XFILLER_73_198 VPWR VGND sg13g2_fill_2
X_0680_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit17.Q net25
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG4 _0161_ net632
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit16.Q Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG11
+ VPWR VGND sg13g2_mux4_1
X_1301_ net771 net693 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
X_1232_ net206 net714 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
X_1094_ net98 net665 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
X_1163_ net211 net741 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
X_0947_ net84 net722 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_118_167 VPWR VGND sg13g2_decap_8
X_0878_ net806 net744 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_70_146 VPWR VGND sg13g2_fill_1
XFILLER_75_96 VPWR VGND sg13g2_fill_1
XFILLER_61_146 VPWR VGND sg13g2_decap_4
XFILLER_91_84 VPWR VGND sg13g2_fill_2
X_0801_ _0238_ VPWR _0239_ VGND _0031_ _0159_ sg13g2_o21ai_1
XFILLER_115_159 VPWR VGND sg13g2_decap_4
X_0594_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit26.Q _0149_
+ _0150_ VPWR VGND sg13g2_nor2_1
X_0732_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit26.Q net145
+ net187 net180 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG15
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit27.Q net301 VPWR
+ VGND sg13g2_mux4_1
X_0663_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit12.Q net225
+ net245 _0067_ net140 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit13.Q
+ _0159_ VPWR VGND sg13g2_mux4_1
X_1146_ net787 net652 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_1_60 VPWR VGND sg13g2_decap_8
XFILLER_1_71 VPWR VGND sg13g2_fill_2
X_1215_ net221 net727 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
X_1077_ net782 net679 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_106_126 VPWR VGND sg13g2_fill_1
XFILLER_121_129 VPWR VGND sg13g2_decap_8
XFILLER_29_67 VPWR VGND sg13g2_fill_2
XFILLER_45_33 VPWR VGND sg13g2_fill_1
XFILLER_61_65 VPWR VGND sg13g2_decap_4
XFILLER_6_16 VPWR VGND sg13g2_fill_1
XFILLER_112_129 VPWR VGND sg13g2_fill_2
XFILLER_6_27 VPWR VGND sg13g2_fill_1
X_1000_ net799 net700 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_19_121 VPWR VGND sg13g2_decap_4
XFILLER_19_165 VPWR VGND sg13g2_fill_1
X_0715_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit24.Q net144
+ net186 net179 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG14
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit25.Q net267 VPWR
+ VGND sg13g2_mux4_1
XFILLER_103_107 VPWR VGND sg13g2_fill_2
X_0577_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit18.Q net34
+ net69 net60 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit19.Q
+ _0135_ VPWR VGND sg13g2_mux4_1
X_0646_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit2.Q net28
+ net32 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG11 net637
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit3.Q Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG4
+ VPWR VGND sg13g2_mux4_1
X_1695_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb4 net549 VPWR
+ VGND sg13g2_buf_1
X_1129_ net800 net655 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_15_47 VPWR VGND sg13g2_fill_1
Xinput135 Tile_X0Y0_S4END[1] net135 VPWR VGND sg13g2_buf_1
Xinput124 Tile_X0Y0_S2END[6] net124 VPWR VGND sg13g2_buf_1
Xinput102 Tile_X0Y0_FrameData[28] net102 VPWR VGND sg13g2_buf_1
Xinput113 Tile_X0Y0_FrameData[9] net113 VPWR VGND sg13g2_buf_1
Xinput157 Tile_X0Y1_E2MID[3] net157 VPWR VGND sg13g2_buf_1
Xinput146 Tile_X0Y1_E2END[0] net146 VPWR VGND sg13g2_buf_1
Xinput179 Tile_X0Y1_EE4END[14] net179 VPWR VGND sg13g2_buf_1
Xinput168 Tile_X0Y1_E6END[4] net168 VPWR VGND sg13g2_buf_1
XFILLER_56_10 VPWR VGND sg13g2_fill_1
XFILLER_56_32 VPWR VGND sg13g2_fill_1
XFILLER_72_75 VPWR VGND sg13g2_fill_1
XFILLER_31_105 VPWR VGND sg13g2_fill_1
XFILLER_31_127 VPWR VGND sg13g2_fill_2
XFILLER_72_97 VPWR VGND sg13g2_decap_8
X_0500_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit12.Q net79
+ net72 net63 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG7 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit13.Q
+ net310 VPWR VGND sg13g2_mux4_1
XFILLER_97_83 VPWR VGND sg13g2_fill_1
X_1480_ net785 net356 VPWR VGND sg13g2_buf_1
X_0362_ _0061_ _0060_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit26.Q
+ VPWR VGND sg13g2_nand2b_1
X_0431_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit11.Q net142
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG12 net168 _0091_
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit10.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END0
+ VPWR VGND sg13g2_mux4_1
XFILLER_11_4 VPWR VGND sg13g2_fill_2
XFILLER_87_0 VPWR VGND sg13g2_fill_1
X_1678_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S4BEG3 net523 VPWR
+ VGND sg13g2_buf_1
Xfanout803 net92 net803 VPWR VGND sg13g2_buf_1
X_0629_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit2.Q net28
+ net6 net637 net635 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit3.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG4 VPWR VGND sg13g2_mux4_1
X_0980_ net83 net712 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_16_90 VPWR VGND sg13g2_fill_2
Xoutput406 net406 Tile_X0Y0_N4BEG[15] VPWR VGND sg13g2_buf_1
Xoutput439 net439 Tile_X0Y0_W6BEG[11] VPWR VGND sg13g2_buf_1
X_1532_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG2 net386 VPWR
+ VGND sg13g2_buf_1
X_1601_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG6 net461 VPWR
+ VGND sg13g2_buf_1
Xoutput428 net428 Tile_X0Y0_W2BEG[7] VPWR VGND sg13g2_buf_1
Xoutput417 net417 Tile_X0Y0_W1BEG[0] VPWR VGND sg13g2_buf_1
X_0414_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit14.Q net36
+ net47 net39 net624 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit15.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG6 VPWR VGND sg13g2_mux4_1
X_1463_ net773 net646 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
X_1394_ net767 net658 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
X_0345_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit29.Q Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit30.Q
+ _0045_ VPWR VGND sg13g2_nor2_1
XFILLER_94_196 VPWR VGND sg13g2_fill_1
XFILLER_10_108 VPWR VGND sg13g2_decap_8
Xfanout633 _0083_ net633 VPWR VGND sg13g2_buf_1
Xfanout644 net645 net644 VPWR VGND sg13g2_buf_1
Xfanout655 net656 net655 VPWR VGND sg13g2_buf_1
Xfanout666 net667 net666 VPWR VGND sg13g2_buf_1
Xfanout677 net678 net677 VPWR VGND sg13g2_buf_1
Xfanout699 net702 net699 VPWR VGND sg13g2_buf_1
Xfanout688 net689 net688 VPWR VGND sg13g2_buf_1
XFILLER_53_66 VPWR VGND sg13g2_fill_1
XFILLER_68_108 VPWR VGND sg13g2_decap_4
XFILLER_94_84 VPWR VGND sg13g2_fill_1
XFILLER_32_200 VPWR VGND sg13g2_fill_1
X_0963_ net101 net712 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
X_0894_ net813 net743 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
X_1515_ net644 net379 VPWR VGND sg13g2_buf_1
Xoutput258 net258 ADDR_SRAM7 VPWR VGND sg13g2_buf_1
Xoutput269 net269 BM_SRAM16 VPWR VGND sg13g2_buf_1
XFILLER_67_196 VPWR VGND sg13g2_fill_1
X_1377_ net752 net671 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
X_1446_ net759 net650 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
X_0328_ VPWR _0031_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit12.Q
+ VGND sg13g2_inv_1
XFILLER_2_126 VPWR VGND sg13g2_decap_8
X_1162_ net213 net740 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
X_1300_ net769 net693 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
X_1231_ net207 net714 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_49_163 VPWR VGND sg13g2_fill_1
X_1093_ net99 net665 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_118_146 VPWR VGND sg13g2_decap_8
X_0946_ net85 net720 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
X_0877_ net805 net744 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
X_1429_ net200 net650 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_55_133 VPWR VGND sg13g2_fill_2
XFILLER_50_12 VPWR VGND sg13g2_fill_2
XFILLER_115_82 VPWR VGND sg13g2_fill_1
XFILLER_46_100 VPWR VGND sg13g2_fill_1
XFILLER_61_103 VPWR VGND sg13g2_decap_8
XFILLER_46_199 VPWR VGND sg13g2_fill_2
X_0800_ VPWR _0238_ _0237_ VGND sg13g2_inv_1
X_0731_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit24.Q net144
+ net186 net179 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG14
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit25.Q net300 VPWR
+ VGND sg13g2_mux4_1
X_0593_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit25.Q net36
+ net62 net71 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG2 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit24.Q
+ _0149_ VPWR VGND sg13g2_mux4_1
X_0662_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit18.Q net2
+ net6 _0158_ net637 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit19.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG12 VPWR VGND sg13g2_mux4_1
X_1145_ net786 net652 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
X_1214_ net780 net726 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
X_1076_ net812 net677 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
X_0929_ net792 net720 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_121_108 VPWR VGND sg13g2_decap_8
XFILLER_101_62 VPWR VGND sg13g2_fill_1
XFILLER_120_174 VPWR VGND sg13g2_decap_8
XFILLER_86_85 VPWR VGND sg13g2_fill_1
XFILLER_13_8 VPWR VGND sg13g2_fill_2
XFILLER_19_199 VPWR VGND sg13g2_fill_2
X_0714_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit22.Q net143
+ net185 net178 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG13
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit23.Q net266 VPWR
+ VGND sg13g2_mux4_1
X_1694_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb3 net548 VPWR
+ VGND sg13g2_buf_1
X_0645_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit30.Q net226
+ net246 _0074_ net141 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit31.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG11 VPWR VGND sg13g2_mux4_1
X_0576_ VGND VPWR _0015_ _0130_ _0134_ _0133_ sg13g2_a21oi_1
XFILLER_32_0 VPWR VGND sg13g2_fill_2
X_1128_ net96 net655 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
X_1059_ net794 net677 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
Xinput125 Tile_X0Y0_S2END[7] net125 VPWR VGND sg13g2_buf_1
Xinput114 Tile_X0Y0_S1END[0] net114 VPWR VGND sg13g2_buf_1
Xinput136 Tile_X0Y0_S4END[2] net136 VPWR VGND sg13g2_buf_1
Xinput103 Tile_X0Y0_FrameData[29] net103 VPWR VGND sg13g2_buf_1
Xinput158 Tile_X0Y1_E2MID[4] net158 VPWR VGND sg13g2_buf_1
Xinput147 Tile_X0Y1_E2END[1] net147 VPWR VGND sg13g2_buf_1
Xinput169 Tile_X0Y1_E6END[5] net169 VPWR VGND sg13g2_buf_1
XFILLER_56_99 VPWR VGND sg13g2_decap_4
X_0361_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit28.Q net35
+ net65 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG13 _0059_
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit29.Q _0060_ VPWR
+ VGND sg13g2_mux4_1
X_0430_ VGND VPWR _0090_ _0089_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit25.Q
+ _0010_ _0091_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit24.Q
+ sg13g2_a221oi_1
XFILLER_117_39 VPWR VGND sg13g2_decap_8
Xfanout804 net91 net804 VPWR VGND sg13g2_buf_1
X_0628_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit0.Q net25
+ net5 net637 net636 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit1.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG3 VPWR VGND sg13g2_mux4_1
X_1677_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S4BEG2 net522 VPWR
+ VGND sg13g2_buf_1
X_0559_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit22.Q VPWR
+ _0119_ VGND _0117_ _0118_ sg13g2_o21ai_1
XFILLER_21_194 VPWR VGND sg13g2_fill_2
XFILLER_107_94 VPWR VGND sg13g2_decap_8
XFILLER_88_194 VPWR VGND sg13g2_fill_2
XFILLER_67_21 VPWR VGND sg13g2_decap_4
XFILLER_12_172 VPWR VGND sg13g2_fill_2
Xoutput407 net407 Tile_X0Y0_N4BEG[1] VPWR VGND sg13g2_buf_1
X_1531_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG1 net385 VPWR
+ VGND sg13g2_buf_1
X_1600_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG5 net460 VPWR
+ VGND sg13g2_buf_1
Xoutput429 net429 Tile_X0Y0_W2BEGb[0] VPWR VGND sg13g2_buf_1
Xoutput418 net418 Tile_X0Y0_W1BEG[1] VPWR VGND sg13g2_buf_1
X_1462_ net772 net641 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
X_0413_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit8.Q net48
+ net40 net58 net625 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit9.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG5 VPWR VGND sg13g2_mux4_1
X_0344_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit29.Q VPWR
+ _0044_ VGND Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit30.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG0 sg13g2_o21ai_1
X_1393_ net766 net661 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
Xfanout656 net657 net656 VPWR VGND sg13g2_buf_1
Xfanout623 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG7 net623
+ VPWR VGND sg13g2_buf_1
Xfanout667 net668 net667 VPWR VGND sg13g2_buf_1
Xfanout645 net646 net645 VPWR VGND sg13g2_buf_1
Xfanout634 _0082_ net634 VPWR VGND sg13g2_buf_1
Xfanout689 net690 net689 VPWR VGND sg13g2_buf_1
Xfanout678 Tile_X0Y1_FrameStrobe[6] net678 VPWR VGND sg13g2_buf_1
XFILLER_53_23 VPWR VGND sg13g2_fill_1
X_0962_ net102 net712 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
X_0893_ net802 net743 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
X_1514_ net654 net378 VPWR VGND sg13g2_buf_1
Xoutput259 net259 ADDR_SRAM8 VPWR VGND sg13g2_buf_1
X_1445_ net756 net649 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
X_1376_ net751 net670 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
X_0327_ VPWR _0030_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit10.Q
+ VGND sg13g2_inv_1
XFILLER_2_105 VPWR VGND sg13g2_decap_8
XFILLER_73_145 VPWR VGND sg13g2_fill_2
XFILLER_120_83 VPWR VGND sg13g2_decap_8
XFILLER_80_43 VPWR VGND sg13g2_fill_2
XFILLER_80_21 VPWR VGND sg13g2_fill_1
XFILLER_89_74 VPWR VGND sg13g2_fill_1
XFILLER_43_8 VPWR VGND sg13g2_fill_2
X_1092_ net100 net665 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_1_193 VPWR VGND sg13g2_decap_8
X_1161_ net214 net740 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
X_1230_ net763 net717 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_118_125 VPWR VGND sg13g2_decap_8
X_0945_ net86 net720 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
X_0876_ net804 net743 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_62_0 VPWR VGND sg13g2_decap_8
X_1428_ net769 net651 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
X_1359_ net764 net673 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_109_169 VPWR VGND sg13g2_fill_2
XFILLER_1_4 VPWR VGND sg13g2_fill_1
XFILLER_91_31 VPWR VGND sg13g2_fill_1
X_0730_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit22.Q net143
+ net185 net178 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG13
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit23.Q net299 VPWR
+ VGND sg13g2_mux4_1
X_0661_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit14.Q net226
+ net246 _0074_ net141 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit15.Q
+ _0158_ VPWR VGND sg13g2_mux4_1
X_0592_ VGND VPWR _0017_ _0144_ _0148_ _0147_ sg13g2_a21oi_1
X_1213_ net779 net726 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
X_1075_ net811 net677 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
X_1144_ net785 net652 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_37_112 VPWR VGND sg13g2_fill_2
XFILLER_60_192 VPWR VGND sg13g2_fill_1
X_0928_ net790 net722 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
X_0859_ net149 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit5.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit6.Q _0294_ VPWR
+ VGND sg13g2_nor3_1
XFILLER_29_47 VPWR VGND sg13g2_fill_2
XFILLER_120_153 VPWR VGND sg13g2_decap_8
XFILLER_103_109 VPWR VGND sg13g2_fill_1
X_1693_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb2 net547 VPWR
+ VGND sg13g2_buf_1
X_0644_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit0.Q net25
+ net9 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG12 net635 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit1.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG3 VPWR VGND sg13g2_mux4_1
X_0713_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit20.Q net142
+ net184 net177 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG12
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit21.Q net265 VPWR
+ VGND sg13g2_mux4_1
X_0575_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit20.Q VPWR
+ _0133_ VGND _0131_ _0132_ sg13g2_o21ai_1
X_1127_ net97 net654 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
X_1058_ net793 net678 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_40_118 VPWR VGND sg13g2_decap_8
XFILLER_31_37 VPWR VGND sg13g2_fill_2
Xinput126 Tile_X0Y0_S2MID[0] net126 VPWR VGND sg13g2_buf_1
Xinput115 Tile_X0Y0_S1END[1] net115 VPWR VGND sg13g2_buf_1
Xinput104 Tile_X0Y0_FrameData[2] net104 VPWR VGND sg13g2_buf_1
Xinput137 Tile_X0Y0_S4END[3] net137 VPWR VGND sg13g2_buf_1
Xinput159 Tile_X0Y1_E2MID[5] net159 VPWR VGND sg13g2_buf_1
Xinput148 Tile_X0Y1_E2END[2] net148 VPWR VGND sg13g2_buf_1
XFILLER_72_22 VPWR VGND sg13g2_fill_1
X_0360_ VGND VPWR _0057_ _0058_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit27.Q
+ _0003_ _0059_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit26.Q
+ sg13g2_a221oi_1
XFILLER_11_6 VPWR VGND sg13g2_fill_1
X_0558_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit21.Q VPWR
+ _0118_ VGND Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit20.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG14 sg13g2_o21ai_1
Xfanout805 net90 net805 VPWR VGND sg13g2_buf_1
X_0627_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit30.Q net14
+ net4 net638 net634 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit31.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG2 VPWR VGND sg13g2_mux4_1
X_1676_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S4BEG1 net521 VPWR
+ VGND sg13g2_buf_1
X_0489_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit23.Q net10
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG7 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG3
+ net626 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit22.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG8
+ VPWR VGND sg13g2_mux4_1
XFILLER_26_37 VPWR VGND sg13g2_fill_2
XFILLER_88_162 VPWR VGND sg13g2_fill_1
Xoutput408 net408 Tile_X0Y0_N4BEG[2] VPWR VGND sg13g2_buf_1
X_1530_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG0 net384 VPWR
+ VGND sg13g2_buf_1
Xoutput419 net419 Tile_X0Y0_W1BEG[2] VPWR VGND sg13g2_buf_1
X_0412_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit19.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb5
+ net131 net240 net123 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit18.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG5 VPWR VGND sg13g2_mux4_1
X_1392_ net765 net659 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
X_1461_ net771 net641 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
X_0343_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit9.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb0
+ net126 net235 net118 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit8.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG0 VPWR VGND sg13g2_mux4_1
Xfanout624 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG6 net624
+ VPWR VGND sg13g2_buf_1
Xfanout657 net222 net657 VPWR VGND sg13g2_buf_1
Xfanout679 Tile_X0Y1_FrameStrobe[6] net679 VPWR VGND sg13g2_buf_1
Xfanout668 Tile_X0Y1_FrameStrobe[7] net668 VPWR VGND sg13g2_buf_1
Xfanout646 Tile_X0Y1_FrameStrobe[9] net646 VPWR VGND sg13g2_buf_1
X_1659_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG4 net513 VPWR
+ VGND sg13g2_buf_1
Xfanout635 net636 net635 VPWR VGND sg13g2_buf_1
XFILLER_118_83 VPWR VGND sg13g2_decap_8
XFILLER_78_21 VPWR VGND sg13g2_fill_2
X_0961_ net103 net712 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
X_0892_ net791 net744 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
X_1513_ net667 net377 VPWR VGND sg13g2_buf_1
XFILLER_4_73 VPWR VGND sg13g2_decap_8
X_1375_ net750 net670 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
X_1444_ net755 net649 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_82_113 VPWR VGND sg13g2_fill_2
X_0326_ VPWR _0029_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit9.Q
+ VGND sg13g2_inv_1
XFILLER_120_62 VPWR VGND sg13g2_decap_8
XFILLER_80_88 VPWR VGND sg13g2_fill_2
XFILLER_1_172 VPWR VGND sg13g2_decap_8
X_1091_ net794 net664 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
X_1160_ net799 net645 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_118_104 VPWR VGND sg13g2_decap_8
X_0944_ net808 net723 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
X_0875_ net803 net743 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
X_1427_ net768 net651 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
X_1358_ net763 net670 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
X_0309_ VPWR _0012_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit18.Q
+ VGND sg13g2_inv_1
X_1289_ net757 net695 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_59_67 VPWR VGND sg13g2_fill_2
Xoutput580 net580 Tile_X0Y1_WW4BEG[9] VPWR VGND sg13g2_buf_1
XFILLER_115_95 VPWR VGND sg13g2_fill_1
XFILLER_46_146 VPWR VGND sg13g2_fill_2
X_0591_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit26.Q VPWR
+ _0147_ VGND _0145_ _0146_ sg13g2_o21ai_1
X_0660_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit16.Q net31
+ net5 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG4 net635 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit17.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG11 VPWR VGND sg13g2_mux4_1
X_1212_ net778 net725 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_27_4 VPWR VGND sg13g2_fill_2
X_1074_ net810 net676 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
X_1143_ net784 net652 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_52_127 VPWR VGND sg13g2_fill_2
X_0927_ net789 net722 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_60_171 VPWR VGND sg13g2_decap_4
XFILLER_20_17 VPWR VGND sg13g2_fill_1
XFILLER_20_39 VPWR VGND sg13g2_fill_1
X_0789_ VPWR _0228_ _0227_ VGND sg13g2_inv_1
X_0858_ VGND VPWR net128 _0037_ _0293_ _0292_ sg13g2_a21oi_1
XFILLER_43_105 VPWR VGND sg13g2_decap_8
XFILLER_120_132 VPWR VGND sg13g2_decap_8
XFILLER_10_61 VPWR VGND sg13g2_decap_4
X_0574_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit19.Q VPWR
+ _0132_ VGND Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit18.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG12 sg13g2_o21ai_1
X_1692_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb1 net546 VPWR
+ VGND sg13g2_buf_1
X_0643_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit30.Q net14
+ net8 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG13 net634 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit31.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG2 VPWR VGND sg13g2_mux4_1
X_0712_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit18.Q net183
+ net176 net164 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG11
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit19.Q net264 VPWR
+ VGND sg13g2_mux4_1
XFILLER_111_198 VPWR VGND sg13g2_fill_2
X_1126_ net797 net654 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_18_0 VPWR VGND sg13g2_fill_1
X_1057_ net792 net678 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
Xinput116 Tile_X0Y0_S1END[2] net116 VPWR VGND sg13g2_buf_1
Xinput138 Tile_X0Y0_S4END[4] net138 VPWR VGND sg13g2_buf_1
Xinput127 Tile_X0Y0_S2MID[1] net127 VPWR VGND sg13g2_buf_1
Xinput105 Tile_X0Y0_FrameData[30] net105 VPWR VGND sg13g2_buf_1
Xinput149 Tile_X0Y1_E2END[3] net149 VPWR VGND sg13g2_buf_1
XFILLER_102_198 VPWR VGND sg13g2_fill_2
XFILLER_62_200 VPWR VGND sg13g2_fill_1
X_0557_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG2 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit20.Q
+ _0117_ VPWR VGND sg13g2_nor2b_1
Xfanout806 net89 net806 VPWR VGND sg13g2_buf_1
X_0626_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit28.Q net3
+ net33 net639 net633 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit29.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG1 VPWR VGND sg13g2_mux4_1
X_1675_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S4BEG0 net520 VPWR
+ VGND sg13g2_buf_1
X_1109_ net782 net666 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
X_0488_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit20.Q net18
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG4 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG8
+ net628 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit21.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG7
+ VPWR VGND sg13g2_mux4_1
XFILLER_21_196 VPWR VGND sg13g2_fill_1
XFILLER_88_196 VPWR VGND sg13g2_fill_1
XFILLER_44_200 VPWR VGND sg13g2_fill_1
XFILLER_66_8 VPWR VGND sg13g2_fill_1
XFILLER_8_178 VPWR VGND sg13g2_fill_2
XFILLER_8_112 VPWR VGND sg13g2_decap_4
Xoutput409 net409 Tile_X0Y0_N4BEG[3] VPWR VGND sg13g2_buf_1
X_1391_ net764 net659 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
X_1460_ net202 net641 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
X_0342_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit18.Q net161
+ net153 net171 net640 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit19.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb0 VPWR VGND sg13g2_mux4_1
X_0411_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit29.Q net156
+ net166 net148 _0082_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit28.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb5 VPWR VGND sg13g2_mux4_1
XFILLER_35_200 VPWR VGND sg13g2_fill_1
X_1658_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG3 net512 VPWR
+ VGND sg13g2_buf_1
X_1589_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG6 net445 VPWR
+ VGND sg13g2_buf_1
Xfanout625 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG5 net625
+ VPWR VGND sg13g2_buf_1
Xfanout636 _0081_ net636 VPWR VGND sg13g2_buf_1
Xfanout658 net661 net658 VPWR VGND sg13g2_buf_1
Xfanout669 net672 net669 VPWR VGND sg13g2_buf_1
X_0609_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit14.Q net142
+ net172 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG12 _0091_
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit15.Q Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S1BEG0
+ VPWR VGND sg13g2_mux4_1
Xfanout647 net651 net647 VPWR VGND sg13g2_buf_1
XFILLER_118_62 VPWR VGND sg13g2_decap_4
XFILLER_76_199 VPWR VGND sg13g2_fill_2
X_0960_ net790 net709 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
X_0891_ net788 net747 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
X_1512_ net678 net376 VPWR VGND sg13g2_buf_1
X_1374_ net780 net669 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_4_41 VPWR VGND sg13g2_decap_8
X_1443_ net754 net648 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
X_0325_ VPWR _0028_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit7.Q
+ VGND sg13g2_inv_1
XFILLER_90_191 VPWR VGND sg13g2_fill_2
XFILLER_58_166 VPWR VGND sg13g2_fill_2
XFILLER_58_155 VPWR VGND sg13g2_decap_8
XFILLER_58_133 VPWR VGND sg13g2_fill_1
XFILLER_120_41 VPWR VGND sg13g2_decap_8
XFILLER_80_45 VPWR VGND sg13g2_fill_1
XFILLER_64_46 VPWR VGND sg13g2_decap_8
XFILLER_1_151 VPWR VGND sg13g2_decap_8
X_1090_ net793 net664 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_64_103 VPWR VGND sg13g2_fill_1
XFILLER_49_199 VPWR VGND sg13g2_fill_2
X_0943_ net807 net723 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
X_0874_ net801 net744 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
X_0308_ VPWR _0011_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit15.Q
+ VGND sg13g2_inv_1
X_1357_ net762 net669 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
X_1426_ net204 net647 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
X_1288_ net781 net703 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_34_49 VPWR VGND sg13g2_fill_2
Xoutput581 net581 WEN_SRAM VPWR VGND sg13g2_buf_1
Xoutput570 net570 Tile_X0Y1_WW4BEG[14] VPWR VGND sg13g2_buf_1
XFILLER_75_56 VPWR VGND sg13g2_fill_2
XFILLER_61_139 VPWR VGND sg13g2_decap_8
XFILLER_61_117 VPWR VGND sg13g2_decap_4
X_0590_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit25.Q VPWR
+ _0146_ VGND Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit24.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG14 sg13g2_o21ai_1
X_1142_ net783 net652 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
X_1211_ net777 net725 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_1_20 VPWR VGND sg13g2_fill_1
XFILLER_1_53 VPWR VGND sg13g2_decap_8
XFILLER_37_114 VPWR VGND sg13g2_fill_1
X_1073_ net809 net675 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
X_0926_ net82 net732 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
X_0857_ VGND VPWR _0001_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit5.Q
+ _0292_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit6.Q sg13g2_a21oi_1
X_0788_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit10.Q VPWR
+ _0227_ VGND net169 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit9.Q
+ sg13g2_o21ai_1
XFILLER_29_49 VPWR VGND sg13g2_fill_1
X_1409_ net219 net662 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_61_69 VPWR VGND sg13g2_fill_1
XFILLER_61_58 VPWR VGND sg13g2_decap_8
XFILLER_120_111 VPWR VGND sg13g2_decap_8
XFILLER_19_82 VPWR VGND sg13g2_fill_1
X_1691_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb0 net545 VPWR
+ VGND sg13g2_buf_1
X_0711_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit16.Q net182
+ net175 net163 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG10
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit17.Q net263 VPWR
+ VGND sg13g2_mux4_1
X_0573_ net626 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit18.Q
+ _0131_ VPWR VGND sg13g2_nor2b_1
X_0642_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit28.Q net3
+ net7 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG14 net633 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit29.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG1 VPWR VGND sg13g2_mux4_1
X_1125_ net99 net654 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
X_1056_ net790 net675 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_15_29 VPWR VGND sg13g2_fill_1
XFILLER_40_109 VPWR VGND sg13g2_fill_1
X_0909_ net805 net731 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
Xinput139 Tile_X0Y0_S4END[5] net139 VPWR VGND sg13g2_buf_1
Xinput128 Tile_X0Y0_S2MID[2] net128 VPWR VGND sg13g2_buf_1
Xinput117 Tile_X0Y0_S1END[3] net117 VPWR VGND sg13g2_buf_1
Xinput106 Tile_X0Y0_FrameData[31] net106 VPWR VGND sg13g2_buf_1
XFILLER_62_90 VPWR VGND sg13g2_fill_1
X_1674_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S4BEG3 net519 VPWR
+ VGND sg13g2_buf_1
X_0625_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit26.Q net2
+ net32 net640 net632 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit27.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG0 VPWR VGND sg13g2_mux4_1
XFILLER_7_41 VPWR VGND sg13g2_fill_1
X_0556_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG6 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG10
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit20.Q _0116_ VPWR
+ VGND sg13g2_mux2_1
X_0487_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit18.Q net17
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG5 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG9
+ net629 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit19.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG6
+ VPWR VGND sg13g2_mux4_1
Xfanout807 net88 net807 VPWR VGND sg13g2_buf_1
XFILLER_30_0 VPWR VGND sg13g2_fill_1
X_1039_ net807 net685 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
X_1108_ net812 net663 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_83_56 VPWR VGND sg13g2_fill_2
X_0410_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit18.Q net240
+ net232 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG5 net131 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit19.Q
+ _0082_ VPWR VGND sg13g2_mux4_1
X_1390_ net763 net658 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
X_0341_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit8.Q net235
+ net227 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG0 net126 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit9.Q
+ _0043_ VPWR VGND sg13g2_mux4_1
X_1588_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG5 net444 VPWR
+ VGND sg13g2_buf_1
X_1657_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG2 net511 VPWR
+ VGND sg13g2_buf_1
X_0608_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit23.Q net34
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG12 net60 _0087_
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit22.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1BEG0
+ VPWR VGND sg13g2_mux4_1
X_1726_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG15 net571 VPWR
+ VGND sg13g2_buf_1
X_0539_ VGND VPWR Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit6.Q
+ _0100_ _0101_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit7.Q
+ net260 _0042_ sg13g2_a221oi_1
Xfanout626 net627 net626 VPWR VGND sg13g2_buf_1
Xfanout659 net660 net659 VPWR VGND sg13g2_buf_1
Xfanout648 net651 net648 VPWR VGND sg13g2_buf_1
Xfanout637 _0080_ net637 VPWR VGND sg13g2_buf_1
XFILLER_118_41 VPWR VGND sg13g2_decap_8
XFILLER_78_23 VPWR VGND sg13g2_fill_1
XFILLER_76_123 VPWR VGND sg13g2_fill_2
XFILLER_91_148 VPWR VGND sg13g2_fill_2
X_0890_ net787 net746 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
X_1511_ net687 net375 VPWR VGND sg13g2_buf_1
XFILLER_4_171 VPWR VGND sg13g2_decap_8
XFILLER_4_20 VPWR VGND sg13g2_decap_8
X_1442_ net753 net648 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_82_115 VPWR VGND sg13g2_fill_1
X_1373_ net779 net669 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
X_0324_ VPWR _0027_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit6.Q
+ VGND sg13g2_inv_1
XFILLER_2_119 VPWR VGND sg13g2_decap_8
X_1709_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG10 net554 VPWR
+ VGND sg13g2_buf_1
XFILLER_120_97 VPWR VGND sg13g2_decap_8
XFILLER_120_20 VPWR VGND sg13g2_decap_8
XFILLER_81_170 VPWR VGND sg13g2_fill_1
XFILLER_8_0 VPWR VGND sg13g2_fill_2
XFILLER_118_139 VPWR VGND sg13g2_decap_8
X_0942_ net806 net721 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
X_0873_ net800 net744 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
X_1425_ net205 net647 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_70_107 VPWR VGND sg13g2_decap_4
X_1356_ net761 net671 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_18_18 VPWR VGND sg13g2_fill_1
X_0307_ VPWR _0010_ net162 VGND sg13g2_inv_1
X_1287_ net770 net703 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_117_183 VPWR VGND sg13g2_decap_4
XFILLER_117_161 VPWR VGND sg13g2_decap_4
XFILLER_59_69 VPWR VGND sg13g2_fill_1
Xoutput571 net571 Tile_X0Y1_WW4BEG[15] VPWR VGND sg13g2_buf_1
Xoutput560 net560 Tile_X0Y1_W6BEG[5] VPWR VGND sg13g2_buf_1
XFILLER_108_150 VPWR VGND sg13g2_fill_1
XFILLER_40_82 VPWR VGND sg13g2_fill_1
X_1141_ net782 net652 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
X_1072_ net808 net678 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_27_6 VPWR VGND sg13g2_fill_1
X_1210_ net195 net728 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_52_129 VPWR VGND sg13g2_fill_1
X_0925_ net93 net732 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_60_0 VPWR VGND sg13g2_decap_4
X_0787_ VGND VPWR _0219_ _0221_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S4BEG0
+ _0226_ sg13g2_a21oi_1
X_0856_ _0288_ _0289_ _0290_ _0291_ VPWR VGND sg13g2_nor3_1
X_1408_ net751 net662 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
X_1339_ net777 net682 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_51_173 VPWR VGND sg13g2_fill_2
Xoutput390 net390 Tile_X0Y0_N2BEG[6] VPWR VGND sg13g2_buf_1
XFILLER_120_167 VPWR VGND sg13g2_decap_8
X_0641_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit26.Q net2
+ net6 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG15 net632 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit27.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG0 VPWR VGND sg13g2_mux4_1
X_1690_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG7 net544 VPWR
+ VGND sg13g2_buf_1
X_0710_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit14.Q net181
+ net189 net173 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG9
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit15.Q net292 VPWR
+ VGND sg13g2_mux4_1
XFILLER_51_70 VPWR VGND sg13g2_fill_2
X_0572_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG4 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG8
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit18.Q _0130_ VPWR
+ VGND sg13g2_mux2_1
X_1055_ net789 net675 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
X_1124_ net795 net657 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_102_101 VPWR VGND sg13g2_fill_2
X_0908_ net91 net732 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
X_0839_ _0275_ net151 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit2.Q
+ VPWR VGND sg13g2_nand2b_1
Xinput118 Tile_X0Y0_S2END[0] net118 VPWR VGND sg13g2_buf_1
Xinput129 Tile_X0Y0_S2MID[3] net129 VPWR VGND sg13g2_buf_1
Xinput107 Tile_X0Y0_FrameData[3] net107 VPWR VGND sg13g2_buf_1
XFILLER_16_118 VPWR VGND sg13g2_decap_4
XFILLER_108_0 VPWR VGND sg13g2_fill_2
XFILLER_21_95 VPWR VGND sg13g2_fill_1
X_1673_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S4BEG2 net518 VPWR
+ VGND sg13g2_buf_1
X_0624_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit25.Q net226
+ net3 _0074_ net28 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit24.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W1BEG3 VPWR VGND sg13g2_mux4_1
X_0555_ _0113_ _0115_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N4BEG1
+ VPWR VGND sg13g2_nor2_1
Xfanout808 net87 net808 VPWR VGND sg13g2_buf_1
X_0486_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit17.Q net16
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG10 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG6
+ net630 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit16.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG5
+ VPWR VGND sg13g2_mux4_1
XFILLER_23_0 VPWR VGND sg13g2_fill_1
X_1038_ net89 net687 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
X_1107_ net811 net663 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_88_187 VPWR VGND sg13g2_fill_2
X_0340_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit2.Q net53
+ net45 net64 net631 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit3.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG0 VPWR VGND sg13g2_mux4_1
X_1725_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG14 net570 VPWR
+ VGND sg13g2_buf_1
X_1587_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG4 net443 VPWR
+ VGND sg13g2_buf_1
X_0538_ _0101_ net42 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit7.Q
+ VPWR VGND sg13g2_nand2b_1
X_1656_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG1 net510 VPWR
+ VGND sg13g2_buf_1
Xfanout627 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG4 net627
+ VPWR VGND sg13g2_buf_1
Xfanout649 net650 net649 VPWR VGND sg13g2_buf_1
Xfanout638 _0079_ net638 VPWR VGND sg13g2_buf_1
X_0607_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit6.Q net226
+ net246 _0074_ net141 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit7.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG15 VPWR VGND sg13g2_mux4_1
X_0469_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit18.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END1
+ net248 net115 net135 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit19.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG5 VPWR VGND sg13g2_mux4_1
XFILLER_118_20 VPWR VGND sg13g2_decap_8
XFILLER_118_97 VPWR VGND sg13g2_decap_8
XFILLER_94_56 VPWR VGND sg13g2_fill_1
XFILLER_27_83 VPWR VGND sg13g2_fill_2
X_1510_ net701 net374 VPWR VGND sg13g2_buf_1
XFILLER_64_7 VPWR VGND sg13g2_fill_2
X_1441_ net752 net648 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
X_1372_ net778 net669 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
X_0323_ VPWR _0026_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit12.Q
+ VGND sg13g2_inv_1
XFILLER_90_0 VPWR VGND sg13g2_fill_2
X_1708_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG9 net564 VPWR
+ VGND sg13g2_buf_1
X_1639_ net761 net485 VPWR VGND sg13g2_buf_1
XFILLER_48_38 VPWR VGND sg13g2_fill_2
XFILLER_64_26 VPWR VGND sg13g2_fill_2
XFILLER_120_76 VPWR VGND sg13g2_decap_8
XFILLER_1_186 VPWR VGND sg13g2_decap_8
XFILLER_49_102 VPWR VGND sg13g2_fill_1
X_0941_ net805 net721 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_118_118 VPWR VGND sg13g2_decap_8
X_0872_ net799 net743 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
X_1355_ net760 net671 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
X_1424_ net765 net647 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_63_182 VPWR VGND sg13g2_decap_8
X_1286_ net759 net703 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
X_0306_ VPWR _0009_ net165 VGND sg13g2_inv_1
XFILLER_109_118 VPWR VGND sg13g2_fill_2
Xoutput572 net572 Tile_X0Y1_WW4BEG[1] VPWR VGND sg13g2_buf_1
Xoutput550 net550 Tile_X0Y1_W2BEGb[5] VPWR VGND sg13g2_buf_1
Xoutput561 net561 Tile_X0Y1_W6BEG[6] VPWR VGND sg13g2_buf_1
XFILLER_24_62 VPWR VGND sg13g2_fill_1
X_1140_ net812 net652 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
X_1071_ net807 net678 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_1_77 VPWR VGND sg13g2_decap_4
X_0924_ net104 net733 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
X_0786_ VGND VPWR _0028_ _0224_ _0226_ _0225_ sg13g2_a21oi_1
X_0855_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit4.Q VPWR
+ _0290_ VGND net129 _0283_ sg13g2_o21ai_1
XFILLER_53_0 VPWR VGND sg13g2_fill_2
XFILLER_114_198 VPWR VGND sg13g2_fill_2
X_1338_ net776 net682 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
X_1407_ net750 net660 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
X_1269_ net200 net706 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
Xoutput391 net391 Tile_X0Y0_N2BEG[7] VPWR VGND sg13g2_buf_1
XFILLER_120_146 VPWR VGND sg13g2_decap_8
Xoutput380 net380 Tile_X0Y0_N1BEG[0] VPWR VGND sg13g2_buf_1
XFILLER_74_200 VPWR VGND sg13g2_fill_1
XFILLER_42_152 VPWR VGND sg13g2_fill_2
X_0571_ _0127_ _0129_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N4BEG3
+ VPWR VGND sg13g2_nor2_1
X_0640_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit24.Q net31
+ net9 net640 net632 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit25.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb7 VPWR VGND sg13g2_mux4_1
XFILLER_111_113 VPWR VGND sg13g2_fill_2
X_1054_ net813 net690 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
X_1123_ net794 net657 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
X_0907_ net92 net733 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
Xinput108 Tile_X0Y0_FrameData[4] net108 VPWR VGND sg13g2_buf_1
X_0769_ net145 net183 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit11.Q
+ _0210_ VPWR VGND sg13g2_mux2_1
X_0838_ _0271_ _0272_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit0.Q
+ _0274_ VPWR VGND _0273_ sg13g2_nand4_1
Xinput119 Tile_X0Y0_S2END[1] net119 VPWR VGND sg13g2_buf_1
XFILLER_72_48 VPWR VGND sg13g2_decap_4
XFILLER_97_12 VPWR VGND sg13g2_fill_2
XFILLER_47_200 VPWR VGND sg13g2_fill_1
XFILLER_15_174 VPWR VGND sg13g2_fill_1
XFILLER_15_196 VPWR VGND sg13g2_fill_1
Xfanout809 net86 net809 VPWR VGND sg13g2_buf_1
X_0554_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit19.Q _0114_
+ _0115_ VPWR VGND sg13g2_nor2_1
X_1672_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S4BEG1 net532 VPWR
+ VGND sg13g2_buf_1
X_0623_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit23.Q net225
+ net2 _0067_ net29 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit22.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W1BEG2 VPWR VGND sg13g2_mux4_1
X_0485_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit15.Q net15
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG11 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG7
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit14.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG4 VPWR VGND sg13g2_mux4_1
X_1106_ net810 net665 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
X_1037_ net90 net688 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_21_100 VPWR VGND sg13g2_decap_8
Xinput90 Tile_X0Y0_FrameData[17] net90 VPWR VGND sg13g2_buf_1
XFILLER_29_200 VPWR VGND sg13g2_fill_1
XFILLER_83_58 VPWR VGND sg13g2_fill_1
XFILLER_16_96 VPWR VGND sg13g2_fill_1
XFILLER_79_199 VPWR VGND sg13g2_fill_2
XFILLER_92_4 VPWR VGND sg13g2_fill_2
X_1724_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG13 net569 VPWR
+ VGND sg13g2_buf_1
X_0537_ net50 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit6.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit7.Q _0100_ VPWR
+ VGND sg13g2_nor3_1
XFILLER_85_114 VPWR VGND sg13g2_decap_4
X_1586_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG3 net442 VPWR
+ VGND sg13g2_buf_1
Xfanout628 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG3 net628
+ VPWR VGND sg13g2_buf_1
X_1655_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG0 net509 VPWR
+ VGND sg13g2_buf_1
X_0606_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit4.Q net225
+ net245 _0067_ net140 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit5.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG14 VPWR VGND sg13g2_mux4_1
Xfanout639 _0078_ net639 VPWR VGND sg13g2_buf_1
X_0399_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit8.Q net50
+ net42 net56 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG3 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit9.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG3 VPWR VGND sg13g2_mux4_1
X_0468_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit24.Q net16
+ net20 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG6 net624 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit25.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG9 VPWR VGND sg13g2_mux4_1
XFILLER_118_76 VPWR VGND sg13g2_decap_8
X_1371_ net777 net671 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_4_55 VPWR VGND sg13g2_fill_1
X_1440_ net751 net650 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
X_0322_ VPWR _0025_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit11.Q
+ VGND sg13g2_inv_1
XFILLER_90_161 VPWR VGND sg13g2_fill_1
X_1638_ net209 net484 VPWR VGND sg13g2_buf_1
X_1707_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG8 net563 VPWR
+ VGND sg13g2_buf_1
X_1569_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG2 net423 VPWR
+ VGND sg13g2_buf_1
XFILLER_120_55 VPWR VGND sg13g2_decap_8
XFILLER_13_31 VPWR VGND sg13g2_fill_1
XFILLER_1_165 VPWR VGND sg13g2_decap_8
XFILLER_64_117 VPWR VGND sg13g2_fill_1
X_0940_ net804 net721 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
X_0871_ net798 net743 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
X_1285_ net756 net703 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
X_1354_ net758 net671 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
X_1423_ net764 net647 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
X_0305_ VPWR _0008_ net166 VGND sg13g2_inv_1
XFILLER_117_130 VPWR VGND sg13g2_decap_8
Xoutput573 net573 Tile_X0Y1_WW4BEG[2] VPWR VGND sg13g2_buf_1
Xoutput551 net551 Tile_X0Y1_W2BEGb[6] VPWR VGND sg13g2_buf_1
Xoutput540 net540 Tile_X0Y1_W2BEG[3] VPWR VGND sg13g2_buf_1
Xoutput562 net562 Tile_X0Y1_W6BEG[7] VPWR VGND sg13g2_buf_1
XFILLER_115_55 VPWR VGND sg13g2_decap_4
XFILLER_115_33 VPWR VGND sg13g2_fill_1
XFILLER_123_199 VPWR VGND sg13g2_fill_2
X_1070_ net89 net678 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_1_67 VPWR VGND sg13g2_decap_4
X_0923_ net107 net733 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
X_0854_ net150 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit5.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit6.Q _0289_ VPWR
+ VGND sg13g2_nor3_1
X_0785_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit8.Q VPWR
+ _0225_ VGND _0222_ _0223_ sg13g2_o21ai_1
X_1337_ net775 net682 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
X_1406_ net780 net660 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
X_1268_ net769 net706 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_28_106 VPWR VGND sg13g2_fill_2
X_1199_ net764 net727 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_51_175 VPWR VGND sg13g2_fill_1
Xoutput392 net392 Tile_X0Y0_N2BEGb[0] VPWR VGND sg13g2_buf_1
Xoutput370 net370 Tile_X0Y0_FrameStrobe_O[19] VPWR VGND sg13g2_buf_1
Xoutput381 net381 Tile_X0Y0_N1BEG[1] VPWR VGND sg13g2_buf_1
XFILLER_120_125 VPWR VGND sg13g2_decap_8
XFILLER_105_199 VPWR VGND sg13g2_fill_2
XFILLER_10_65 VPWR VGND sg13g2_fill_1
XFILLER_19_63 VPWR VGND sg13g2_fill_2
XFILLER_51_72 VPWR VGND sg13g2_fill_1
X_0570_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit25.Q _0128_
+ _0129_ VPWR VGND sg13g2_nor2_1
X_1122_ net793 net653 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
X_1053_ net802 net690 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_25_109 VPWR VGND sg13g2_decap_4
X_0906_ net94 net735 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
X_0837_ VGND VPWR _0273_ _0258_ net129 sg13g2_or2_1
Xinput109 Tile_X0Y0_FrameData[5] net109 VPWR VGND sg13g2_buf_1
X_0699_ VGND VPWR net150 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit26.Q
+ _0176_ _0175_ sg13g2_a21oi_1
X_0768_ _0208_ VPWR _0209_ VGND _0025_ _0158_ sg13g2_o21ai_1
XFILLER_112_89 VPWR VGND sg13g2_fill_2
XFILLER_108_2 VPWR VGND sg13g2_fill_1
X_1671_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S4BEG0 net531 VPWR
+ VGND sg13g2_buf_1
X_0553_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit18.Q net35
+ net65 net73 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG1 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit17.Q
+ _0114_ VPWR VGND sg13g2_mux4_1
XFILLER_97_112 VPWR VGND sg13g2_decap_4
X_0484_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit12.Q net250
+ net137 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG8 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG12
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit13.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG3
+ VPWR VGND sg13g2_mux4_1
X_0622_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit21.Q net224
+ net25 _0060_ net30 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit20.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W1BEG1 VPWR VGND sg13g2_mux4_1
X_1105_ net809 net665 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
X_1036_ net804 net687 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
Xinput91 Tile_X0Y0_FrameData[18] net91 VPWR VGND sg13g2_buf_1
Xinput80 Tile_X0Y0_EE4END[8] net80 VPWR VGND sg13g2_buf_1
XFILLER_88_189 VPWR VGND sg13g2_fill_1
XFILLER_88_167 VPWR VGND sg13g2_fill_2
XFILLER_16_42 VPWR VGND sg13g2_fill_2
XFILLER_32_41 VPWR VGND sg13g2_fill_2
XFILLER_57_82 VPWR VGND sg13g2_fill_1
X_1723_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG12 net568 VPWR
+ VGND sg13g2_buf_1
X_1654_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG7 net508 VPWR
+ VGND sg13g2_buf_1
X_1585_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG2 net441 VPWR
+ VGND sg13g2_buf_1
X_0467_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit20.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END2
+ net249 net116 net136 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit21.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG6 VPWR VGND sg13g2_mux4_1
Xfanout629 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG2 net629
+ VPWR VGND sg13g2_buf_1
X_0536_ VGND VPWR Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit4.Q
+ _0098_ _0099_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit5.Q
+ net259 _0041_ sg13g2_a221oi_1
X_0605_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit2.Q net224
+ net244 _0060_ net139 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit3.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG13 VPWR VGND sg13g2_mux4_1
X_0398_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit2.Q net51
+ net43 net61 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG2 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit3.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG2 VPWR VGND sg13g2_mux4_1
X_1019_ net788 net702 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_118_66 VPWR VGND sg13g2_fill_2
XFILLER_118_55 VPWR VGND sg13g2_decap_8
XFILLER_91_129 VPWR VGND sg13g2_fill_2
XFILLER_91_107 VPWR VGND sg13g2_fill_1
XFILLER_76_159 VPWR VGND sg13g2_fill_2
XFILLER_57_8 VPWR VGND sg13g2_decap_8
XFILLER_4_185 VPWR VGND sg13g2_decap_4
XFILLER_4_34 VPWR VGND sg13g2_decap_8
X_1370_ net776 net670 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
X_0321_ VPWR _0024_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit9.Q
+ VGND sg13g2_inv_1
XFILLER_75_181 VPWR VGND sg13g2_fill_1
XFILLER_90_2 VPWR VGND sg13g2_fill_1
X_1706_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG7 net562 VPWR
+ VGND sg13g2_buf_1
X_1637_ net208 net483 VPWR VGND sg13g2_buf_1
X_0519_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit18.Q net74
+ net67 net55 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG10 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit19.Q
+ net280 VPWR VGND sg13g2_mux4_1
X_1499_ net99 net345 VPWR VGND sg13g2_buf_1
X_1568_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG1 net422 VPWR
+ VGND sg13g2_buf_1
XFILLER_120_34 VPWR VGND sg13g2_decap_8
XFILLER_64_28 VPWR VGND sg13g2_fill_1
X_0870_ net797 net748 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_54_83 VPWR VGND sg13g2_decap_4
X_1422_ net208 net649 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
X_0304_ VPWR _0007_ net167 VGND sg13g2_inv_1
X_1353_ net757 net672 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
X_1284_ net755 net706 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_55_129 VPWR VGND sg13g2_decap_4
X_0999_ net798 net700 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
Xoutput552 net552 Tile_X0Y1_W2BEGb[7] VPWR VGND sg13g2_buf_1
Xoutput574 net574 Tile_X0Y1_WW4BEG[3] VPWR VGND sg13g2_buf_1
Xoutput541 net541 Tile_X0Y1_W2BEG[4] VPWR VGND sg13g2_buf_1
Xoutput530 net530 Tile_X0Y1_S4BEG[7] VPWR VGND sg13g2_buf_1
Xoutput563 net563 Tile_X0Y1_W6BEG[8] VPWR VGND sg13g2_buf_1
XFILLER_115_78 VPWR VGND sg13g2_decap_4
XFILLER_54_195 VPWR VGND sg13g2_fill_2
XFILLER_123_145 VPWR VGND sg13g2_decap_4
Xfanout790 net105 net790 VPWR VGND sg13g2_buf_1
XFILLER_1_13 VPWR VGND sg13g2_fill_1
XFILLER_45_140 VPWR VGND sg13g2_fill_2
X_0922_ net787 net731 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
X_0853_ _0037_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit6.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG0 _0288_ VPWR VGND sg13g2_nor3_1
X_1405_ net779 net660 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
X_0784_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG4 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG8
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit6.Q _0224_ VPWR
+ VGND sg13g2_mux2_1
XFILLER_39_0 VPWR VGND sg13g2_fill_2
Xinput1 CONFIGURED_top net1 VPWR VGND sg13g2_buf_1
X_1198_ net763 net725 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
X_1336_ net774 net681 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
X_1267_ net768 net706 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_10_55 VPWR VGND sg13g2_fill_2
Xoutput371 net371 Tile_X0Y0_FrameStrobe_O[1] VPWR VGND sg13g2_buf_1
Xoutput360 net360 Tile_X0Y0_FrameStrobe_O[0] VPWR VGND sg13g2_buf_1
Xoutput393 net393 Tile_X0Y0_N2BEGb[1] VPWR VGND sg13g2_buf_1
Xoutput382 net382 Tile_X0Y0_N1BEG[2] VPWR VGND sg13g2_buf_1
XFILLER_120_104 VPWR VGND sg13g2_decap_8
XFILLER_105_167 VPWR VGND sg13g2_fill_2
XFILLER_42_154 VPWR VGND sg13g2_fill_1
XFILLER_111_115 VPWR VGND sg13g2_fill_1
X_1121_ net792 net653 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
X_1052_ net791 net690 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
X_0905_ net95 net734 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
X_0767_ VPWR _0208_ _0207_ VGND sg13g2_inv_1
X_0836_ net150 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit1.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit2.Q _0272_ VPWR
+ VGND sg13g2_or3_1
X_0698_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit26.Q net158
+ _0175_ VPWR VGND sg13g2_nor2b_1
X_1319_ net201 net696 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_21_21 VPWR VGND sg13g2_fill_1
XFILLER_97_14 VPWR VGND sg13g2_fill_1
XFILLER_15_121 VPWR VGND sg13g2_fill_1
XFILLER_30_124 VPWR VGND sg13g2_fill_2
X_1670_ Tile_X0Y0_S4END[15] net530 VPWR VGND sg13g2_buf_1
X_0621_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit19.Q net223
+ net14 _0088_ net31 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit18.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W1BEG0 VPWR VGND sg13g2_mux4_1
X_0483_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit10.Q net249
+ net136 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG9 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG13
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit11.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG2
+ VPWR VGND sg13g2_mux4_1
X_0552_ VGND VPWR _0012_ _0109_ _0113_ _0112_ sg13g2_a21oi_1
X_1104_ net808 net664 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
X_1035_ net803 net687 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
Xinput92 Tile_X0Y0_FrameData[19] net92 VPWR VGND sg13g2_buf_1
Xinput81 Tile_X0Y0_EE4END[9] net81 VPWR VGND sg13g2_buf_1
Xinput70 Tile_X0Y0_EE4END[13] net70 VPWR VGND sg13g2_buf_1
XFILLER_88_113 VPWR VGND sg13g2_fill_1
X_0819_ VGND VPWR _0034_ _0254_ _0256_ _0255_ sg13g2_a21oi_1
XFILLER_12_146 VPWR VGND sg13g2_fill_1
XFILLER_106_0 VPWR VGND sg13g2_fill_2
XFILLER_92_6 VPWR VGND sg13g2_fill_1
X_1584_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG1 net440 VPWR
+ VGND sg13g2_buf_1
XFILLER_7_194 VPWR VGND sg13g2_fill_2
X_1722_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG11 net567 VPWR
+ VGND sg13g2_buf_1
X_0604_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit0.Q net223
+ net243 _0088_ net138 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit1.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG12 VPWR VGND sg13g2_mux4_1
X_1653_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG6 net507 VPWR
+ VGND sg13g2_buf_1
X_0466_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit22.Q net15
+ net19 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG7 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG7
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit23.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG8
+ VPWR VGND sg13g2_mux4_1
X_0535_ _0099_ net41 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit5.Q
+ VPWR VGND sg13g2_nand2b_1
X_0397_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit12.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb2
+ net237 net128 net120 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit13.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG2 VPWR VGND sg13g2_mux4_1
X_1018_ net787 net697 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_118_34 VPWR VGND sg13g2_decap_8
XFILLER_4_164 VPWR VGND sg13g2_decap_8
X_0320_ VPWR _0023_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit8.Q
+ VGND sg13g2_inv_1
X_1705_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG6 net561 VPWR
+ VGND sg13g2_buf_1
X_0518_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit16.Q net73
+ net81 net65 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG9 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit17.Q
+ net279 VPWR VGND sg13g2_mux4_1
X_1567_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG0 net421 VPWR
+ VGND sg13g2_buf_1
X_1636_ net764 net482 VPWR VGND sg13g2_buf_1
X_1498_ net98 net344 VPWR VGND sg13g2_buf_1
X_0449_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit0.Q net16
+ net24 net629 net625 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit1.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb5 VPWR VGND sg13g2_mux4_1
XFILLER_81_196 VPWR VGND sg13g2_fill_1
XFILLER_1_112 VPWR VGND sg13g2_decap_8
XFILLER_64_108 VPWR VGND sg13g2_fill_1
XFILLER_57_171 VPWR VGND sg13g2_fill_2
XFILLER_62_7 VPWR VGND sg13g2_decap_8
X_1421_ net209 net649 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
X_0303_ VPWR _0006_ net54 VGND sg13g2_inv_1
X_1352_ net781 net691 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
X_1283_ net754 net706 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_117_176 VPWR VGND sg13g2_decap_8
XFILLER_117_154 VPWR VGND sg13g2_decap_8
X_0998_ net797 net701 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
Xoutput520 net520 Tile_X0Y1_S4BEG[12] VPWR VGND sg13g2_buf_1
XFILLER_117_187 VPWR VGND sg13g2_fill_2
XFILLER_86_200 VPWR VGND sg13g2_fill_1
XFILLER_59_29 VPWR VGND sg13g2_fill_1
XFILLER_59_18 VPWR VGND sg13g2_decap_8
Xoutput553 net553 Tile_X0Y1_W6BEG[0] VPWR VGND sg13g2_buf_1
X_1619_ net751 net495 VPWR VGND sg13g2_buf_1
Xoutput575 net575 Tile_X0Y1_WW4BEG[4] VPWR VGND sg13g2_buf_1
Xoutput542 net542 Tile_X0Y1_W2BEG[5] VPWR VGND sg13g2_buf_1
Xoutput531 net531 Tile_X0Y1_S4BEG[8] VPWR VGND sg13g2_buf_1
Xoutput564 net564 Tile_X0Y1_W6BEG[9] VPWR VGND sg13g2_buf_1
XFILLER_39_182 VPWR VGND sg13g2_fill_1
XFILLER_24_21 VPWR VGND sg13g2_fill_2
Xfanout791 net104 net791 VPWR VGND sg13g2_buf_1
XFILLER_37_119 VPWR VGND sg13g2_decap_4
Xfanout780 net191 net780 VPWR VGND sg13g2_buf_1
X_0921_ net786 net731 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_81_93 VPWR VGND sg13g2_fill_2
X_0783_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit7.Q VPWR
+ _0223_ VGND Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit6.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG12 sg13g2_o21ai_1
X_0852_ _0286_ VPWR _0287_ VGND _0037_ _0279_ sg13g2_o21ai_1
XFILLER_68_200 VPWR VGND sg13g2_fill_1
X_1335_ net773 net681 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
X_1404_ net193 net662 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
Xinput2 DOUT_SRAM0 net2 VPWR VGND sg13g2_buf_1
X_1266_ net767 net703 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
X_1197_ net762 net726 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_28_108 VPWR VGND sg13g2_fill_1
XFILLER_36_130 VPWR VGND sg13g2_decap_4
XFILLER_36_196 VPWR VGND sg13g2_fill_1
Xoutput361 net361 Tile_X0Y0_FrameStrobe_O[10] VPWR VGND sg13g2_buf_1
Xoutput350 net350 Tile_X0Y0_FrameData_O[2] VPWR VGND sg13g2_buf_1
Xoutput372 net372 Tile_X0Y0_FrameStrobe_O[2] VPWR VGND sg13g2_buf_1
Xoutput394 net394 Tile_X0Y0_N2BEGb[2] VPWR VGND sg13g2_buf_1
Xoutput383 net383 Tile_X0Y0_N1BEG[3] VPWR VGND sg13g2_buf_1
XFILLER_113_190 VPWR VGND sg13g2_fill_2
XFILLER_35_20 VPWR VGND sg13g2_fill_2
XFILLER_42_199 VPWR VGND sg13g2_fill_2
X_1120_ net105 net655 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
X_1051_ net788 net690 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_18_141 VPWR VGND sg13g2_fill_2
X_0904_ net96 net734 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_33_199 VPWR VGND sg13g2_fill_2
X_0697_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit27.Q net635
+ _0174_ VPWR VGND Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit26.Q
+ sg13g2_nand3b_1
X_0766_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit12.Q VPWR
+ _0207_ VGND net164 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit11.Q
+ sg13g2_o21ai_1
X_0835_ _0271_ _0257_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG0
+ VPWR VGND sg13g2_nand2b_1
X_1318_ net759 net692 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
X_1249_ net752 net716 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_24_155 VPWR VGND sg13g2_fill_1
XFILLER_21_55 VPWR VGND sg13g2_fill_2
X_0551_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit19.Q VPWR
+ _0112_ VGND _0110_ _0111_ sg13g2_o21ai_1
X_0620_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit5.Q net145
+ net146 net154 net632 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit4.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG7 VPWR VGND sg13g2_mux4_1
X_0482_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit8.Q net248
+ net135 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG10 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG14
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit9.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG1
+ VPWR VGND sg13g2_mux4_1
X_1103_ net807 net664 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
X_1034_ net801 net686 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_99_0 VPWR VGND sg13g2_fill_2
Xinput93 Tile_X0Y0_FrameData[1] net93 VPWR VGND sg13g2_buf_1
Xinput82 Tile_X0Y0_FrameData[0] net82 VPWR VGND sg13g2_buf_1
Xinput60 Tile_X0Y0_E6END[4] net60 VPWR VGND sg13g2_buf_1
Xinput71 Tile_X0Y0_EE4END[14] net71 VPWR VGND sg13g2_buf_1
XFILLER_107_58 VPWR VGND sg13g2_fill_2
X_0749_ _0021_ net639 _0192_ VPWR VGND sg13g2_nor2_1
X_0818_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit17.Q VPWR
+ _0255_ VGND _0252_ _0253_ sg13g2_o21ai_1
XFILLER_88_169 VPWR VGND sg13g2_fill_1
X_1721_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG10 net566 VPWR
+ VGND sg13g2_buf_1
X_0603_ _0155_ _0157_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S4BEG3
+ VPWR VGND sg13g2_nor2_1
X_1583_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG0 net437 VPWR
+ VGND sg13g2_buf_1
X_0534_ net49 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit4.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit5.Q _0098_ VPWR
+ VGND sg13g2_nor3_1
X_1652_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG5 net506 VPWR
+ VGND sg13g2_buf_1
X_0465_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit22.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END3
+ net250 net117 net137 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit23.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG7 VPWR VGND sg13g2_mux4_1
XFILLER_78_180 VPWR VGND sg13g2_fill_1
X_0396_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit23.Q net159
+ net169 net151 _0079_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit22.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb2 VPWR VGND sg13g2_mux4_1
X_1017_ net786 net697 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_68_83 VPWR VGND sg13g2_fill_1
Xinput250 Tile_X0Y1_N4END[7] net250 VPWR VGND sg13g2_buf_1
X_1704_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG5 net560 VPWR
+ VGND sg13g2_buf_1
X_1497_ net97 net343 VPWR VGND sg13g2_buf_1
X_1566_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W1BEG3 net420 VPWR
+ VGND sg13g2_buf_1
X_0517_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit14.Q net66
+ net80 net64 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG8 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit15.Q
+ net278 VPWR VGND sg13g2_mux4_1
X_1635_ net765 net481 VPWR VGND sg13g2_buf_1
X_0379_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit30.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit31.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END3 _0072_ VPWR VGND sg13g2_nor3_1
X_0448_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit30.Q net15
+ net23 net628 net626 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit31.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb4 VPWR VGND sg13g2_mux4_1
XFILLER_66_194 VPWR VGND sg13g2_fill_2
XFILLER_120_69 VPWR VGND sg13g2_decap_8
XFILLER_1_179 VPWR VGND sg13g2_decap_8
XFILLER_70_51 VPWR VGND sg13g2_fill_1
X_0302_ VPWR _0005_ net59 VGND sg13g2_inv_1
X_1351_ net770 net691 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
X_1420_ net210 net649 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
X_1282_ net753 net703 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_48_161 VPWR VGND sg13g2_fill_1
XFILLER_63_175 VPWR VGND sg13g2_decap_8
X_0997_ net796 net700 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
Xoutput543 net543 Tile_X0Y1_W2BEG[6] VPWR VGND sg13g2_buf_1
Xoutput510 net510 Tile_X0Y1_S2BEGb[1] VPWR VGND sg13g2_buf_1
Xoutput532 net532 Tile_X0Y1_S4BEG[9] VPWR VGND sg13g2_buf_1
Xoutput521 net521 Tile_X0Y1_S4BEG[13] VPWR VGND sg13g2_buf_1
Xoutput554 net554 Tile_X0Y1_W6BEG[10] VPWR VGND sg13g2_buf_1
X_1618_ net219 net494 VPWR VGND sg13g2_buf_1
X_1549_ Tile_X0Y1_N4END[11] net409 VPWR VGND sg13g2_buf_1
Xoutput576 net576 Tile_X0Y1_WW4BEG[5] VPWR VGND sg13g2_buf_1
Xoutput565 net565 Tile_X0Y1_WW4BEG[0] VPWR VGND sg13g2_buf_1
XFILLER_40_87 VPWR VGND sg13g2_fill_1
Xfanout792 net103 net792 VPWR VGND sg13g2_buf_1
Xfanout770 net201 net770 VPWR VGND sg13g2_buf_1
Xfanout781 net190 net781 VPWR VGND sg13g2_buf_1
X_0920_ net110 net732 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
X_0782_ _0027_ net636 _0222_ VPWR VGND sg13g2_nor2_1
X_0851_ _0286_ _0284_ _0285_ _0282_ _0280_ VPWR VGND sg13g2_a22oi_1
X_1265_ net766 net703 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
X_1334_ net772 net684 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
X_1403_ net194 net668 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
X_1196_ net761 net725 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
Xinput3 DOUT_SRAM1 net3 VPWR VGND sg13g2_buf_1
Xoutput373 net373 Tile_X0Y0_FrameStrobe_O[3] VPWR VGND sg13g2_buf_1
Xoutput384 net384 Tile_X0Y0_N2BEG[0] VPWR VGND sg13g2_buf_1
Xoutput362 net362 Tile_X0Y0_FrameStrobe_O[11] VPWR VGND sg13g2_buf_1
Xoutput395 net395 Tile_X0Y0_N2BEGb[3] VPWR VGND sg13g2_buf_1
XFILLER_105_169 VPWR VGND sg13g2_fill_1
XFILLER_105_125 VPWR VGND sg13g2_fill_2
XFILLER_105_103 VPWR VGND sg13g2_fill_1
Xoutput351 net351 Tile_X0Y0_FrameData_O[30] VPWR VGND sg13g2_buf_1
Xoutput340 net340 Tile_X0Y0_FrameData_O[20] VPWR VGND sg13g2_buf_1
XFILLER_120_139 VPWR VGND sg13g2_decap_8
XFILLER_19_22 VPWR VGND sg13g2_fill_2
XFILLER_42_112 VPWR VGND sg13g2_decap_4
X_1050_ net787 net686 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
X_0903_ net97 net734 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
X_0834_ _0266_ _0269_ _0264_ _0270_ VPWR VGND sg13g2_nand3_1
X_0765_ VGND VPWR _0199_ _0201_ Tile_X0Y0_IHP_SRAM_top.N4BEG_outbuf_10.A _0206_ sg13g2_a21oi_1
X_0696_ _0171_ VPWR net254 VGND Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit25.Q
+ _0173_ sg13g2_o21ai_1
XFILLER_102_128 VPWR VGND sg13g2_fill_2
X_1317_ net756 net692 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_2_91 VPWR VGND sg13g2_decap_8
X_1248_ net751 net715 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
X_1179_ net777 net740 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_62_85 VPWR VGND sg13g2_fill_1
X_0550_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit18.Q VPWR
+ _0111_ VGND Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit17.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG13 sg13g2_o21ai_1
X_1102_ net806 net664 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
X_0481_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit6.Q net247
+ net134 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG11 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG15
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit7.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG0
+ VPWR VGND sg13g2_mux4_1
X_1033_ net800 net686 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
Xinput61 Tile_X0Y0_E6END[5] net61 VPWR VGND sg13g2_buf_1
Xinput72 Tile_X0Y0_EE4END[15] net72 VPWR VGND sg13g2_buf_1
Xinput50 Tile_X0Y0_E2MID[4] net50 VPWR VGND sg13g2_buf_1
X_0817_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG7 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG11
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit15.Q _0254_ VPWR
+ VGND sg13g2_mux2_1
Xinput94 Tile_X0Y0_FrameData[20] net94 VPWR VGND sg13g2_buf_1
Xinput83 Tile_X0Y0_FrameData[10] net83 VPWR VGND sg13g2_buf_1
X_0679_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit15.Q net14
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG5 _0160_ net633
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit14.Q Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG10
+ VPWR VGND sg13g2_mux4_1
X_0748_ VGND VPWR _0022_ _0190_ _0191_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit7.Q
+ sg13g2_a21oi_1
XFILLER_16_12 VPWR VGND sg13g2_fill_1
XFILLER_106_2 VPWR VGND sg13g2_fill_1
XFILLER_79_148 VPWR VGND sg13g2_fill_1
XFILLER_73_62 VPWR VGND sg13g2_decap_4
X_1720_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG9 net580 VPWR
+ VGND sg13g2_buf_1
X_1651_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG4 net505 VPWR
+ VGND sg13g2_buf_1
X_0533_ VGND VPWR Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit2.Q
+ _0096_ _0097_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit3.Q
+ net258 _0040_ sg13g2_a221oi_1
X_0602_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit29.Q _0156_
+ _0157_ VPWR VGND sg13g2_nor2_1
XFILLER_85_107 VPWR VGND sg13g2_decap_8
X_1582_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb7 net436 VPWR
+ VGND sg13g2_buf_1
X_0464_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit20.Q net18
+ net22 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG8 net631 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit21.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG7 VPWR VGND sg13g2_mux4_1
XFILLER_7_196 VPWR VGND sg13g2_fill_1
XFILLER_85_118 VPWR VGND sg13g2_fill_1
X_0395_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit13.Q net237
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG2 net229 net128 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit12.Q
+ _0079_ VPWR VGND sg13g2_mux4_1
X_1016_ net785 net697 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_43_10 VPWR VGND sg13g2_fill_1
XFILLER_4_48 VPWR VGND sg13g2_decap_8
Xinput240 Tile_X0Y1_N2MID[5] net240 VPWR VGND sg13g2_buf_1
X_1703_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG4 net559 VPWR
+ VGND sg13g2_buf_1
X_1634_ net205 net480 VPWR VGND sg13g2_buf_1
X_1496_ net96 net342 VPWR VGND sg13g2_buf_1
X_0516_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit12.Q net79
+ net72 net63 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG7 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit13.Q
+ net277 VPWR VGND sg13g2_mux4_1
X_1565_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W1BEG2 net419 VPWR
+ VGND sg13g2_buf_1
X_0447_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit28.Q net13
+ net22 net628 net626 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit29.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb3 VPWR VGND sg13g2_mux4_1
XFILLER_58_129 VPWR VGND sg13g2_decap_4
XFILLER_120_48 VPWR VGND sg13g2_decap_8
X_0378_ _0071_ net117 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit30.Q
+ VPWR VGND sg13g2_nand2b_1
XFILLER_13_57 VPWR VGND sg13g2_fill_2
XFILLER_1_158 VPWR VGND sg13g2_decap_8
XFILLER_57_195 VPWR VGND sg13g2_fill_2
XFILLER_57_173 VPWR VGND sg13g2_fill_1
XFILLER_55_8 VPWR VGND sg13g2_fill_1
X_0301_ VPWR _0004_ net58 VGND sg13g2_inv_1
X_1350_ net759 net680 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_0_180 VPWR VGND sg13g2_decap_8
X_1281_ net752 net703 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
X_0996_ net795 net698 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_74_0 VPWR VGND sg13g2_fill_2
XFILLER_117_123 VPWR VGND sg13g2_decap_8
Xoutput577 net577 Tile_X0Y1_WW4BEG[6] VPWR VGND sg13g2_buf_1
Xoutput544 net544 Tile_X0Y1_W2BEG[7] VPWR VGND sg13g2_buf_1
Xoutput533 net533 Tile_X0Y1_W1BEG[0] VPWR VGND sg13g2_buf_1
Xoutput500 net500 Tile_X0Y1_S1BEG[3] VPWR VGND sg13g2_buf_1
Xoutput511 net511 Tile_X0Y1_S2BEGb[2] VPWR VGND sg13g2_buf_1
Xoutput522 net522 Tile_X0Y1_S4BEG[14] VPWR VGND sg13g2_buf_1
Xoutput566 net566 Tile_X0Y1_WW4BEG[10] VPWR VGND sg13g2_buf_1
Xoutput555 net555 Tile_X0Y1_W6BEG[11] VPWR VGND sg13g2_buf_1
X_1617_ net218 net493 VPWR VGND sg13g2_buf_1
X_1548_ Tile_X0Y1_N4END[10] net408 VPWR VGND sg13g2_buf_1
XFILLER_115_59 VPWR VGND sg13g2_fill_2
X_1479_ net786 net355 VPWR VGND sg13g2_buf_1
XFILLER_91_29 VPWR VGND sg13g2_fill_2
XFILLER_24_23 VPWR VGND sg13g2_fill_1
Xfanout760 net211 net760 VPWR VGND sg13g2_buf_1
Xfanout793 net102 net793 VPWR VGND sg13g2_buf_1
XFILLER_105_81 VPWR VGND sg13g2_fill_1
Xfanout782 net113 net782 VPWR VGND sg13g2_buf_1
Xfanout771 net200 net771 VPWR VGND sg13g2_buf_1
XFILLER_121_80 VPWR VGND sg13g2_decap_8
X_0850_ VGND VPWR net160 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit4.Q
+ _0285_ _0283_ sg13g2_a21oi_1
X_0781_ VGND VPWR _0028_ _0220_ _0221_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit8.Q
+ sg13g2_a21oi_1
X_1402_ net195 net662 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
Xinput4 DOUT_SRAM10 net4 VPWR VGND sg13g2_buf_1
X_1333_ net771 net684 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_36_110 VPWR VGND sg13g2_fill_2
X_1264_ net765 net707 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_101_17 VPWR VGND sg13g2_fill_2
X_1195_ net760 net725 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_51_113 VPWR VGND sg13g2_decap_4
X_0979_ net84 net712 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
Xoutput363 net363 Tile_X0Y0_FrameStrobe_O[12] VPWR VGND sg13g2_buf_1
Xoutput374 net374 Tile_X0Y0_FrameStrobe_O[4] VPWR VGND sg13g2_buf_1
Xoutput396 net396 Tile_X0Y0_N2BEGb[4] VPWR VGND sg13g2_buf_1
Xoutput385 net385 Tile_X0Y0_N2BEG[1] VPWR VGND sg13g2_buf_1
XFILLER_120_118 VPWR VGND sg13g2_decap_8
XFILLER_113_192 VPWR VGND sg13g2_fill_1
Xoutput352 net352 Tile_X0Y0_FrameData_O[31] VPWR VGND sg13g2_buf_1
Xoutput341 net341 Tile_X0Y0_FrameData_O[21] VPWR VGND sg13g2_buf_1
Xoutput330 net330 Tile_X0Y0_FrameData_O[11] VPWR VGND sg13g2_buf_1
XFILLER_27_143 VPWR VGND sg13g2_fill_1
XFILLER_18_143 VPWR VGND sg13g2_fill_1
XFILLER_33_168 VPWR VGND sg13g2_fill_2
X_0902_ net797 net731 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
X_0833_ _0269_ _0268_ _0257_ _0261_ _0259_ VPWR VGND sg13g2_a22oi_1
XFILLER_37_0 VPWR VGND sg13g2_fill_2
X_0764_ VGND VPWR _0024_ _0204_ _0206_ _0205_ sg13g2_a21oi_1
X_0695_ VGND VPWR net149 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit24.Q
+ _0173_ _0172_ sg13g2_a21oi_1
X_1316_ net755 net692 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_2_70 VPWR VGND sg13g2_decap_8
X_1247_ net750 net714 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
X_1178_ net776 net741 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_101_140 VPWR VGND sg13g2_fill_1
XFILLER_15_146 VPWR VGND sg13g2_fill_2
XFILLER_46_98 VPWR VGND sg13g2_fill_2
XFILLER_62_31 VPWR VGND sg13g2_decap_4
XFILLER_7_59 VPWR VGND sg13g2_fill_1
XFILLER_97_116 VPWR VGND sg13g2_fill_2
XFILLER_97_105 VPWR VGND sg13g2_decap_8
X_0480_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit4.Q net13
+ net27 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG0 net631 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit5.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG15 VPWR VGND sg13g2_mux4_1
XFILLER_11_90 VPWR VGND sg13g2_decap_8
X_1101_ net805 net664 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
X_1032_ net799 net686 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
Xinput95 Tile_X0Y0_FrameData[21] net95 VPWR VGND sg13g2_buf_1
Xinput84 Tile_X0Y0_FrameData[11] net84 VPWR VGND sg13g2_buf_1
Xinput62 Tile_X0Y0_E6END[6] net62 VPWR VGND sg13g2_buf_1
Xinput73 Tile_X0Y0_EE4END[1] net73 VPWR VGND sg13g2_buf_1
Xinput51 Tile_X0Y0_E2MID[5] net51 VPWR VGND sg13g2_buf_1
Xinput40 Tile_X0Y0_E2END[2] net40 VPWR VGND sg13g2_buf_1
X_0747_ net143 net181 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit5.Q
+ _0190_ VPWR VGND sg13g2_mux2_1
X_0816_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit16.Q VPWR
+ _0253_ VGND Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit15.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG15 sg13g2_o21ai_1
X_0678_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit13.Q net3
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG6 _0159_ net634
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit12.Q Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG9
+ VPWR VGND sg13g2_mux4_1
XFILLER_12_127 VPWR VGND sg13g2_fill_2
XFILLER_94_119 VPWR VGND sg13g2_fill_2
XFILLER_57_64 VPWR VGND sg13g2_fill_1
X_0601_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit28.Q net37
+ net63 net72 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG3 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit27.Q
+ _0156_ VPWR VGND sg13g2_mux4_1
X_1581_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb6 net435 VPWR
+ VGND sg13g2_buf_1
X_1650_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG3 net504 VPWR
+ VGND sg13g2_buf_1
X_0532_ _0097_ net40 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit3.Q
+ VPWR VGND sg13g2_nand2b_1
XFILLER_98_93 VPWR VGND sg13g2_fill_1
X_0394_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit6.Q net51
+ net43 net55 net629 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit7.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG2 VPWR VGND sg13g2_mux4_1
X_0463_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit24.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END0
+ net247 net114 net134 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit25.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG8 VPWR VGND sg13g2_mux4_1
XFILLER_93_163 VPWR VGND sg13g2_fill_2
X_1015_ net784 net700 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_118_48 VPWR VGND sg13g2_decap_8
XFILLER_4_178 VPWR VGND sg13g2_decap_8
XFILLER_4_27 VPWR VGND sg13g2_decap_8
Xinput241 Tile_X0Y1_N2MID[6] net241 VPWR VGND sg13g2_buf_1
Xinput230 Tile_X0Y1_N2END[3] net230 VPWR VGND sg13g2_buf_1
X_1564_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W1BEG1 net418 VPWR
+ VGND sg13g2_buf_1
X_1702_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG3 net558 VPWR
+ VGND sg13g2_buf_1
X_1633_ net204 net479 VPWR VGND sg13g2_buf_1
X_0515_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit10.Q net78
+ net71 net62 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG6 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit11.Q
+ net276 VPWR VGND sg13g2_mux4_1
X_1495_ net800 net341 VPWR VGND sg13g2_buf_1
X_0377_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit26.Q net36
+ net62 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG14 _0066_
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit27.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1BEG2
+ VPWR VGND sg13g2_mux4_1
X_0446_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit26.Q net12
+ net21 net629 net625 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit27.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb2 VPWR VGND sg13g2_mux4_1
XFILLER_120_27 VPWR VGND sg13g2_decap_8
XFILLER_66_196 VPWR VGND sg13g2_fill_1
XFILLER_89_200 VPWR VGND sg13g2_fill_1
XFILLER_54_87 VPWR VGND sg13g2_fill_1
XFILLER_119_80 VPWR VGND sg13g2_decap_8
X_0300_ VPWR _0003_ net57 VGND sg13g2_inv_1
X_1280_ net751 net707 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_117_102 VPWR VGND sg13g2_decap_4
X_0995_ net794 net698 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
Xoutput556 net556 Tile_X0Y1_W6BEG[1] VPWR VGND sg13g2_buf_1
Xoutput545 net545 Tile_X0Y1_W2BEGb[0] VPWR VGND sg13g2_buf_1
Xoutput578 net578 Tile_X0Y1_WW4BEG[7] VPWR VGND sg13g2_buf_1
X_1547_ Tile_X0Y1_N4END[9] net407 VPWR VGND sg13g2_buf_1
Xoutput534 net534 Tile_X0Y1_W1BEG[1] VPWR VGND sg13g2_buf_1
Xoutput501 net501 Tile_X0Y1_S2BEG[0] VPWR VGND sg13g2_buf_1
Xoutput512 net512 Tile_X0Y1_S2BEGb[3] VPWR VGND sg13g2_buf_1
Xoutput523 net523 Tile_X0Y1_S4BEG[15] VPWR VGND sg13g2_buf_1
Xoutput567 net567 Tile_X0Y1_WW4BEG[11] VPWR VGND sg13g2_buf_1
X_1616_ net217 net492 VPWR VGND sg13g2_buf_1
X_1478_ net787 net354 VPWR VGND sg13g2_buf_1
X_0429_ _0090_ _0088_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit24.Q
+ VPWR VGND sg13g2_nand2b_1
XFILLER_123_149 VPWR VGND sg13g2_fill_2
Xfanout794 net101 net794 VPWR VGND sg13g2_buf_1
Xfanout783 net112 net783 VPWR VGND sg13g2_buf_1
Xfanout750 net221 net750 VPWR VGND sg13g2_buf_1
Xfanout761 net210 net761 VPWR VGND sg13g2_buf_1
XFILLER_49_98 VPWR VGND sg13g2_decap_4
Xfanout772 net199 net772 VPWR VGND sg13g2_buf_1
XFILLER_65_75 VPWR VGND sg13g2_decap_4
X_0780_ net142 net177 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit6.Q
+ _0220_ VPWR VGND sg13g2_mux2_1
XFILLER_114_116 VPWR VGND sg13g2_fill_2
X_1401_ net196 net662 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
X_1332_ net769 net681 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
Xinput5 DOUT_SRAM11 net5 VPWR VGND sg13g2_buf_1
XFILLER_36_144 VPWR VGND sg13g2_fill_2
X_1263_ net764 net707 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
X_1194_ net213 net728 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
X_0978_ net85 net710 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
Xoutput375 net375 Tile_X0Y0_FrameStrobe_O[5] VPWR VGND sg13g2_buf_1
Xoutput386 net386 Tile_X0Y0_N2BEG[2] VPWR VGND sg13g2_buf_1
Xoutput364 net364 Tile_X0Y0_FrameStrobe_O[13] VPWR VGND sg13g2_buf_1
Xoutput397 net397 Tile_X0Y0_N2BEGb[5] VPWR VGND sg13g2_buf_1
XFILLER_105_127 VPWR VGND sg13g2_fill_1
Xoutput342 net342 Tile_X0Y0_FrameData_O[22] VPWR VGND sg13g2_buf_1
Xoutput331 net331 Tile_X0Y0_FrameData_O[12] VPWR VGND sg13g2_buf_1
Xoutput353 net353 Tile_X0Y0_FrameData_O[3] VPWR VGND sg13g2_buf_1
Xoutput320 net320 DIN_SRAM4 VPWR VGND sg13g2_buf_1
XFILLER_19_24 VPWR VGND sg13g2_fill_1
XFILLER_116_81 VPWR VGND sg13g2_decap_8
XFILLER_76_96 VPWR VGND sg13g2_fill_2
XFILLER_18_199 VPWR VGND sg13g2_fill_2
X_0901_ net796 net731 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
X_0763_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit10.Q VPWR
+ _0205_ VGND _0202_ _0203_ sg13g2_o21ai_1
X_0832_ VGND VPWR net230 _0035_ _0268_ _0267_ sg13g2_a21oi_1
XFILLER_110_141 VPWR VGND sg13g2_fill_2
X_1315_ net754 net692 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
X_0694_ _0000_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit24.Q
+ _0172_ VPWR VGND sg13g2_nor2_1
X_1246_ net780 net717 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
X_1177_ net775 net740 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_62_21 VPWR VGND sg13g2_decap_4
X_1031_ net798 net685 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
X_1100_ net804 net663 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_21_128 VPWR VGND sg13g2_decap_8
XFILLER_21_139 VPWR VGND sg13g2_fill_1
Xinput96 Tile_X0Y0_FrameData[22] net96 VPWR VGND sg13g2_buf_1
Xinput85 Tile_X0Y0_FrameData[12] net85 VPWR VGND sg13g2_buf_1
Xinput63 Tile_X0Y0_E6END[7] net63 VPWR VGND sg13g2_buf_1
Xinput74 Tile_X0Y0_EE4END[2] net74 VPWR VGND sg13g2_buf_1
Xinput41 Tile_X0Y0_E2END[3] net41 VPWR VGND sg13g2_buf_1
Xinput52 Tile_X0Y0_E2MID[6] net52 VPWR VGND sg13g2_buf_1
Xinput30 DOUT_SRAM6 net30 VPWR VGND sg13g2_buf_1
X_0746_ _0188_ VPWR _0189_ VGND _0021_ _0160_ sg13g2_o21ai_1
X_0815_ _0033_ _0084_ _0252_ VPWR VGND sg13g2_nor2_1
XFILLER_96_194 VPWR VGND sg13g2_fill_2
XFILLER_88_139 VPWR VGND sg13g2_fill_2
X_0677_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit11.Q net2
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG7 _0158_ net635
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit10.Q Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG8
+ VPWR VGND sg13g2_mux4_1
X_1229_ net762 net717 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
X_0531_ net48 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit2.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit3.Q _0096_ VPWR
+ VGND sg13g2_nor3_1
X_0600_ VGND VPWR _0018_ _0151_ _0155_ _0154_ sg13g2_a21oi_1
X_1580_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb5 net434 VPWR
+ VGND sg13g2_buf_1
XFILLER_22_90 VPWR VGND sg13g2_decap_8
X_0393_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit0.Q net52
+ net44 net62 net630 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit1.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG1 VPWR VGND sg13g2_mux4_1
X_0462_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit18.Q net17
+ net21 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG9 net630 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit19.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG6 VPWR VGND sg13g2_mux4_1
X_1014_ net783 net700 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_118_27 VPWR VGND sg13g2_decap_8
X_0729_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit20.Q net142
+ net184 net177 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG12
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit21.Q net298 VPWR
+ VGND sg13g2_mux4_1
XFILLER_43_45 VPWR VGND sg13g2_fill_1
XFILLER_4_157 VPWR VGND sg13g2_decap_8
Xinput242 Tile_X0Y1_N2MID[7] net242 VPWR VGND sg13g2_buf_1
Xinput231 Tile_X0Y1_N2END[4] net231 VPWR VGND sg13g2_buf_1
Xinput220 Tile_X0Y1_FrameData[8] net220 VPWR VGND sg13g2_buf_1
X_1701_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG2 net557 VPWR
+ VGND sg13g2_buf_1
X_1494_ net801 net340 VPWR VGND sg13g2_buf_1
X_1563_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W1BEG0 net417 VPWR
+ VGND sg13g2_buf_1
X_0514_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit8.Q net77
+ net70 net61 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG5 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit9.Q
+ net275 VPWR VGND sg13g2_mux4_1
XFILLER_69_4 VPWR VGND sg13g2_fill_1
X_1632_ net203 net478 VPWR VGND sg13g2_buf_1
X_0376_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit4.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END2
+ net249 net116 net136 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit5.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG14 VPWR VGND sg13g2_mux4_1
XFILLER_81_112 VPWR VGND sg13g2_fill_2
X_0445_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit24.Q net11
+ net20 net630 net624 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit25.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb1 VPWR VGND sg13g2_mux4_1
XFILLER_13_59 VPWR VGND sg13g2_fill_1
XFILLER_1_105 VPWR VGND sg13g2_decap_8
XFILLER_72_167 VPWR VGND sg13g2_fill_1
XFILLER_57_153 VPWR VGND sg13g2_fill_1
X_0994_ net793 net697 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_74_2 VPWR VGND sg13g2_fill_1
Xoutput502 net502 Tile_X0Y1_S2BEG[1] VPWR VGND sg13g2_buf_1
X_1546_ Tile_X0Y1_N4END[8] net400 VPWR VGND sg13g2_buf_1
XFILLER_117_169 VPWR VGND sg13g2_decap_8
X_1477_ net788 net353 VPWR VGND sg13g2_buf_1
Xoutput568 net568 Tile_X0Y1_WW4BEG[12] VPWR VGND sg13g2_buf_1
Xoutput546 net546 Tile_X0Y1_W2BEGb[1] VPWR VGND sg13g2_buf_1
Xoutput579 net579 Tile_X0Y1_WW4BEG[8] VPWR VGND sg13g2_buf_1
X_1615_ net755 net491 VPWR VGND sg13g2_buf_1
Xoutput535 net535 Tile_X0Y1_W1BEG[2] VPWR VGND sg13g2_buf_1
Xoutput513 net513 Tile_X0Y1_S2BEGb[4] VPWR VGND sg13g2_buf_1
Xoutput524 net524 Tile_X0Y1_S4BEG[1] VPWR VGND sg13g2_buf_1
Xoutput557 net557 Tile_X0Y1_W6BEG[2] VPWR VGND sg13g2_buf_1
X_0359_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit26.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit27.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END1 _0058_ VPWR VGND sg13g2_nor3_1
X_0428_ net223 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit24.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit25.Q _0089_ VPWR
+ VGND sg13g2_nor3_1
XFILLER_116_180 VPWR VGND sg13g2_decap_4
XFILLER_108_125 VPWR VGND sg13g2_decap_4
XFILLER_40_68 VPWR VGND sg13g2_fill_2
Xfanout795 net100 net795 VPWR VGND sg13g2_buf_1
Xfanout784 net111 net784 VPWR VGND sg13g2_buf_1
XFILLER_65_32 VPWR VGND sg13g2_fill_2
XFILLER_1_18 VPWR VGND sg13g2_fill_2
Xfanout751 net220 net751 VPWR VGND sg13g2_buf_1
Xfanout740 net741 net740 VPWR VGND sg13g2_buf_1
Xfanout773 net198 net773 VPWR VGND sg13g2_buf_1
Xfanout762 net209 net762 VPWR VGND sg13g2_buf_1
X_1331_ net768 net681 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
X_1400_ net774 net662 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
X_1262_ net208 net708 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
Xinput6 DOUT_SRAM12 net6 VPWR VGND sg13g2_buf_1
XFILLER_36_112 VPWR VGND sg13g2_fill_1
XFILLER_36_134 VPWR VGND sg13g2_fill_1
X_1193_ net214 net728 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_51_137 VPWR VGND sg13g2_fill_2
X_0977_ net86 net710 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
Xoutput343 net343 Tile_X0Y0_FrameData_O[23] VPWR VGND sg13g2_buf_1
Xoutput332 net332 Tile_X0Y0_FrameData_O[13] VPWR VGND sg13g2_buf_1
Xoutput310 net310 DIN_SRAM23 VPWR VGND sg13g2_buf_1
Xoutput321 net321 DIN_SRAM5 VPWR VGND sg13g2_buf_1
Xoutput376 net376 Tile_X0Y0_FrameStrobe_O[6] VPWR VGND sg13g2_buf_1
Xoutput398 net398 Tile_X0Y0_N2BEGb[6] VPWR VGND sg13g2_buf_1
Xoutput387 net387 Tile_X0Y0_N2BEG[3] VPWR VGND sg13g2_buf_1
Xoutput365 net365 Tile_X0Y0_FrameStrobe_O[14] VPWR VGND sg13g2_buf_1
X_1529_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1BEG3 net383 VPWR
+ VGND sg13g2_buf_1
Xoutput354 net354 Tile_X0Y0_FrameData_O[4] VPWR VGND sg13g2_buf_1
XFILLER_19_58 VPWR VGND sg13g2_fill_1
XFILLER_27_178 VPWR VGND sg13g2_fill_2
XFILLER_51_12 VPWR VGND sg13g2_fill_2
XFILLER_116_60 VPWR VGND sg13g2_decap_8
XFILLER_18_101 VPWR VGND sg13g2_fill_1
XFILLER_18_123 VPWR VGND sg13g2_fill_1
X_0900_ net795 net732 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_92_74 VPWR VGND sg13g2_fill_2
X_0762_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG6 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG10
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit8.Q _0204_ VPWR
+ VGND sg13g2_mux2_1
X_0693_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit25.Q net637
+ _0171_ VPWR VGND Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit24.Q
+ sg13g2_nand3b_1
X_0831_ net154 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit0.Q
+ _0267_ VPWR VGND sg13g2_and2_1
X_1314_ net753 net693 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
X_1245_ net779 net717 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
X_1176_ net774 net740 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_24_126 VPWR VGND sg13g2_fill_2
XFILLER_102_95 VPWR VGND sg13g2_fill_2
XFILLER_15_148 VPWR VGND sg13g2_fill_1
XFILLER_87_85 VPWR VGND sg13g2_fill_1
XFILLER_87_63 VPWR VGND sg13g2_fill_1
X_1030_ net797 net688 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
Xinput31 DOUT_SRAM7 net31 VPWR VGND sg13g2_buf_1
Xinput20 DOUT_SRAM25 net20 VPWR VGND sg13g2_buf_1
XFILLER_21_107 VPWR VGND sg13g2_decap_4
X_0814_ VGND VPWR _0034_ _0250_ _0251_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit17.Q
+ sg13g2_a21oi_1
Xinput97 Tile_X0Y0_FrameData[23] net97 VPWR VGND sg13g2_buf_1
Xinput86 Tile_X0Y0_FrameData[13] net86 VPWR VGND sg13g2_buf_1
Xinput64 Tile_X0Y0_E6END[8] net64 VPWR VGND sg13g2_buf_1
Xinput75 Tile_X0Y0_EE4END[3] net75 VPWR VGND sg13g2_buf_1
Xinput42 Tile_X0Y0_E2END[4] net42 VPWR VGND sg13g2_buf_1
Xinput53 Tile_X0Y0_E2MID[7] net53 VPWR VGND sg13g2_buf_1
X_0676_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit8.Q net31
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG4 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG8
+ net637 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit9.Q Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG7
+ VPWR VGND sg13g2_mux4_1
X_0745_ VPWR _0188_ _0187_ VGND sg13g2_inv_1
X_1228_ net761 net718 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
X_1159_ net798 net645 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_32_47 VPWR VGND sg13g2_fill_1
XFILLER_11_173 VPWR VGND sg13g2_fill_1
X_0530_ VGND VPWR Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit0.Q
+ _0094_ _0095_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit1.Q
+ net257 _0039_ sg13g2_a221oi_1
XFILLER_11_195 VPWR VGND sg13g2_fill_2
X_0461_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit26.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END1
+ net248 net115 net135 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit27.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG9 VPWR VGND sg13g2_mux4_1
X_0392_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit11.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb1
+ net127 net236 net119 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit10.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG1 VPWR VGND sg13g2_mux4_1
XFILLER_93_176 VPWR VGND sg13g2_fill_2
XFILLER_93_165 VPWR VGND sg13g2_fill_1
X_1013_ net782 net700 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
X_0659_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit16.Q net223
+ net243 _0088_ net138 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit17.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG4 VPWR VGND sg13g2_mux4_1
X_0728_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit18.Q net183
+ net176 net164 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG11
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit19.Q net297 VPWR
+ VGND sg13g2_mux4_1
XFILLER_84_143 VPWR VGND sg13g2_fill_1
Xinput243 Tile_X0Y1_N4END[0] net243 VPWR VGND sg13g2_buf_1
Xinput232 Tile_X0Y1_N2END[5] net232 VPWR VGND sg13g2_buf_1
Xinput221 Tile_X0Y1_FrameData[9] net221 VPWR VGND sg13g2_buf_1
Xinput210 Tile_X0Y1_FrameData[28] net210 VPWR VGND sg13g2_buf_1
X_1700_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG1 net556 VPWR
+ VGND sg13g2_buf_1
X_1631_ net202 net477 VPWR VGND sg13g2_buf_1
X_1562_ Tile_X0Y1_UserCLK net416 VPWR VGND sg13g2_buf_1
X_1493_ net92 net338 VPWR VGND sg13g2_buf_1
X_0444_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit22.Q net10
+ net19 net631 net623 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit23.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb0 VPWR VGND sg13g2_mux4_1
X_0513_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit6.Q net76
+ net69 net60 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG4 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit7.Q
+ net274 VPWR VGND sg13g2_mux4_1
XFILLER_66_176 VPWR VGND sg13g2_fill_1
X_0375_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit15.Q net144
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG14 net170 _0070_
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit14.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END2
+ VPWR VGND sg13g2_mux4_1
XFILLER_81_168 VPWR VGND sg13g2_fill_2
XFILLER_57_121 VPWR VGND sg13g2_decap_4
XFILLER_54_12 VPWR VGND sg13g2_fill_2
XFILLER_110_40 VPWR VGND sg13g2_fill_2
XFILLER_95_96 VPWR VGND sg13g2_fill_2
XFILLER_0_161 VPWR VGND sg13g2_decap_8
XFILLER_0_194 VPWR VGND sg13g2_decap_8
X_0993_ net792 net699 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_81_4 VPWR VGND sg13g2_fill_1
X_1614_ net756 net490 VPWR VGND sg13g2_buf_1
Xoutput536 net536 Tile_X0Y1_W1BEG[3] VPWR VGND sg13g2_buf_1
Xoutput503 net503 Tile_X0Y1_S2BEG[2] VPWR VGND sg13g2_buf_1
Xoutput514 net514 Tile_X0Y1_S2BEGb[5] VPWR VGND sg13g2_buf_1
Xoutput525 net525 Tile_X0Y1_S4BEG[2] VPWR VGND sg13g2_buf_1
X_0427_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit27.Q net34
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG12 net64 _0087_
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit26.Q _0088_ VPWR
+ VGND sg13g2_mux4_1
X_1476_ net791 net350 VPWR VGND sg13g2_buf_1
Xoutput558 net558 Tile_X0Y1_W6BEG[3] VPWR VGND sg13g2_buf_1
Xoutput569 net569 Tile_X0Y1_WW4BEG[13] VPWR VGND sg13g2_buf_1
Xoutput547 net547 Tile_X0Y1_W2BEGb[2] VPWR VGND sg13g2_buf_1
XFILLER_39_110 VPWR VGND sg13g2_fill_2
X_1545_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb7 net399 VPWR
+ VGND sg13g2_buf_1
X_0358_ _0057_ net115 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit26.Q
+ VPWR VGND sg13g2_nand2b_1
XFILLER_108_148 VPWR VGND sg13g2_fill_2
XFILLER_108_137 VPWR VGND sg13g2_fill_2
XFILLER_49_12 VPWR VGND sg13g2_fill_1
Xfanout796 net99 net796 VPWR VGND sg13g2_buf_1
Xfanout785 net110 net785 VPWR VGND sg13g2_buf_1
Xfanout752 net219 net752 VPWR VGND sg13g2_buf_1
Xfanout730 net737 net730 VPWR VGND sg13g2_buf_1
Xfanout741 net742 net741 VPWR VGND sg13g2_buf_1
Xfanout774 net197 net774 VPWR VGND sg13g2_buf_1
Xfanout763 net208 net763 VPWR VGND sg13g2_buf_1
XFILLER_121_94 VPWR VGND sg13g2_decap_8
X_1261_ net209 net708 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
X_1330_ net767 net683 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
Xinput7 DOUT_SRAM13 net7 VPWR VGND sg13g2_buf_1
X_1192_ net781 net739 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
X_0976_ net808 net713 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
Xoutput377 net377 Tile_X0Y0_FrameStrobe_O[7] VPWR VGND sg13g2_buf_1
Xoutput366 net366 Tile_X0Y0_FrameStrobe_O[15] VPWR VGND sg13g2_buf_1
Xoutput344 net344 Tile_X0Y0_FrameData_O[24] VPWR VGND sg13g2_buf_1
Xoutput355 net355 Tile_X0Y0_FrameData_O[5] VPWR VGND sg13g2_buf_1
Xoutput333 net333 Tile_X0Y0_FrameData_O[14] VPWR VGND sg13g2_buf_1
Xoutput311 net311 DIN_SRAM24 VPWR VGND sg13g2_buf_1
Xoutput300 net300 DIN_SRAM14 VPWR VGND sg13g2_buf_1
Xoutput322 net322 DIN_SRAM6 VPWR VGND sg13g2_buf_1
XFILLER_10_28 VPWR VGND sg13g2_fill_2
Xoutput388 net388 Tile_X0Y0_N2BEG[4] VPWR VGND sg13g2_buf_1
Xoutput399 net399 Tile_X0Y0_N2BEGb[7] VPWR VGND sg13g2_buf_1
X_1528_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1BEG2 net382 VPWR
+ VGND sg13g2_buf_1
X_1459_ net203 net641 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_42_105 VPWR VGND sg13g2_decap_8
XFILLER_42_116 VPWR VGND sg13g2_fill_2
XFILLER_51_35 VPWR VGND sg13g2_decap_4
XFILLER_76_21 VPWR VGND sg13g2_fill_1
XFILLER_33_127 VPWR VGND sg13g2_fill_2
X_0830_ _0265_ VPWR _0266_ VGND _0000_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit0.Q
+ sg13g2_o21ai_1
X_0692_ _0168_ VPWR net253 VGND Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit23.Q
+ _0170_ sg13g2_o21ai_1
X_0761_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit9.Q VPWR
+ _0203_ VGND Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit8.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG14 sg13g2_o21ai_1
XFILLER_110_143 VPWR VGND sg13g2_fill_1
XFILLER_2_84 VPWR VGND sg13g2_decap_8
X_1313_ net752 net695 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
X_1244_ net778 net715 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
X_1175_ net773 net740 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
X_0959_ net789 net709 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_46_35 VPWR VGND sg13g2_fill_2
Xinput54 Tile_X0Y0_E6END[0] net54 VPWR VGND sg13g2_buf_1
Xinput43 Tile_X0Y0_E2END[5] net43 VPWR VGND sg13g2_buf_1
Xinput32 DOUT_SRAM8 net32 VPWR VGND sg13g2_buf_1
Xinput10 DOUT_SRAM16 net10 VPWR VGND sg13g2_buf_1
Xinput21 DOUT_SRAM26 net21 VPWR VGND sg13g2_buf_1
X_0813_ net145 net180 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit15.Q
+ _0250_ VPWR VGND sg13g2_mux2_1
Xinput98 Tile_X0Y0_FrameData[24] net98 VPWR VGND sg13g2_buf_1
Xinput87 Tile_X0Y0_FrameData[14] net87 VPWR VGND sg13g2_buf_1
Xinput65 Tile_X0Y0_E6END[9] net65 VPWR VGND sg13g2_buf_1
Xinput76 Tile_X0Y0_EE4END[4] net76 VPWR VGND sg13g2_buf_1
X_0675_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit6.Q net30
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG5 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG9
+ net638 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit7.Q Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG6
+ VPWR VGND sg13g2_mux4_1
X_0744_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit6.Q VPWR
+ _0187_ VGND net173 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit5.Q
+ sg13g2_o21ai_1
XFILLER_35_0 VPWR VGND sg13g2_fill_2
X_1158_ net98 net644 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_96_196 VPWR VGND sg13g2_fill_1
X_1227_ net760 net718 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
X_1089_ net792 net664 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_79_108 VPWR VGND sg13g2_fill_2
XFILLER_57_56 VPWR VGND sg13g2_fill_2
XFILLER_73_88 VPWR VGND sg13g2_fill_2
XFILLER_73_66 VPWR VGND sg13g2_fill_1
X_0460_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit16.Q net16
+ net19 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG10 net629
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit17.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG5
+ VPWR VGND sg13g2_mux4_1
XFILLER_7_189 VPWR VGND sg13g2_fill_1
X_1012_ net812 net701 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_93_111 VPWR VGND sg13g2_fill_1
X_0391_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit20.Q net160
+ net152 net170 _0078_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit21.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb1 VPWR VGND sg13g2_mux4_1
XFILLER_93_199 VPWR VGND sg13g2_fill_2
XFILLER_8_94 VPWR VGND sg13g2_fill_1
XFILLER_8_72 VPWR VGND sg13g2_decap_4
X_0727_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit16.Q net182
+ net175 net163 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG10
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit17.Q net296 VPWR
+ VGND sg13g2_mux4_1
X_0589_ net624 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit24.Q
+ _0145_ VPWR VGND sg13g2_nor2b_1
X_0658_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit14.Q net30
+ net4 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG5 net634 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit15.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG10 VPWR VGND sg13g2_mux4_1
XFILLER_84_199 VPWR VGND sg13g2_fill_2
XFILLER_111_4 VPWR VGND sg13g2_fill_1
XFILLER_68_11 VPWR VGND sg13g2_fill_2
XFILLER_68_77 VPWR VGND sg13g2_fill_1
XFILLER_68_55 VPWR VGND sg13g2_fill_1
Xinput233 Tile_X0Y1_N2END[6] net233 VPWR VGND sg13g2_buf_1
Xinput244 Tile_X0Y1_N4END[1] net244 VPWR VGND sg13g2_buf_1
Xinput222 Tile_X0Y1_FrameStrobe[8] net222 VPWR VGND sg13g2_buf_1
Xinput200 Tile_X0Y1_FrameData[19] net200 VPWR VGND sg13g2_buf_1
Xinput211 Tile_X0Y1_FrameData[29] net211 VPWR VGND sg13g2_buf_1
XFILLER_75_199 VPWR VGND sg13g2_fill_2
XFILLER_16_200 VPWR VGND sg13g2_fill_1
XFILLER_83_8 VPWR VGND sg13g2_fill_2
X_1630_ net771 net475 VPWR VGND sg13g2_buf_1
X_1492_ net804 net337 VPWR VGND sg13g2_buf_1
X_0512_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit4.Q net75
+ net68 net59 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG3 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit5.Q
+ net272 VPWR VGND sg13g2_mux4_1
X_1561_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N4BEG3 net406 VPWR
+ VGND sg13g2_buf_1
X_0443_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit20.Q net18
+ net27 net631 net623 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit21.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG7 VPWR VGND sg13g2_mux4_1
XFILLER_3_192 VPWR VGND sg13g2_fill_1
XFILLER_3_181 VPWR VGND sg13g2_decap_8
X_0374_ VGND VPWR _0069_ _0068_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit29.Q
+ _0008_ _0070_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit28.Q
+ sg13g2_a221oi_1
XFILLER_66_122 VPWR VGND sg13g2_fill_2
XFILLER_119_94 VPWR VGND sg13g2_decap_8
XFILLER_63_136 VPWR VGND sg13g2_fill_1
XFILLER_0_173 VPWR VGND sg13g2_decap_8
X_0992_ net790 net698 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_44_90 VPWR VGND sg13g2_fill_1
Xoutput559 net559 Tile_X0Y1_W6BEG[4] VPWR VGND sg13g2_buf_1
Xoutput548 net548 Tile_X0Y1_W2BEGb[3] VPWR VGND sg13g2_buf_1
XFILLER_5_40 VPWR VGND sg13g2_fill_2
Xoutput537 net537 Tile_X0Y1_W2BEG[0] VPWR VGND sg13g2_buf_1
Xoutput504 net504 Tile_X0Y1_S2BEG[3] VPWR VGND sg13g2_buf_1
Xoutput515 net515 Tile_X0Y1_S2BEGb[6] VPWR VGND sg13g2_buf_1
Xoutput526 net526 Tile_X0Y1_S4BEG[3] VPWR VGND sg13g2_buf_1
X_1613_ net759 net487 VPWR VGND sg13g2_buf_1
X_1544_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb6 net398 VPWR
+ VGND sg13g2_buf_1
X_0426_ VGND VPWR _0085_ _0086_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit25.Q
+ _0006_ _0087_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit24.Q
+ sg13g2_a221oi_1
X_1475_ net802 net339 VPWR VGND sg13g2_buf_1
X_0357_ VGND VPWR Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit31.Q
+ _0052_ net326 _0056_ sg13g2_a21oi_1
Xfanout720 net724 net720 VPWR VGND sg13g2_buf_1
Xfanout742 net749 net742 VPWR VGND sg13g2_buf_1
Xfanout731 net737 net731 VPWR VGND sg13g2_buf_1
Xfanout786 net109 net786 VPWR VGND sg13g2_buf_1
Xfanout797 net98 net797 VPWR VGND sg13g2_buf_1
XFILLER_65_12 VPWR VGND sg13g2_fill_2
Xfanout753 net218 net753 VPWR VGND sg13g2_buf_1
Xfanout775 net196 net775 VPWR VGND sg13g2_buf_1
Xfanout764 net207 net764 VPWR VGND sg13g2_buf_1
XFILLER_121_73 VPWR VGND sg13g2_decap_8
XFILLER_60_117 VPWR VGND sg13g2_fill_2
XFILLER_14_71 VPWR VGND sg13g2_fill_2
Xinput8 DOUT_SRAM14 net8 VPWR VGND sg13g2_buf_1
X_1191_ net770 net739 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
X_1260_ net761 net706 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_46_8 VPWR VGND sg13g2_fill_2
XFILLER_51_106 VPWR VGND sg13g2_decap_8
XFILLER_51_117 VPWR VGND sg13g2_fill_1
XFILLER_51_139 VPWR VGND sg13g2_fill_1
X_0975_ net807 net713 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
Xoutput378 net378 Tile_X0Y0_FrameStrobe_O[8] VPWR VGND sg13g2_buf_1
Xoutput389 net389 Tile_X0Y0_N2BEG[5] VPWR VGND sg13g2_buf_1
Xoutput367 net367 Tile_X0Y0_FrameStrobe_O[16] VPWR VGND sg13g2_buf_1
XFILLER_113_130 VPWR VGND sg13g2_decap_8
Xoutput345 net345 Tile_X0Y0_FrameData_O[25] VPWR VGND sg13g2_buf_1
Xoutput334 net334 Tile_X0Y0_FrameData_O[15] VPWR VGND sg13g2_buf_1
X_1527_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1BEG1 net381 VPWR
+ VGND sg13g2_buf_1
Xoutput356 net356 Tile_X0Y0_FrameData_O[6] VPWR VGND sg13g2_buf_1
Xoutput312 net312 DIN_SRAM25 VPWR VGND sg13g2_buf_1
Xoutput301 net301 DIN_SRAM15 VPWR VGND sg13g2_buf_1
Xoutput323 net323 DIN_SRAM7 VPWR VGND sg13g2_buf_1
X_0409_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit12.Q net35
+ net48 net40 net625 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit13.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG5 VPWR VGND sg13g2_mux4_1
X_1389_ net762 net658 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
X_1458_ net204 net642 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_116_95 VPWR VGND sg13g2_decap_8
XFILLER_92_76 VPWR VGND sg13g2_fill_1
XFILLER_92_54 VPWR VGND sg13g2_fill_2
XFILLER_76_77 VPWR VGND sg13g2_fill_2
XFILLER_41_150 VPWR VGND sg13g2_fill_1
X_0760_ _0023_ _0079_ _0202_ VPWR VGND sg13g2_nor2_1
X_0691_ VGND VPWR net148 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit22.Q
+ _0170_ _0169_ sg13g2_a21oi_1
XFILLER_110_199 VPWR VGND sg13g2_fill_2
X_1174_ net772 net739 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_2_63 VPWR VGND sg13g2_decap_8
X_1312_ net751 net692 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
X_1243_ net777 net715 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
X_0958_ net813 net722 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
X_0889_ net109 net746 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_15_139 VPWR VGND sg13g2_decap_8
XFILLER_11_83 VPWR VGND sg13g2_decap_8
XFILLER_36_80 VPWR VGND sg13g2_fill_1
Xinput88 Tile_X0Y0_FrameData[15] net88 VPWR VGND sg13g2_buf_1
Xinput77 Tile_X0Y0_EE4END[5] net77 VPWR VGND sg13g2_buf_1
Xinput55 Tile_X0Y0_E6END[10] net55 VPWR VGND sg13g2_buf_1
Xinput66 Tile_X0Y0_EE4END[0] net66 VPWR VGND sg13g2_buf_1
Xinput44 Tile_X0Y0_E2END[6] net44 VPWR VGND sg13g2_buf_1
Xinput11 DOUT_SRAM17 net11 VPWR VGND sg13g2_buf_1
Xinput33 DOUT_SRAM9 net33 VPWR VGND sg13g2_buf_1
XFILLER_14_194 VPWR VGND sg13g2_fill_2
Xinput22 DOUT_SRAM27 net22 VPWR VGND sg13g2_buf_1
X_0743_ VGND VPWR _0179_ _0181_ Tile_X0Y0_IHP_SRAM_top.N4BEG_outbuf_8.A _0186_ sg13g2_a21oi_1
X_0812_ _0248_ VPWR _0249_ VGND _0033_ _0158_ sg13g2_o21ai_1
Xinput99 Tile_X0Y0_FrameData[25] net99 VPWR VGND sg13g2_buf_1
X_0674_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit5.Q net29
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG10 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG6
+ net639 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit4.Q Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG5
+ VPWR VGND sg13g2_mux4_1
X_1157_ net796 net644 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
X_1226_ net213 net718 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
X_1088_ net790 net667 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
X_0390_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit10.Q net236
+ net228 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG1 net127 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit11.Q
+ _0078_ VPWR VGND sg13g2_mux4_1
X_1011_ net811 net701 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_93_101 VPWR VGND sg13g2_decap_4
X_0726_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit14.Q net181
+ net189 net173 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG9
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit15.Q net325 VPWR
+ VGND sg13g2_mux4_1
X_0588_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG6 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG10
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit24.Q _0144_ VPWR
+ VGND sg13g2_mux2_1
X_0657_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit18.Q net224
+ net244 _0060_ net139 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit19.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG5 VPWR VGND sg13g2_mux4_1
X_1209_ net196 net728 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_104_4 VPWR VGND sg13g2_fill_1
Xinput201 Tile_X0Y1_FrameData[1] net201 VPWR VGND sg13g2_buf_1
XFILLER_90_137 VPWR VGND sg13g2_fill_1
XFILLER_90_115 VPWR VGND sg13g2_fill_1
Xinput223 Tile_X0Y1_N1END[0] net223 VPWR VGND sg13g2_buf_1
Xinput234 Tile_X0Y1_N2END[7] net234 VPWR VGND sg13g2_buf_1
Xinput245 Tile_X0Y1_N4END[2] net245 VPWR VGND sg13g2_buf_1
Xinput212 Tile_X0Y1_FrameData[2] net212 VPWR VGND sg13g2_buf_1
XFILLER_90_159 VPWR VGND sg13g2_fill_2
X_0511_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit2.Q net74
+ net67 net58 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG2 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit3.Q
+ net271 VPWR VGND sg13g2_mux4_1
X_1560_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N4BEG2 net405 VPWR
+ VGND sg13g2_buf_1
X_1491_ net805 net336 VPWR VGND sg13g2_buf_1
X_0442_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit18.Q net17
+ net26 net630 net624 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit19.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG6 VPWR VGND sg13g2_mux4_1
XFILLER_3_160 VPWR VGND sg13g2_decap_8
X_0373_ _0069_ _0067_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit28.Q
+ VPWR VGND sg13g2_nand2b_1
XFILLER_95_0 VPWR VGND sg13g2_fill_1
X_1689_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG6 net543 VPWR
+ VGND sg13g2_buf_1
X_0709_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit12.Q net174
+ net188 net172 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG8
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit13.Q net291 VPWR
+ VGND sg13g2_mux4_1
XFILLER_72_104 VPWR VGND sg13g2_decap_4
XFILLER_110_64 VPWR VGND sg13g2_fill_1
XFILLER_119_73 VPWR VGND sg13g2_decap_8
XFILLER_119_62 VPWR VGND sg13g2_decap_8
XFILLER_48_123 VPWR VGND sg13g2_fill_2
XFILLER_48_156 VPWR VGND sg13g2_fill_1
X_0991_ net789 net698 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_71_192 VPWR VGND sg13g2_fill_1
X_1474_ net813 net328 VPWR VGND sg13g2_buf_1
X_1543_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb5 net397 VPWR
+ VGND sg13g2_buf_1
Xoutput549 net549 Tile_X0Y1_W2BEGb[4] VPWR VGND sg13g2_buf_1
Xoutput538 net538 Tile_X0Y1_W2BEG[1] VPWR VGND sg13g2_buf_1
Xoutput505 net505 Tile_X0Y1_S2BEG[4] VPWR VGND sg13g2_buf_1
Xoutput516 net516 Tile_X0Y1_S2BEGb[7] VPWR VGND sg13g2_buf_1
Xoutput527 net527 Tile_X0Y1_S4BEG[4] VPWR VGND sg13g2_buf_1
X_1612_ net201 net476 VPWR VGND sg13g2_buf_1
X_0425_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit24.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit25.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END0 _0086_ VPWR VGND sg13g2_nor3_1
X_0356_ net1 VPWR _0056_ VGND Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit31.Q
+ _0055_ sg13g2_o21ai_1
XFILLER_116_161 VPWR VGND sg13g2_fill_2
Xfanout710 net713 net710 VPWR VGND sg13g2_buf_1
Xfanout721 net724 net721 VPWR VGND sg13g2_buf_1
Xfanout732 net736 net732 VPWR VGND sg13g2_buf_1
Xfanout743 net748 net743 VPWR VGND sg13g2_buf_1
Xfanout754 net217 net754 VPWR VGND sg13g2_buf_1
Xfanout776 net195 net776 VPWR VGND sg13g2_buf_1
Xfanout765 net206 net765 VPWR VGND sg13g2_buf_1
XFILLER_121_52 VPWR VGND sg13g2_decap_8
Xfanout787 net108 net787 VPWR VGND sg13g2_buf_1
Xfanout798 net97 net798 VPWR VGND sg13g2_buf_1
XFILLER_65_79 VPWR VGND sg13g2_fill_1
XFILLER_65_68 VPWR VGND sg13g2_decap_8
XFILLER_14_94 VPWR VGND sg13g2_decap_8
XFILLER_107_161 VPWR VGND sg13g2_fill_2
Xinput9 DOUT_SRAM15 net9 VPWR VGND sg13g2_buf_1
X_1190_ net759 net739 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
X_0974_ net806 net711 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
Xoutput379 net379 Tile_X0Y0_FrameStrobe_O[9] VPWR VGND sg13g2_buf_1
Xoutput368 net368 Tile_X0Y0_FrameStrobe_O[17] VPWR VGND sg13g2_buf_1
Xoutput346 net346 Tile_X0Y0_FrameData_O[26] VPWR VGND sg13g2_buf_1
Xoutput335 net335 Tile_X0Y0_FrameData_O[16] VPWR VGND sg13g2_buf_1
Xoutput357 net357 Tile_X0Y0_FrameData_O[7] VPWR VGND sg13g2_buf_1
X_1526_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1BEG0 net380 VPWR
+ VGND sg13g2_buf_1
Xoutput313 net313 DIN_SRAM26 VPWR VGND sg13g2_buf_1
Xoutput302 net302 DIN_SRAM16 VPWR VGND sg13g2_buf_1
Xoutput324 net324 DIN_SRAM8 VPWR VGND sg13g2_buf_1
X_1457_ net205 net642 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
X_0339_ VPWR _0042_ net627 VGND sg13g2_inv_1
X_0408_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit6.Q net49
+ net41 net59 net627 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit7.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG4 VPWR VGND sg13g2_mux4_1
X_1388_ net761 net658 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_27_126 VPWR VGND sg13g2_decap_4
XFILLER_35_27 VPWR VGND sg13g2_fill_2
XFILLER_116_74 VPWR VGND sg13g2_decap_8
XFILLER_104_142 VPWR VGND sg13g2_fill_1
X_0690_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit22.Q net156
+ _0169_ VPWR VGND sg13g2_nor2b_1
X_1311_ net750 net693 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
X_1173_ net771 net739 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_2_42 VPWR VGND sg13g2_decap_8
X_1242_ net776 net716 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_32_140 VPWR VGND sg13g2_fill_1
X_0957_ net802 net722 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
X_0888_ net110 net745 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
X_1509_ net710 net373 VPWR VGND sg13g2_buf_1
XFILLER_102_65 VPWR VGND sg13g2_fill_1
XFILLER_62_25 VPWR VGND sg13g2_fill_2
XFILLER_62_14 VPWR VGND sg13g2_decap_8
XFILLER_46_37 VPWR VGND sg13g2_fill_1
Xinput89 Tile_X0Y0_FrameData[16] net89 VPWR VGND sg13g2_buf_1
Xinput56 Tile_X0Y0_E6END[11] net56 VPWR VGND sg13g2_buf_1
Xinput78 Tile_X0Y0_EE4END[6] net78 VPWR VGND sg13g2_buf_1
Xinput45 Tile_X0Y0_E2END[7] net45 VPWR VGND sg13g2_buf_1
Xinput67 Tile_X0Y0_EE4END[10] net67 VPWR VGND sg13g2_buf_1
Xinput34 Tile_X0Y0_E1END[0] net34 VPWR VGND sg13g2_buf_1
X_0673_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit3.Q net28
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG11 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG7
+ net640 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit2.Q Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG4
+ VPWR VGND sg13g2_mux4_1
Xinput12 DOUT_SRAM18 net12 VPWR VGND sg13g2_buf_1
Xinput23 DOUT_SRAM28 net23 VPWR VGND sg13g2_buf_1
X_0742_ VGND VPWR _0020_ _0184_ _0186_ _0185_ sg13g2_a21oi_1
X_0811_ VPWR _0248_ _0247_ VGND sg13g2_inv_1
XFILLER_35_2 VPWR VGND sg13g2_fill_1
X_1156_ net795 net644 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
X_1087_ net789 net667 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
X_1225_ net214 net718 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_87_198 VPWR VGND sg13g2_fill_2
XFILLER_113_97 VPWR VGND sg13g2_fill_2
XFILLER_98_21 VPWR VGND sg13g2_fill_1
XFILLER_11_154 VPWR VGND sg13g2_fill_2
X_1010_ net810 net697 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_78_198 VPWR VGND sg13g2_fill_2
X_0656_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit12.Q net29
+ net33 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG6 net633 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit13.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG9 VPWR VGND sg13g2_mux4_1
X_0725_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit12.Q net174
+ net188 net172 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG8
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit13.Q net324 VPWR
+ VGND sg13g2_mux4_1
X_0587_ _0141_ _0143_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S4BEG1
+ VPWR VGND sg13g2_nor2_1
XFILLER_69_198 VPWR VGND sg13g2_fill_2
X_1208_ net774 net730 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
X_1139_ net811 net652 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_108_20 VPWR VGND sg13g2_fill_2
XFILLER_4_128 VPWR VGND sg13g2_decap_4
XFILLER_108_86 VPWR VGND sg13g2_fill_1
XFILLER_68_35 VPWR VGND sg13g2_fill_2
XFILLER_68_13 VPWR VGND sg13g2_fill_1
Xinput213 Tile_X0Y1_FrameData[30] net213 VPWR VGND sg13g2_buf_1
Xinput224 Tile_X0Y1_N1END[1] net224 VPWR VGND sg13g2_buf_1
Xinput235 Tile_X0Y1_N2MID[0] net235 VPWR VGND sg13g2_buf_1
Xinput202 Tile_X0Y1_FrameData[20] net202 VPWR VGND sg13g2_buf_1
XFILLER_75_146 VPWR VGND sg13g2_fill_1
Xinput246 Tile_X0Y1_N4END[3] net246 VPWR VGND sg13g2_buf_1
XFILLER_33_71 VPWR VGND sg13g2_fill_1
X_0510_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit0.Q net73
+ net81 net57 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG1 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit1.Q
+ net270 VPWR VGND sg13g2_mux4_1
X_1490_ net806 net335 VPWR VGND sg13g2_buf_1
X_0441_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit16.Q net16
+ net24 net629 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG5 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit17.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG5 VPWR VGND sg13g2_mux4_1
XFILLER_66_124 VPWR VGND sg13g2_fill_1
X_0372_ net225 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit28.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit29.Q _0068_ VPWR
+ VGND sg13g2_nor3_1
X_0639_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit22.Q net30
+ net8 net639 net633 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit23.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb6 VPWR VGND sg13g2_mux4_1
X_1688_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG5 net542 VPWR
+ VGND sg13g2_buf_1
X_0708_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit10.Q net187
+ net180 net171 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG7
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit11.Q net290 VPWR
+ VGND sg13g2_mux4_1
XFILLER_57_113 VPWR VGND sg13g2_decap_4
XFILLER_119_41 VPWR VGND sg13g2_decap_8
XFILLER_48_146 VPWR VGND sg13g2_fill_2
X_0990_ net813 net712 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_60_91 VPWR VGND sg13g2_decap_4
X_1611_ net781 net465 VPWR VGND sg13g2_buf_1
X_1473_ Tile_X0Y1_UserCLK net293 VPWR VGND sg13g2_buf_1
X_0424_ _0085_ net114 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit24.Q
+ VPWR VGND sg13g2_nand2b_1
X_1542_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb4 net396 VPWR
+ VGND sg13g2_buf_1
XFILLER_5_97 VPWR VGND sg13g2_fill_2
XFILLER_5_31 VPWR VGND sg13g2_fill_1
Xoutput539 net539 Tile_X0Y1_W2BEG[2] VPWR VGND sg13g2_buf_1
Xoutput506 net506 Tile_X0Y1_S2BEG[5] VPWR VGND sg13g2_buf_1
Xoutput517 net517 Tile_X0Y1_S4BEG[0] VPWR VGND sg13g2_buf_1
Xoutput528 net528 Tile_X0Y1_S4BEG[5] VPWR VGND sg13g2_buf_1
X_0355_ _0054_ _0053_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit30.Q
+ _0055_ VPWR VGND sg13g2_mux2_1
XFILLER_116_184 VPWR VGND sg13g2_fill_1
Xfanout711 net713 net711 VPWR VGND sg13g2_buf_1
Xfanout788 net107 net788 VPWR VGND sg13g2_buf_1
Xfanout722 net724 net722 VPWR VGND sg13g2_buf_1
Xfanout733 net736 net733 VPWR VGND sg13g2_buf_1
Xfanout700 net701 net700 VPWR VGND sg13g2_buf_1
Xfanout799 net96 net799 VPWR VGND sg13g2_buf_1
Xfanout744 net747 net744 VPWR VGND sg13g2_buf_1
Xfanout755 net216 net755 VPWR VGND sg13g2_buf_1
Xfanout777 net194 net777 VPWR VGND sg13g2_buf_1
Xfanout766 net205 net766 VPWR VGND sg13g2_buf_1
XFILLER_121_31 VPWR VGND sg13g2_decap_8
XFILLER_65_25 VPWR VGND sg13g2_decap_8
XFILLER_60_119 VPWR VGND sg13g2_fill_1
XFILLER_91_200 VPWR VGND sg13g2_fill_1
X_0973_ net805 net711 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
Xoutput314 net314 DIN_SRAM27 VPWR VGND sg13g2_buf_1
Xoutput303 net303 DIN_SRAM17 VPWR VGND sg13g2_buf_1
Xoutput325 net325 DIN_SRAM9 VPWR VGND sg13g2_buf_1
X_1525_ Tile_X0Y1_FrameStrobe[19] net370 VPWR VGND sg13g2_buf_1
Xoutput369 net369 Tile_X0Y0_FrameStrobe_O[18] VPWR VGND sg13g2_buf_1
Xoutput336 net336 Tile_X0Y0_FrameData_O[17] VPWR VGND sg13g2_buf_1
Xoutput347 net347 Tile_X0Y0_FrameData_O[27] VPWR VGND sg13g2_buf_1
Xoutput358 net358 Tile_X0Y0_FrameData_O[8] VPWR VGND sg13g2_buf_1
X_0407_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit17.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb4
+ net130 net239 net122 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit16.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG4 VPWR VGND sg13g2_mux4_1
X_1387_ net760 net661 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
X_1456_ net765 net642 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_82_200 VPWR VGND sg13g2_fill_1
X_0338_ VPWR _0041_ net628 VGND sg13g2_inv_1
XFILLER_50_174 VPWR VGND sg13g2_fill_2
XFILLER_116_53 VPWR VGND sg13g2_decap_8
XFILLER_104_198 VPWR VGND sg13g2_fill_2
XFILLER_76_68 VPWR VGND sg13g2_fill_1
XFILLER_73_200 VPWR VGND sg13g2_fill_1
XFILLER_92_56 VPWR VGND sg13g2_fill_1
X_1310_ net780 net692 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
X_1241_ net775 net716 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
X_1172_ net769 net738 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_2_98 VPWR VGND sg13g2_decap_8
X_0956_ net104 net721 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_70_0 VPWR VGND sg13g2_fill_2
X_0887_ net111 net746 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
X_1508_ net721 net372 VPWR VGND sg13g2_buf_1
X_1439_ net750 net650 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
Xinput13 DOUT_SRAM19 net13 VPWR VGND sg13g2_buf_1
XFILLER_14_196 VPWR VGND sg13g2_fill_1
X_0810_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit16.Q VPWR
+ _0247_ VGND net171 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit15.Q
+ sg13g2_o21ai_1
Xinput57 Tile_X0Y0_E6END[1] net57 VPWR VGND sg13g2_buf_1
Xinput68 Tile_X0Y0_EE4END[11] net68 VPWR VGND sg13g2_buf_1
Xinput79 Tile_X0Y0_EE4END[7] net79 VPWR VGND sg13g2_buf_1
Xinput35 Tile_X0Y0_E1END[1] net35 VPWR VGND sg13g2_buf_1
Xinput46 Tile_X0Y0_E2MID[0] net46 VPWR VGND sg13g2_buf_1
Xinput24 DOUT_SRAM29 net24 VPWR VGND sg13g2_buf_1
X_0741_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit4.Q VPWR
+ _0185_ VGND _0182_ _0183_ sg13g2_o21ai_1
X_0672_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit0.Q net246
+ net141 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG8 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG12
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit1.Q Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG3
+ VPWR VGND sg13g2_mux4_1
XFILLER_96_133 VPWR VGND sg13g2_fill_2
XFILLER_96_111 VPWR VGND sg13g2_fill_1
X_1224_ net781 net729 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
X_1155_ net101 net644 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
X_1086_ net813 net679 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
X_0939_ net803 net721 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_20_166 VPWR VGND sg13g2_fill_2
XFILLER_57_15 VPWR VGND sg13g2_fill_1
XFILLER_7_115 VPWR VGND sg13g2_decap_4
XFILLER_0_0 VPWR VGND sg13g2_fill_1
X_0586_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit23.Q _0142_
+ _0143_ VPWR VGND sg13g2_nor2_1
X_0724_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit10.Q net187
+ net180 net171 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG7
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit11.Q net323 VPWR
+ VGND sg13g2_mux4_1
X_0655_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit20.Q net225
+ net245 _0067_ net140 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit21.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG6 VPWR VGND sg13g2_mux4_1
XFILLER_33_0 VPWR VGND sg13g2_fill_2
X_1207_ net773 net730 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
X_1138_ net810 net657 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
X_1069_ net90 net678 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_75_114 VPWR VGND sg13g2_decap_4
Xinput214 Tile_X0Y1_FrameData[31] net214 VPWR VGND sg13g2_buf_1
Xinput236 Tile_X0Y1_N2MID[1] net236 VPWR VGND sg13g2_buf_1
Xinput247 Tile_X0Y1_N4END[4] net247 VPWR VGND sg13g2_buf_1
Xinput225 Tile_X0Y1_N1END[2] net225 VPWR VGND sg13g2_buf_1
Xinput203 Tile_X0Y1_FrameData[21] net203 VPWR VGND sg13g2_buf_1
XFILLER_17_95 VPWR VGND sg13g2_fill_2
X_0440_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit14.Q net15
+ net23 net628 net627 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit15.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG4 VPWR VGND sg13g2_mux4_1
X_0371_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit30.Q net36
+ net55 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG14 _0066_
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit31.Q _0067_ VPWR
+ VGND sg13g2_mux4_1
X_0707_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit8.Q net186
+ net179 net170 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG6
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit9.Q net289 VPWR
+ VGND sg13g2_mux4_1
X_0569_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit24.Q net37
+ net56 net75 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG3 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit23.Q
+ _0128_ VPWR VGND sg13g2_mux4_1
X_0638_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit20.Q net29
+ net7 net638 net634 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit21.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb5 VPWR VGND sg13g2_mux4_1
X_1687_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG4 net541 VPWR
+ VGND sg13g2_buf_1
XFILLER_57_125 VPWR VGND sg13g2_fill_2
XFILLER_119_20 VPWR VGND sg13g2_decap_8
XFILLER_119_171 VPWR VGND sg13g2_decap_8
XFILLER_0_187 VPWR VGND sg13g2_decap_8
X_1610_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG15 net455 VPWR
+ VGND sg13g2_buf_1
Xoutput507 net507 Tile_X0Y1_S2BEG[6] VPWR VGND sg13g2_buf_1
Xoutput518 net518 Tile_X0Y1_S4BEG[10] VPWR VGND sg13g2_buf_1
X_0423_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit12.Q net46
+ net38 net54 net623 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit13.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG7 VPWR VGND sg13g2_mux4_1
X_1541_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb3 net395 VPWR
+ VGND sg13g2_buf_1
Xoutput529 net529 Tile_X0Y1_S4BEG[6] VPWR VGND sg13g2_buf_1
X_0354_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit28.Q net241
+ net229 net230 net154 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit29.Q
+ _0054_ VPWR VGND sg13g2_mux4_1
Xfanout712 net713 net712 VPWR VGND sg13g2_buf_1
Xfanout734 net736 net734 VPWR VGND sg13g2_buf_1
Xfanout789 net106 net789 VPWR VGND sg13g2_buf_1
Xfanout701 net702 net701 VPWR VGND sg13g2_buf_1
Xfanout723 net724 net723 VPWR VGND sg13g2_buf_1
Xfanout745 net747 net745 VPWR VGND sg13g2_buf_1
Xfanout756 net215 net756 VPWR VGND sg13g2_buf_1
Xfanout778 net193 net778 VPWR VGND sg13g2_buf_1
Xfanout767 net204 net767 VPWR VGND sg13g2_buf_1
XFILLER_121_87 VPWR VGND sg13g2_decap_8
XFILLER_53_194 VPWR VGND sg13g2_fill_2
XFILLER_30_51 VPWR VGND sg13g2_fill_2
X_0972_ net804 net711 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
X_1524_ Tile_X0Y1_FrameStrobe[18] net369 VPWR VGND sg13g2_buf_1
Xoutput348 net348 Tile_X0Y0_FrameData_O[28] VPWR VGND sg13g2_buf_1
Xoutput337 net337 Tile_X0Y0_FrameData_O[18] VPWR VGND sg13g2_buf_1
Xoutput359 net359 Tile_X0Y0_FrameData_O[9] VPWR VGND sg13g2_buf_1
Xoutput326 net326 MEN_SRAM VPWR VGND sg13g2_buf_1
Xoutput315 net315 DIN_SRAM28 VPWR VGND sg13g2_buf_1
XFILLER_72_4 VPWR VGND sg13g2_fill_1
Xoutput304 net304 DIN_SRAM18 VPWR VGND sg13g2_buf_1
XFILLER_113_144 VPWR VGND sg13g2_decap_8
X_0337_ VPWR _0040_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG2
+ VGND sg13g2_inv_1
X_1386_ net758 net658 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_27_106 VPWR VGND sg13g2_fill_2
X_1455_ net764 net642 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
X_0406_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit26.Q net157
+ net149 net167 net636 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit27.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb4 VPWR VGND sg13g2_mux4_1
X_1171_ net768 net738 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_2_77 VPWR VGND sg13g2_decap_8
XFILLER_44_8 VPWR VGND sg13g2_fill_1
X_1240_ net197 net714 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
X_0955_ net107 net721 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_82_90 VPWR VGND sg13g2_fill_2
X_0886_ net783 net743 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
X_1507_ net734 net371 VPWR VGND sg13g2_buf_1
XFILLER_63_0 VPWR VGND sg13g2_decap_8
X_1369_ net775 net672 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
X_1438_ net191 net222 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_23_131 VPWR VGND sg13g2_fill_2
XFILLER_11_97 VPWR VGND sg13g2_fill_2
Xinput36 Tile_X0Y0_E1END[2] net36 VPWR VGND sg13g2_buf_1
Xinput25 DOUT_SRAM3 net25 VPWR VGND sg13g2_buf_1
Xinput14 DOUT_SRAM2 net14 VPWR VGND sg13g2_buf_1
X_0740_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG4 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG8
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit2.Q _0184_ VPWR
+ VGND sg13g2_mux2_1
Xinput58 Tile_X0Y0_E6END[2] net58 VPWR VGND sg13g2_buf_1
Xinput69 Tile_X0Y0_EE4END[12] net69 VPWR VGND sg13g2_buf_1
Xinput47 Tile_X0Y0_E2MID[1] net47 VPWR VGND sg13g2_buf_1
X_0671_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit30.Q net245
+ net140 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG9 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG13
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit31.Q Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG2
+ VPWR VGND sg13g2_mux4_1
X_1154_ net102 net644 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
X_1223_ net770 net729 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
X_1085_ net802 net679 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
X_0938_ net94 net720 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
X_0869_ net796 net748 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_78_178 VPWR VGND sg13g2_fill_2
XFILLER_8_76 VPWR VGND sg13g2_fill_1
XFILLER_8_54 VPWR VGND sg13g2_fill_1
X_0723_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit8.Q net186
+ net179 net170 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG6
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit9.Q net322 VPWR
+ VGND sg13g2_mux4_1
X_0585_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit22.Q net35
+ net61 net70 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG1 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit21.Q
+ _0142_ VPWR VGND sg13g2_mux4_1
X_0654_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit10.Q net28
+ net32 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG7 net632 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit11.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG8 VPWR VGND sg13g2_mux4_1
X_1137_ net809 net657 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
X_1206_ net772 net725 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
X_1068_ net804 net679 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_68_37 VPWR VGND sg13g2_fill_1
Xinput226 Tile_X0Y1_N1END[3] net226 VPWR VGND sg13g2_buf_1
Xinput237 Tile_X0Y1_N2MID[2] net237 VPWR VGND sg13g2_buf_1
Xinput248 Tile_X0Y1_N4END[5] net248 VPWR VGND sg13g2_buf_1
Xinput215 Tile_X0Y1_FrameData[3] net215 VPWR VGND sg13g2_buf_1
Xinput204 Tile_X0Y1_FrameData[22] net204 VPWR VGND sg13g2_buf_1
X_0370_ VGND VPWR _0064_ _0065_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit29.Q
+ _0004_ _0066_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit28.Q
+ sg13g2_a221oi_1
XFILLER_3_174 VPWR VGND sg13g2_decap_8
XFILLER_81_118 VPWR VGND sg13g2_decap_4
X_0706_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit6.Q net185
+ net178 net169 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG5
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit7.Q net288 VPWR
+ VGND sg13g2_mux4_1
X_1686_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG3 net540 VPWR
+ VGND sg13g2_buf_1
X_0499_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit10.Q net78
+ net71 net62 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG6 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit11.Q
+ net309 VPWR VGND sg13g2_mux4_1
X_0568_ VGND VPWR _0014_ _0123_ _0127_ _0126_ sg13g2_a21oi_1
XFILLER_57_148 VPWR VGND sg13g2_fill_1
X_0637_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit18.Q net28
+ net6 net637 net635 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit19.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb4 VPWR VGND sg13g2_mux4_1
XFILLER_119_150 VPWR VGND sg13g2_decap_8
XFILLER_70_49 VPWR VGND sg13g2_fill_2
XFILLER_119_87 VPWR VGND sg13g2_decap_8
XFILLER_79_47 VPWR VGND sg13g2_fill_2
XFILLER_63_129 VPWR VGND sg13g2_decap_8
XFILLER_56_181 VPWR VGND sg13g2_fill_1
Xoutput508 net508 Tile_X0Y1_S2BEG[7] VPWR VGND sg13g2_buf_1
Xoutput519 net519 Tile_X0Y1_S4BEG[11] VPWR VGND sg13g2_buf_1
X_1540_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb2 net394 VPWR
+ VGND sg13g2_buf_1
X_0422_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit23.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb7
+ net133 net242 net125 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit22.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG7 VPWR VGND sg13g2_mux4_1
XFILLER_5_99 VPWR VGND sg13g2_fill_1
X_0353_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit28.Q net157
+ net160 net147 net148 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit29.Q
+ _0053_ VPWR VGND sg13g2_mux4_1
XFILLER_62_173 VPWR VGND sg13g2_fill_2
XFILLER_62_140 VPWR VGND sg13g2_fill_1
X_1669_ Tile_X0Y0_S4END[14] net529 VPWR VGND sg13g2_buf_1
Xfanout713 Tile_X0Y1_FrameStrobe[3] net713 VPWR VGND sg13g2_buf_1
Xfanout724 Tile_X0Y1_FrameStrobe[2] net724 VPWR VGND sg13g2_buf_1
Xfanout702 Tile_X0Y1_FrameStrobe[4] net702 VPWR VGND sg13g2_buf_1
Xfanout735 net736 net735 VPWR VGND sg13g2_buf_1
Xfanout746 net747 net746 VPWR VGND sg13g2_buf_1
Xfanout768 net203 net768 VPWR VGND sg13g2_buf_1
Xfanout757 net214 net757 VPWR VGND sg13g2_buf_1
Xfanout779 net192 net779 VPWR VGND sg13g2_buf_1
XFILLER_121_66 VPWR VGND sg13g2_decap_8
XFILLER_81_26 VPWR VGND sg13g2_fill_2
XFILLER_107_131 VPWR VGND sg13g2_fill_2
XFILLER_122_112 VPWR VGND sg13g2_decap_8
XFILLER_44_151 VPWR VGND sg13g2_fill_1
X_0971_ net803 net711 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
X_1523_ Tile_X0Y1_FrameStrobe[17] net368 VPWR VGND sg13g2_buf_1
Xoutput349 net349 Tile_X0Y0_FrameData_O[29] VPWR VGND sg13g2_buf_1
Xoutput338 net338 Tile_X0Y0_FrameData_O[19] VPWR VGND sg13g2_buf_1
Xoutput316 net316 DIN_SRAM29 VPWR VGND sg13g2_buf_1
Xoutput327 net327 REN_SRAM VPWR VGND sg13g2_buf_1
Xoutput305 net305 DIN_SRAM19 VPWR VGND sg13g2_buf_1
X_1454_ net763 net642 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
X_0336_ VPWR _0039_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG1
+ VGND sg13g2_inv_1
X_0405_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit16.Q net239
+ net231 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG4 net130 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit17.Q
+ _0081_ VPWR VGND sg13g2_mux4_1
X_1385_ net757 net658 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_116_88 VPWR VGND sg13g2_decap_8
XFILLER_41_176 VPWR VGND sg13g2_fill_2
XFILLER_41_62 VPWR VGND sg13g2_fill_1
XFILLER_2_56 VPWR VGND sg13g2_decap_8
X_1170_ net767 net738 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
X_0954_ net108 net720 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
X_0885_ net782 net743 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
X_1506_ net746 net360 VPWR VGND sg13g2_buf_1
X_1437_ net192 net651 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
X_1368_ net774 net674 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
X_0319_ VPWR _0022_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit6.Q
+ VGND sg13g2_inv_1
X_1299_ net768 net693 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_23_143 VPWR VGND sg13g2_fill_1
XFILLER_23_176 VPWR VGND sg13g2_fill_2
XFILLER_11_76 VPWR VGND sg13g2_decap_8
XFILLER_11_54 VPWR VGND sg13g2_fill_1
Xinput59 Tile_X0Y0_E6END[3] net59 VPWR VGND sg13g2_buf_1
Xinput48 Tile_X0Y0_E2MID[2] net48 VPWR VGND sg13g2_buf_1
Xinput37 Tile_X0Y0_E1END[3] net37 VPWR VGND sg13g2_buf_1
Xinput15 DOUT_SRAM20 net15 VPWR VGND sg13g2_buf_1
X_0670_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit28.Q net244
+ net139 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG10 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG14
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit29.Q Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG1
+ VPWR VGND sg13g2_mux4_1
Xinput26 DOUT_SRAM30 net26 VPWR VGND sg13g2_buf_1
XFILLER_96_135 VPWR VGND sg13g2_fill_1
X_1153_ net103 net645 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_96_157 VPWR VGND sg13g2_fill_2
X_1084_ net791 net679 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_28_4 VPWR VGND sg13g2_fill_2
X_1222_ net212 net729 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_20_124 VPWR VGND sg13g2_decap_4
X_0937_ net95 net720 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
X_0868_ net795 net744 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
X_0799_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit13.Q VPWR
+ _0237_ VGND net170 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit12.Q
+ sg13g2_o21ai_1
XFILLER_22_64 VPWR VGND sg13g2_fill_1
XFILLER_78_113 VPWR VGND sg13g2_fill_1
XFILLER_22_97 VPWR VGND sg13g2_fill_2
XFILLER_6_172 VPWR VGND sg13g2_decap_4
X_0722_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit6.Q net185
+ net178 net169 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG5
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit7.Q net321 VPWR
+ VGND sg13g2_mux4_1
X_0653_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit22.Q net226
+ net246 _0074_ net141 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit23.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG7 VPWR VGND sg13g2_mux4_1
X_0584_ VGND VPWR _0016_ _0137_ _0141_ _0140_ sg13g2_a21oi_1
XFILLER_33_2 VPWR VGND sg13g2_fill_1
X_1136_ net808 net657 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
X_1067_ net803 net679 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
X_1205_ net771 net726 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_90_108 VPWR VGND sg13g2_decap_8
Xinput238 Tile_X0Y1_N2MID[3] net238 VPWR VGND sg13g2_buf_1
Xinput227 Tile_X0Y1_N2END[0] net227 VPWR VGND sg13g2_buf_1
Xinput249 Tile_X0Y1_N4END[6] net249 VPWR VGND sg13g2_buf_1
Xinput216 Tile_X0Y1_FrameData[4] net216 VPWR VGND sg13g2_buf_1
Xinput205 Tile_X0Y1_FrameData[23] net205 VPWR VGND sg13g2_buf_1
XFILLER_17_97 VPWR VGND sg13g2_fill_1
XFILLER_123_0 VPWR VGND sg13g2_fill_1
XFILLER_3_153 VPWR VGND sg13g2_decap_8
XFILLER_59_190 VPWR VGND sg13g2_fill_2
X_1685_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG2 net539 VPWR
+ VGND sg13g2_buf_1
X_0636_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit16.Q net25
+ net5 net637 net635 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit17.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb3 VPWR VGND sg13g2_mux4_1
X_0705_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit4.Q net184
+ net177 net168 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG4
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit5.Q net287 VPWR
+ VGND sg13g2_mux4_1
X_0567_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit25.Q VPWR
+ _0126_ VGND _0124_ _0125_ sg13g2_o21ai_1
X_0498_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit8.Q net77
+ net70 net61 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG5 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit9.Q
+ net308 VPWR VGND sg13g2_mux4_1
X_1119_ net789 net655 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_80_196 VPWR VGND sg13g2_fill_1
XFILLER_119_55 VPWR VGND sg13g2_decap_8
Xoutput509 net509 Tile_X0Y1_S2BEGb[0] VPWR VGND sg13g2_buf_1
X_1470_ net191 net643 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_10_4 VPWR VGND sg13g2_fill_2
X_0421_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit0.Q net154
+ net146 net162 _0084_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit1.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb7 VPWR VGND sg13g2_mux4_1
X_0352_ _0047_ VPWR _0052_ VGND Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit28.Q
+ _0051_ sg13g2_o21ai_1
X_1668_ Tile_X0Y0_S4END[13] net528 VPWR VGND sg13g2_buf_1
X_1599_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG4 net459 VPWR
+ VGND sg13g2_buf_1
Xfanout747 net748 net747 VPWR VGND sg13g2_buf_1
Xfanout736 net737 net736 VPWR VGND sg13g2_buf_1
Xfanout725 net727 net725 VPWR VGND sg13g2_buf_1
Xfanout714 net715 net714 VPWR VGND sg13g2_buf_1
X_0619_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit2.Q net144
+ net155 net147 _0083_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit3.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG6 VPWR VGND sg13g2_mux4_1
Xfanout758 net213 net758 VPWR VGND sg13g2_buf_1
Xfanout703 net705 net703 VPWR VGND sg13g2_buf_1
Xfanout769 net202 net769 VPWR VGND sg13g2_buf_1
XFILLER_121_45 VPWR VGND sg13g2_decap_8
XFILLER_53_196 VPWR VGND sg13g2_fill_1
XFILLER_122_135 VPWR VGND sg13g2_fill_2
X_0970_ net801 net710 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_113_168 VPWR VGND sg13g2_fill_1
Xoutput328 net328 Tile_X0Y0_FrameData_O[0] VPWR VGND sg13g2_buf_1
Xoutput339 net339 Tile_X0Y0_FrameData_O[1] VPWR VGND sg13g2_buf_1
X_0404_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit11.Q net34
+ net41 net49 net626 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit10.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG4 VPWR VGND sg13g2_mux4_1
X_1522_ Tile_X0Y1_FrameStrobe[16] net367 VPWR VGND sg13g2_buf_1
X_1453_ net762 net642 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
Xoutput306 net306 DIN_SRAM2 VPWR VGND sg13g2_buf_1
Xoutput317 net317 DIN_SRAM3 VPWR VGND sg13g2_buf_1
X_0335_ VPWR _0038_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG0
+ VGND sg13g2_inv_1
X_1384_ net781 net674 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_27_108 VPWR VGND sg13g2_fill_1
XFILLER_50_155 VPWR VGND sg13g2_fill_2
XFILLER_116_67 VPWR VGND sg13g2_decap_8
XFILLER_112_190 VPWR VGND sg13g2_fill_2
XFILLER_92_15 VPWR VGND sg13g2_fill_1
XFILLER_41_199 VPWR VGND sg13g2_fill_2
XFILLER_2_35 VPWR VGND sg13g2_decap_8
XFILLER_17_141 VPWR VGND sg13g2_decap_4
X_0953_ net109 net720 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
X_0884_ net812 net745 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_101_138 VPWR VGND sg13g2_fill_2
X_1505_ net789 net352 VPWR VGND sg13g2_buf_1
X_1367_ net773 net674 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
X_1436_ net193 net651 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
X_0318_ VPWR _0021_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit5.Q
+ VGND sg13g2_inv_1
X_1298_ net767 net694 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_23_199 VPWR VGND sg13g2_fill_2
Xinput49 Tile_X0Y0_E2MID[3] net49 VPWR VGND sg13g2_buf_1
Xinput38 Tile_X0Y0_E2END[0] net38 VPWR VGND sg13g2_buf_1
Xinput16 DOUT_SRAM21 net16 VPWR VGND sg13g2_buf_1
Xinput27 DOUT_SRAM31 net27 VPWR VGND sg13g2_buf_1
X_1221_ net215 net731 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
X_1152_ net105 net644 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
X_1083_ net788 net679 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
X_0936_ net799 net723 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
X_0867_ net794 net747 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
X_0798_ VGND VPWR _0229_ _0231_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S4BEG1
+ _0236_ sg13g2_a21oi_1
XFILLER_87_158 VPWR VGND sg13g2_fill_2
X_1419_ net211 net649 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_63_50 VPWR VGND sg13g2_fill_1
X_0583_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit23.Q VPWR
+ _0140_ VGND _0138_ _0139_ sg13g2_o21ai_1
XFILLER_6_195 VPWR VGND sg13g2_fill_2
X_0652_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit8.Q net31
+ net5 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG8 net640 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit9.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG7 VPWR VGND sg13g2_mux4_1
X_0721_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit4.Q net184
+ net177 net168 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG4
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit5.Q net320 VPWR
+ VGND sg13g2_mux4_1
XFILLER_111_200 VPWR VGND sg13g2_fill_1
XFILLER_84_106 VPWR VGND sg13g2_decap_4
X_1204_ net769 net725 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
X_1135_ net807 net657 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
X_1066_ net801 net676 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
X_0919_ net784 net732 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_102_200 VPWR VGND sg13g2_fill_1
Xinput217 Tile_X0Y1_FrameData[5] net217 VPWR VGND sg13g2_buf_1
Xinput206 Tile_X0Y1_FrameData[24] net206 VPWR VGND sg13g2_buf_1
XFILLER_75_128 VPWR VGND sg13g2_fill_1
Xinput239 Tile_X0Y1_N2MID[4] net239 VPWR VGND sg13g2_buf_1
Xinput228 Tile_X0Y1_N2END[1] net228 VPWR VGND sg13g2_buf_1
XFILLER_3_132 VPWR VGND sg13g2_decap_8
XFILLER_33_97 VPWR VGND sg13g2_fill_1
XFILLER_58_72 VPWR VGND sg13g2_fill_2
XFILLER_74_82 VPWR VGND sg13g2_decap_8
X_0566_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit24.Q VPWR
+ _0125_ VGND Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit23.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG15 sg13g2_o21ai_1
X_0704_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit2.Q net183
+ net176 net167 _0158_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit3.Q
+ net284 VPWR VGND sg13g2_mux4_1
X_1684_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG1 net538 VPWR
+ VGND sg13g2_buf_1
X_0635_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit14.Q net14
+ net4 net638 net634 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit15.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb2 VPWR VGND sg13g2_mux4_1
X_0497_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit6.Q net76
+ net69 net60 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG4 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit7.Q
+ net307 VPWR VGND sg13g2_mux4_1
X_1118_ net813 net666 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
X_1049_ net786 net686 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_119_185 VPWR VGND sg13g2_decap_4
XFILLER_119_34 VPWR VGND sg13g2_decap_8
XFILLER_0_168 VPWR VGND sg13g2_fill_1
XFILLER_28_53 VPWR VGND sg13g2_fill_2
X_0420_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit22.Q net242
+ net234 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG7 net133 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit23.Q
+ _0084_ VPWR VGND sg13g2_mux4_1
XFILLER_60_95 VPWR VGND sg13g2_fill_1
XFILLER_5_24 VPWR VGND sg13g2_decap_8
X_0351_ _0050_ VPWR _0051_ VGND Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit29.Q
+ _0049_ sg13g2_o21ai_1
X_1667_ Tile_X0Y0_S4END[12] net527 VPWR VGND sg13g2_buf_1
X_0549_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG1 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit17.Q
+ _0110_ VPWR VGND sg13g2_nor2b_1
Xfanout737 Tile_X0Y1_FrameStrobe[1] net737 VPWR VGND sg13g2_buf_1
X_1598_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG3 net458 VPWR
+ VGND sg13g2_buf_1
Xfanout748 net749 net748 VPWR VGND sg13g2_buf_1
Xfanout759 net212 net759 VPWR VGND sg13g2_buf_1
Xfanout726 net727 net726 VPWR VGND sg13g2_buf_1
X_0618_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit0.Q net143
+ net156 net148 _0082_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit1.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG5 VPWR VGND sg13g2_mux4_1
Xfanout715 net716 net715 VPWR VGND sg13g2_buf_1
Xfanout704 net705 net704 VPWR VGND sg13g2_buf_1
XFILLER_121_24 VPWR VGND sg13g2_decap_8
XFILLER_65_18 VPWR VGND sg13g2_decap_8
XFILLER_107_133 VPWR VGND sg13g2_fill_1
Xoutput307 net307 DIN_SRAM20 VPWR VGND sg13g2_buf_1
X_1521_ Tile_X0Y1_FrameStrobe[15] net366 VPWR VGND sg13g2_buf_1
Xoutput329 net329 Tile_X0Y0_FrameData_O[10] VPWR VGND sg13g2_buf_1
X_0403_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit4.Q net50
+ net42 net60 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG3 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit5.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG3 VPWR VGND sg13g2_mux4_1
Xoutput318 net318 DIN_SRAM30 VPWR VGND sg13g2_buf_1
X_1383_ net770 net674 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
X_1452_ net761 net641 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
X_0334_ VPWR _0037_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit5.Q
+ VGND sg13g2_inv_1
X_1719_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG8 net579 VPWR
+ VGND sg13g2_buf_1
X_0952_ net785 net723 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
X_1504_ net790 net351 VPWR VGND sg13g2_buf_1
X_0883_ net811 net745 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
X_1366_ net772 net673 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
X_0317_ VPWR _0020_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit3.Q
+ VGND sg13g2_inv_1
X_1435_ net777 net651 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_102_26 VPWR VGND sg13g2_fill_2
X_1297_ net766 net695 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_14_101 VPWR VGND sg13g2_decap_8
XFILLER_52_63 VPWR VGND sg13g2_fill_2
Xinput39 Tile_X0Y0_E2END[1] net39 VPWR VGND sg13g2_buf_1
Xinput28 DOUT_SRAM4 net28 VPWR VGND sg13g2_buf_1
Xinput17 DOUT_SRAM22 net17 VPWR VGND sg13g2_buf_1
X_1151_ net106 net644 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_96_159 VPWR VGND sg13g2_fill_1
XFILLER_77_71 VPWR VGND sg13g2_decap_8
XFILLER_28_6 VPWR VGND sg13g2_fill_1
X_1220_ net216 net729 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
X_1082_ net787 net677 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
X_0866_ net793 net746 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
X_0935_ net798 net723 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_61_0 VPWR VGND sg13g2_decap_8
X_0797_ VGND VPWR _0030_ _0234_ _0236_ _0235_ sg13g2_a21oi_1
XFILLER_113_58 VPWR VGND sg13g2_fill_1
X_1349_ net756 net680 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_3_90 VPWR VGND sg13g2_decap_8
X_1418_ net758 net647 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_7_119 VPWR VGND sg13g2_fill_2
Xoutput490 net490 Tile_X0Y1_FrameData_O[3] VPWR VGND sg13g2_buf_1
X_0720_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit2.Q net183
+ net176 net167 _0158_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit3.Q
+ net317 VPWR VGND sg13g2_mux4_1
X_0582_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit22.Q VPWR
+ _0139_ VGND Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit21.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG13 sg13g2_o21ai_1
XFILLER_69_126 VPWR VGND sg13g2_fill_1
X_0651_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit24.Q net223
+ net243 _0088_ net138 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit25.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG8 VPWR VGND sg13g2_mux4_1
X_1134_ net806 net657 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
X_1203_ net768 net725 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
X_1065_ net800 net676 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
X_0918_ net783 net731 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
X_0849_ _0284_ net157 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit4.Q
+ VPWR VGND sg13g2_nand2b_1
XFILLER_75_118 VPWR VGND sg13g2_fill_2
Xinput229 Tile_X0Y1_N2END[2] net229 VPWR VGND sg13g2_buf_1
Xinput218 Tile_X0Y1_FrameData[6] net218 VPWR VGND sg13g2_buf_1
Xinput207 Tile_X0Y1_FrameData[25] net207 VPWR VGND sg13g2_buf_1
XFILLER_84_28 VPWR VGND sg13g2_fill_2
XFILLER_83_195 VPWR VGND sg13g2_fill_2
XFILLER_59_192 VPWR VGND sg13g2_fill_1
XFILLER_3_188 VPWR VGND sg13g2_decap_4
X_1683_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG0 net537 VPWR
+ VGND sg13g2_buf_1
X_0703_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit0.Q net182
+ net175 net166 _0159_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit1.Q
+ net273 VPWR VGND sg13g2_mux4_1
X_0496_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit4.Q net75
+ net68 net59 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG3 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit5.Q
+ net305 VPWR VGND sg13g2_mux4_1
X_0565_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG3 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit23.Q
+ _0124_ VPWR VGND sg13g2_nor2b_1
X_0634_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit12.Q net3
+ net33 net639 net633 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit13.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb1 VPWR VGND sg13g2_mux4_1
X_1117_ net802 net666 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
X_1048_ net785 net685 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_119_164 VPWR VGND sg13g2_decap_8
XFILLER_100_81 VPWR VGND sg13g2_fill_1
XFILLER_69_83 VPWR VGND sg13g2_fill_1
XFILLER_69_72 VPWR VGND sg13g2_decap_8
X_0350_ net151 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit29.Q
+ _0050_ VPWR VGND Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit30.Q
+ sg13g2_nand3b_1
XFILLER_10_6 VPWR VGND sg13g2_fill_1
XFILLER_39_129 VPWR VGND sg13g2_fill_2
XFILLER_47_173 VPWR VGND sg13g2_fill_1
X_1666_ Tile_X0Y0_S4END[11] net526 VPWR VGND sg13g2_buf_1
X_0548_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG5 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG9
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit17.Q _0109_ VPWR
+ VGND sg13g2_mux2_1
X_1597_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG2 net457 VPWR
+ VGND sg13g2_buf_1
X_0479_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit8.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END0
+ net247 net114 net134 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit9.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG0 VPWR VGND sg13g2_mux4_1
Xfanout749 Tile_X0Y1_FrameStrobe[0] net749 VPWR VGND sg13g2_buf_1
Xfanout738 net749 net738 VPWR VGND sg13g2_buf_1
Xfanout716 net719 net716 VPWR VGND sg13g2_buf_1
Xfanout727 net737 net727 VPWR VGND sg13g2_buf_1
X_0617_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit31.Q net142
+ net149 net157 net635 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit30.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG4 VPWR VGND sg13g2_mux4_1
Xfanout705 net708 net705 VPWR VGND sg13g2_buf_1
XFILLER_107_101 VPWR VGND sg13g2_decap_4
XFILLER_39_75 VPWR VGND sg13g2_fill_1
XFILLER_55_30 VPWR VGND sg13g2_fill_2
XFILLER_71_73 VPWR VGND sg13g2_fill_1
X_1520_ Tile_X0Y1_FrameStrobe[14] net365 VPWR VGND sg13g2_buf_1
Xoutput319 net319 DIN_SRAM31 VPWR VGND sg13g2_buf_1
Xoutput308 net308 DIN_SRAM21 VPWR VGND sg13g2_buf_1
XFILLER_71_95 VPWR VGND sg13g2_fill_2
XFILLER_113_137 VPWR VGND sg13g2_decap_8
X_0402_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit14.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb3
+ net238 net129 net121 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit15.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG3 VPWR VGND sg13g2_mux4_1
X_0333_ VPWR _0036_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit3.Q
+ VGND sg13g2_inv_1
X_1382_ net759 net670 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
X_1451_ net760 net641 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
X_1718_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG7 net578 VPWR
+ VGND sg13g2_buf_1
X_1649_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG2 net503 VPWR
+ VGND sg13g2_buf_1
XFILLER_112_192 VPWR VGND sg13g2_fill_1
XFILLER_17_176 VPWR VGND sg13g2_fill_2
X_0951_ net784 net723 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
X_0882_ net810 net745 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
X_1503_ net792 net349 VPWR VGND sg13g2_buf_1
X_1365_ net771 net673 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
X_1434_ net776 net649 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
X_0316_ VPWR _0019_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit2.Q
+ VGND sg13g2_inv_1
X_1296_ net206 net696 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_23_124 VPWR VGND sg13g2_decap_8
Xinput18 DOUT_SRAM23 net18 VPWR VGND sg13g2_buf_1
Xinput29 DOUT_SRAM5 net29 VPWR VGND sg13g2_buf_1
X_1150_ net82 net654 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
X_1081_ net786 net675 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_20_105 VPWR VGND sg13g2_fill_2
X_0865_ net792 net745 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
X_0934_ net797 net723 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
X_0796_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit11.Q VPWR
+ _0235_ VGND _0232_ _0233_ sg13g2_o21ai_1
X_1417_ net757 net647 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
X_1348_ net755 net680 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
X_1279_ net750 net707 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_22_45 VPWR VGND sg13g2_fill_2
Xoutput480 net480 Tile_X0Y1_FrameData_O[23] VPWR VGND sg13g2_buf_1
Xoutput491 net491 Tile_X0Y1_FrameData_O[4] VPWR VGND sg13g2_buf_1
XFILLER_63_85 VPWR VGND sg13g2_fill_2
XFILLER_47_75 VPWR VGND sg13g2_fill_2
XFILLER_8_36 VPWR VGND sg13g2_fill_1
XFILLER_6_120 VPWR VGND sg13g2_decap_4
XFILLER_88_93 VPWR VGND sg13g2_fill_2
X_0581_ net625 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit21.Q
+ _0138_ VPWR VGND sg13g2_nor2b_1
X_0650_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit6.Q net30
+ net4 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG9 net639 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit7.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG6 VPWR VGND sg13g2_mux4_1
X_1133_ net805 net653 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
X_1064_ net799 net675 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
X_1202_ net767 net728 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_92_196 VPWR VGND sg13g2_fill_1
X_0917_ net782 net731 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
X_0779_ _0218_ VPWR _0219_ VGND _0027_ _0161_ sg13g2_o21ai_1
X_0848_ _0283_ _0037_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit6.Q
+ VPWR VGND sg13g2_nand2_1
XFILLER_75_108 VPWR VGND sg13g2_fill_2
Xinput219 Tile_X0Y1_FrameData[7] net219 VPWR VGND sg13g2_buf_1
Xinput208 Tile_X0Y1_FrameData[26] net208 VPWR VGND sg13g2_buf_1
XFILLER_3_167 VPWR VGND sg13g2_decap_8
XFILLER_59_171 VPWR VGND sg13g2_fill_2
X_0633_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit10.Q net2
+ net32 net640 net632 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit11.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb0 VPWR VGND sg13g2_mux4_1
X_1682_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W1BEG3 net536 VPWR
+ VGND sg13g2_buf_1
X_0702_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit30.Q net181
+ net189 net165 _0160_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit31.Q
+ net262 VPWR VGND sg13g2_mux4_1
X_0495_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit2.Q net74
+ net67 net58 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG2 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit3.Q
+ net304 VPWR VGND sg13g2_mux4_1
X_0564_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG7 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG11
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit23.Q _0123_ VPWR
+ VGND sg13g2_mux2_1
XFILLER_57_108 VPWR VGND sg13g2_fill_1
X_1116_ net791 net664 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
X_1047_ net784 net686 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_80_111 VPWR VGND sg13g2_fill_2
XFILLER_17_0 VPWR VGND sg13g2_fill_2
XFILLER_119_143 VPWR VGND sg13g2_decap_8
XFILLER_95_39 VPWR VGND sg13g2_fill_2
XFILLER_28_55 VPWR VGND sg13g2_fill_1
XFILLER_60_42 VPWR VGND sg13g2_decap_8
XFILLER_62_166 VPWR VGND sg13g2_decap_8
X_1665_ Tile_X0Y0_S4END[10] net525 VPWR VGND sg13g2_buf_1
XFILLER_116_102 VPWR VGND sg13g2_decap_4
X_1596_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG1 net456 VPWR
+ VGND sg13g2_buf_1
X_0616_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit29.Q net158
+ net164 net150 _0080_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit28.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG3 VPWR VGND sg13g2_mux4_1
Xfanout706 net708 net706 VPWR VGND sg13g2_buf_1
X_0547_ _0106_ _0108_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N4BEG0
+ VPWR VGND sg13g2_nor2_1
X_0478_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit2.Q net12
+ net26 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG1 net630 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit3.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG14 VPWR VGND sg13g2_mux4_1
Xfanout739 net749 net739 VPWR VGND sg13g2_buf_1
Xfanout728 net730 net728 VPWR VGND sg13g2_buf_1
Xfanout717 net718 net717 VPWR VGND sg13g2_buf_1
XFILLER_121_59 VPWR VGND sg13g2_decap_8
XFILLER_122_149 VPWR VGND sg13g2_decap_8
XFILLER_122_105 VPWR VGND sg13g2_decap_8
XFILLER_55_53 VPWR VGND sg13g2_fill_1
XFILLER_55_75 VPWR VGND sg13g2_decap_4
XFILLER_55_97 VPWR VGND sg13g2_fill_2
Xoutput309 net309 DIN_SRAM22 VPWR VGND sg13g2_buf_1
XFILLER_65_8 VPWR VGND sg13g2_decap_4
X_1450_ net758 net641 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_121_171 VPWR VGND sg13g2_fill_2
X_1381_ net756 net670 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
X_0401_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit25.Q net158
+ net168 net150 _0080_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit24.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb3 VPWR VGND sg13g2_mux4_1
X_0332_ VPWR _0035_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit0.Q
+ VGND sg13g2_inv_1
XFILLER_84_0 VPWR VGND sg13g2_fill_2
XFILLER_104_116 VPWR VGND sg13g2_fill_1
X_1579_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb4 net433 VPWR
+ VGND sg13g2_buf_1
X_1717_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG6 net577 VPWR
+ VGND sg13g2_buf_1
X_1648_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG1 net502 VPWR
+ VGND sg13g2_buf_1
XFILLER_25_45 VPWR VGND sg13g2_fill_1
XFILLER_41_77 VPWR VGND sg13g2_fill_1
XFILLER_103_160 VPWR VGND sg13g2_fill_1
XFILLER_2_49 VPWR VGND sg13g2_decap_8
XFILLER_17_199 VPWR VGND sg13g2_fill_2
X_0950_ net783 net719 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
X_0881_ net809 net745 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
X_1502_ net793 net348 VPWR VGND sg13g2_buf_1
XFILLER_99_125 VPWR VGND sg13g2_fill_2
X_1433_ net775 net649 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
X_0315_ VPWR _0018_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit28.Q
+ VGND sg13g2_inv_1
X_1364_ net769 net669 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
X_1295_ net207 net696 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_100_141 VPWR VGND sg13g2_fill_2
XFILLER_36_55 VPWR VGND sg13g2_fill_2
Xinput19 DOUT_SRAM24 net19 VPWR VGND sg13g2_buf_1
X_1080_ net785 net676 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_114_200 VPWR VGND sg13g2_fill_1
X_0864_ net790 net745 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
X_0933_ net796 net723 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
X_0795_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG5 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG9
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit9.Q _0234_ VPWR
+ VGND sg13g2_mux2_1
X_1347_ net754 net680 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
X_1416_ net781 net659 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
X_1278_ net191 net705 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
Xoutput470 net470 Tile_X0Y1_FrameData_O[14] VPWR VGND sg13g2_buf_1
Xoutput481 net481 Tile_X0Y1_FrameData_O[24] VPWR VGND sg13g2_buf_1
Xoutput492 net492 Tile_X0Y1_FrameData_O[5] VPWR VGND sg13g2_buf_1
XFILLER_93_109 VPWR VGND sg13g2_fill_2
XFILLER_78_139 VPWR VGND sg13g2_fill_1
XFILLER_10_194 VPWR VGND sg13g2_fill_2
XFILLER_6_176 VPWR VGND sg13g2_fill_2
X_0580_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG5 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG9
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit21.Q _0137_ VPWR
+ VGND sg13g2_mux2_1
X_1201_ net766 net728 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
X_1132_ net91 net653 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_92_164 VPWR VGND sg13g2_fill_2
X_1063_ net798 net675 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_19_4 VPWR VGND sg13g2_fill_1
X_0916_ net812 net732 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
X_0778_ VPWR _0218_ _0217_ VGND sg13g2_inv_1
X_0847_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit5.Q Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit6.Q
+ _0281_ _0282_ VPWR VGND sg13g2_nor3_1
Xinput209 Tile_X0Y1_FrameData[27] net209 VPWR VGND sg13g2_buf_1
XFILLER_3_146 VPWR VGND sg13g2_decap_8
X_0563_ _0120_ _0122_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N4BEG2
+ VPWR VGND sg13g2_nor2_1
X_1681_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W1BEG2 net535 VPWR
+ VGND sg13g2_buf_1
X_0632_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit8.Q net31
+ net9 net640 net632 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit9.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG7 VPWR VGND sg13g2_mux4_1
X_0701_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit28.Q net174
+ net188 net162 _0161_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit29.Q
+ net261 VPWR VGND sg13g2_mux4_1
X_0494_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit0.Q net73
+ net81 net57 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG1 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit1.Q
+ net303 VPWR VGND sg13g2_mux4_1
X_1115_ net788 net665 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
X_1046_ net112 net688 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_80_178 VPWR VGND sg13g2_fill_1
XFILLER_119_122 VPWR VGND sg13g2_decap_8
XFILLER_119_48 VPWR VGND sg13g2_decap_8
XFILLER_86_4 VPWR VGND sg13g2_fill_1
X_1595_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG0 net449 VPWR
+ VGND sg13g2_buf_1
X_0546_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit16.Q _0107_
+ _0108_ VPWR VGND sg13g2_nor2_1
X_1664_ Tile_X0Y0_S4END[9] net524 VPWR VGND sg13g2_buf_1
Xfanout729 net730 net729 VPWR VGND sg13g2_buf_1
Xfanout707 net708 net707 VPWR VGND sg13g2_buf_1
X_0615_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit27.Q net159
+ net163 net151 _0079_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit26.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG2 VPWR VGND sg13g2_mux4_1
Xfanout718 net719 net718 VPWR VGND sg13g2_buf_1
X_0477_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit10.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END1
+ net248 net115 net135 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit11.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG1 VPWR VGND sg13g2_mux4_1
XFILLER_53_101 VPWR VGND sg13g2_decap_4
XFILLER_121_38 VPWR VGND sg13g2_decap_8
X_1029_ net796 net688 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_115_180 VPWR VGND sg13g2_fill_1
XFILLER_29_131 VPWR VGND sg13g2_fill_1
XFILLER_55_32 VPWR VGND sg13g2_fill_1
XFILLER_71_97 VPWR VGND sg13g2_fill_1
XFILLER_71_53 VPWR VGND sg13g2_fill_2
XFILLER_58_8 VPWR VGND sg13g2_decap_8
X_1380_ net755 net669 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
X_0400_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit15.Q net238
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG3 net230 net129 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit14.Q
+ _0080_ VPWR VGND sg13g2_mux4_1
XFILLER_121_150 VPWR VGND sg13g2_decap_8
X_0331_ VPWR _0034_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit16.Q
+ VGND sg13g2_inv_1
XFILLER_50_104 VPWR VGND sg13g2_decap_8
X_1716_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG5 net576 VPWR
+ VGND sg13g2_buf_1
X_0529_ _0095_ net39 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit1.Q
+ VPWR VGND sg13g2_nand2b_1
X_1578_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb3 net432 VPWR
+ VGND sg13g2_buf_1
X_1647_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG0 net501 VPWR
+ VGND sg13g2_buf_1
XFILLER_1_200 VPWR VGND sg13g2_fill_1
XFILLER_66_86 VPWR VGND sg13g2_fill_1
XFILLER_66_42 VPWR VGND sg13g2_decap_4
XFILLER_2_28 VPWR VGND sg13g2_decap_8
XFILLER_17_145 VPWR VGND sg13g2_fill_2
X_0880_ net87 net744 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
X_1501_ net794 net347 VPWR VGND sg13g2_buf_1
X_1363_ net768 net669 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
X_1432_ net774 net648 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
X_0314_ VPWR _0017_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit25.Q
+ VGND sg13g2_inv_1
X_1294_ net763 net694 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_11_15 VPWR VGND sg13g2_fill_1
XFILLER_36_12 VPWR VGND sg13g2_fill_2
XFILLER_36_78 VPWR VGND sg13g2_fill_2
XFILLER_117_81 VPWR VGND sg13g2_decap_8
XFILLER_93_51 VPWR VGND sg13g2_fill_1
X_0932_ net100 net722 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
X_0863_ net106 net745 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
X_0794_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit10.Q VPWR
+ _0233_ VGND Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit9.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG13 sg13g2_o21ai_1
X_1346_ net753 net682 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
X_1415_ net770 net660 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
X_1277_ net192 net704 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
Xoutput482 net482 Tile_X0Y1_FrameData_O[25] VPWR VGND sg13g2_buf_1
Xoutput471 net471 Tile_X0Y1_FrameData_O[15] VPWR VGND sg13g2_buf_1
Xoutput493 net493 Tile_X0Y1_FrameData_O[6] VPWR VGND sg13g2_buf_1
Xoutput460 net460 Tile_X0Y0_WW4BEG[5] VPWR VGND sg13g2_buf_1
XFILLER_47_77 VPWR VGND sg13g2_fill_1
XFILLER_88_95 VPWR VGND sg13g2_fill_1
X_1200_ net765 net727 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
X_1131_ net803 net653 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
X_1062_ net797 net675 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
X_0915_ net811 net732 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
X_0777_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit7.Q VPWR
+ _0217_ VGND net168 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit6.Q
+ sg13g2_o21ai_1
X_0846_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit4.Q net241
+ _0281_ VPWR VGND sg13g2_nor2b_1
X_1329_ net766 net683 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_3_125 VPWR VGND sg13g2_decap_8
Xoutput290 net290 BM_SRAM7 VPWR VGND sg13g2_buf_1
XFILLER_74_198 VPWR VGND sg13g2_fill_2
XFILLER_74_20 VPWR VGND sg13g2_fill_2
XFILLER_90_85 VPWR VGND sg13g2_fill_2
X_0700_ _0174_ VPWR net255 VGND Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit27.Q
+ _0176_ sg13g2_o21ai_1
X_0562_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit22.Q _0121_
+ _0122_ VPWR VGND sg13g2_nor2_1
XFILLER_99_50 VPWR VGND sg13g2_fill_1
X_0631_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit6.Q net30
+ net8 net639 net633 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit7.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG6 VPWR VGND sg13g2_mux4_1
X_1680_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W1BEG1 net534 VPWR
+ VGND sg13g2_buf_1
X_1114_ net787 net666 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
X_0493_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit30.Q net66
+ net80 net54 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit31.Q
+ net302 VPWR VGND sg13g2_mux4_1
XFILLER_65_143 VPWR VGND sg13g2_decap_8
XFILLER_31_4 VPWR VGND sg13g2_fill_2
X_1045_ net113 net688 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_119_178 VPWR VGND sg13g2_decap_8
XFILLER_119_101 VPWR VGND sg13g2_decap_8
XFILLER_119_27 VPWR VGND sg13g2_decap_8
X_0829_ VGND VPWR net160 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit0.Q
+ _0265_ _0258_ sg13g2_a21oi_1
XFILLER_107_0 VPWR VGND sg13g2_fill_2
XFILLER_60_99 VPWR VGND sg13g2_fill_1
X_1663_ Tile_X0Y0_S4END[8] net517 VPWR VGND sg13g2_buf_1
XFILLER_79_4 VPWR VGND sg13g2_fill_1
X_0476_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit0.Q net11
+ net24 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG2 net629 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit1.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG13 VPWR VGND sg13g2_mux4_1
X_0545_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit14.Q net34
+ net66 net64 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit15.Q
+ _0107_ VPWR VGND sg13g2_mux4_1
X_1594_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG11 net439 VPWR
+ VGND sg13g2_buf_1
Xfanout708 Tile_X0Y1_FrameStrobe[3] net708 VPWR VGND sg13g2_buf_1
Xfanout719 net724 net719 VPWR VGND sg13g2_buf_1
X_0614_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit24.Q net160
+ net152 net173 _0078_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit25.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG1 VPWR VGND sg13g2_mux4_1
X_1028_ net795 net687 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_14_37 VPWR VGND sg13g2_fill_1
XFILLER_107_126 VPWR VGND sg13g2_fill_1
XFILLER_39_56 VPWR VGND sg13g2_fill_2
XFILLER_111_61 VPWR VGND sg13g2_fill_1
XFILLER_111_50 VPWR VGND sg13g2_fill_1
XFILLER_55_99 VPWR VGND sg13g2_fill_1
X_0330_ VPWR _0033_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit15.Q
+ VGND sg13g2_inv_1
XFILLER_35_135 VPWR VGND sg13g2_fill_2
XFILLER_84_2 VPWR VGND sg13g2_fill_1
X_1646_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S1BEG3 net500 VPWR
+ VGND sg13g2_buf_1
X_1715_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG4 net575 VPWR
+ VGND sg13g2_buf_1
X_0459_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit28.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END2
+ net249 net116 net136 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit29.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG10 VPWR VGND sg13g2_mux4_1
X_0528_ net47 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit0.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit1.Q _0094_ VPWR
+ VGND sg13g2_nor3_1
X_1577_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb2 net431 VPWR
+ VGND sg13g2_buf_1
XFILLER_25_25 VPWR VGND sg13g2_fill_2
XFILLER_106_72 VPWR VGND sg13g2_fill_1
XFILLER_15_80 VPWR VGND sg13g2_decap_8
XFILLER_32_138 VPWR VGND sg13g2_fill_2
XFILLER_40_171 VPWR VGND sg13g2_fill_2
X_1500_ net795 net346 VPWR VGND sg13g2_buf_1
XFILLER_63_7 VPWR VGND sg13g2_fill_1
X_0313_ VPWR _0016_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit22.Q
+ VGND sg13g2_inv_1
X_1362_ net767 net671 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
X_1431_ net773 net648 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
X_1293_ net762 net694 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
Xinput190 Tile_X0Y1_FrameData[0] net190 VPWR VGND sg13g2_buf_1
XFILLER_23_149 VPWR VGND sg13g2_fill_2
X_1629_ net772 net474 VPWR VGND sg13g2_buf_1
XFILLER_100_143 VPWR VGND sg13g2_fill_1
XFILLER_52_34 VPWR VGND sg13g2_fill_1
XFILLER_22_171 VPWR VGND sg13g2_fill_1
XFILLER_117_60 VPWR VGND sg13g2_decap_8
X_0931_ net101 net722 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
X_0862_ _0296_ VPWR net581 VGND Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit7.Q
+ _0287_ sg13g2_o21ai_1
X_0793_ _0029_ net634 _0232_ VPWR VGND sg13g2_nor2_1
X_1345_ net752 net682 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_3_83 VPWR VGND sg13g2_decap_8
X_1414_ net759 net659 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
X_1276_ net778 net705 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
Xoutput483 net483 Tile_X0Y1_FrameData_O[26] VPWR VGND sg13g2_buf_1
Xoutput494 net494 Tile_X0Y1_FrameData_O[7] VPWR VGND sg13g2_buf_1
Xoutput472 net472 Tile_X0Y1_FrameData_O[16] VPWR VGND sg13g2_buf_1
Xoutput450 net450 Tile_X0Y0_WW4BEG[10] VPWR VGND sg13g2_buf_1
Xoutput461 net461 Tile_X0Y0_WW4BEG[6] VPWR VGND sg13g2_buf_1
XFILLER_10_141 VPWR VGND sg13g2_fill_2
XFILLER_10_196 VPWR VGND sg13g2_fill_1
X_1130_ net801 net655 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_92_166 VPWR VGND sg13g2_fill_1
X_1061_ net796 net675 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
X_0914_ net810 net735 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
X_0845_ _0280_ net229 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit4.Q
+ VPWR VGND sg13g2_nand2_1
X_0776_ VGND VPWR _0209_ _0211_ Tile_X0Y0_IHP_SRAM_top.N4BEG_outbuf_11.A _0216_ sg13g2_a21oi_1
XFILLER_83_177 VPWR VGND sg13g2_fill_1
X_1328_ net765 net681 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
X_1259_ net760 net706 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_58_22 VPWR VGND sg13g2_decap_4
Xoutput291 net291 BM_SRAM8 VPWR VGND sg13g2_buf_1
Xoutput280 net280 BM_SRAM26 VPWR VGND sg13g2_buf_1
XFILLER_90_20 VPWR VGND sg13g2_fill_2
X_0561_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit21.Q net36
+ net55 net74 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG2 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit20.Q
+ _0121_ VPWR VGND sg13g2_mux4_1
X_0492_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit29.Q net13
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG4 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG0
+ net623 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit28.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG11
+ VPWR VGND sg13g2_mux4_1
X_0630_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit4.Q net29
+ net7 net638 net634 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit5.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG5 VPWR VGND sg13g2_mux4_1
X_1113_ net786 net666 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
X_1044_ net812 net687 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_65_188 VPWR VGND sg13g2_fill_1
XFILLER_119_157 VPWR VGND sg13g2_decap_8
X_0759_ VGND VPWR _0024_ _0200_ _0201_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit10.Q
+ sg13g2_a21oi_1
X_0828_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit2.Q _0262_
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit1.Q _0264_ VPWR
+ VGND _0263_ sg13g2_nand4_1
XFILLER_56_199 VPWR VGND sg13g2_fill_2
XFILLER_62_136 VPWR VGND sg13g2_decap_4
X_1662_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG7 net516 VPWR
+ VGND sg13g2_buf_1
X_0613_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit22.Q net161
+ net153 net172 _0043_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit23.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG0 VPWR VGND sg13g2_mux4_1
X_0475_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit12.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END2
+ net249 net116 net136 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit13.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG2 VPWR VGND sg13g2_mux4_1
X_1593_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG10 net438 VPWR
+ VGND sg13g2_buf_1
X_0544_ VGND VPWR _0011_ _0102_ _0106_ _0105_ sg13g2_a21oi_1
Xfanout709 net713 net709 VPWR VGND sg13g2_buf_1
X_1027_ net794 net687 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_38_122 VPWR VGND sg13g2_fill_1
XFILLER_100_8 VPWR VGND sg13g2_fill_2
XFILLER_71_55 VPWR VGND sg13g2_fill_1
X_1576_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb1 net430 VPWR
+ VGND sg13g2_buf_1
XFILLER_6_72 VPWR VGND sg13g2_fill_2
X_1714_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG3 net574 VPWR
+ VGND sg13g2_buf_1
X_1645_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S1BEG2 net499 VPWR
+ VGND sg13g2_buf_1
X_0389_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit4.Q net52
+ net44 net65 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG1 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit5.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG1 VPWR VGND sg13g2_mux4_1
X_0527_ VGND VPWR Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit30.Q
+ _0092_ _0093_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit31.Q
+ net256 _0038_ sg13g2_a221oi_1
X_0458_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit14.Q net15
+ net19 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG11 net628
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit15.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG4
+ VPWR VGND sg13g2_mux4_1
XFILLER_99_106 VPWR VGND sg13g2_fill_2
X_1430_ net199 net650 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
X_0312_ VPWR _0015_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit19.Q
+ VGND sg13g2_inv_1
X_1361_ net766 net671 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
Xinput180 Tile_X0Y1_EE4END[15] net180 VPWR VGND sg13g2_buf_1
X_1292_ net210 net694 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_23_117 VPWR VGND sg13g2_decap_8
Xinput191 Tile_X0Y1_FrameData[10] net191 VPWR VGND sg13g2_buf_1
XFILLER_82_0 VPWR VGND sg13g2_fill_2
X_1559_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N4BEG1 net404 VPWR
+ VGND sg13g2_buf_1
X_1628_ net198 net473 VPWR VGND sg13g2_buf_1
XFILLER_77_65 VPWR VGND sg13g2_fill_2
X_0930_ net793 net720 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
X_0792_ VGND VPWR _0030_ _0230_ _0231_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit11.Q
+ sg13g2_a21oi_1
X_0861_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit7.Q VPWR
+ _0296_ VGND _0291_ _0295_ sg13g2_o21ai_1
X_1413_ net756 net660 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_95_175 VPWR VGND sg13g2_fill_2
XFILLER_3_62 VPWR VGND sg13g2_decap_8
X_1344_ net751 net680 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
X_1275_ net194 net705 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
Xoutput484 net484 Tile_X0Y1_FrameData_O[27] VPWR VGND sg13g2_buf_1
Xoutput473 net473 Tile_X0Y1_FrameData_O[17] VPWR VGND sg13g2_buf_1
Xoutput495 net495 Tile_X0Y1_FrameData_O[8] VPWR VGND sg13g2_buf_1
Xoutput440 net440 Tile_X0Y0_W6BEG[1] VPWR VGND sg13g2_buf_1
Xoutput451 net451 Tile_X0Y0_WW4BEG[11] VPWR VGND sg13g2_buf_1
Xoutput462 net462 Tile_X0Y0_WW4BEG[7] VPWR VGND sg13g2_buf_1
XFILLER_78_109 VPWR VGND sg13g2_decap_4
XFILLER_6_124 VPWR VGND sg13g2_fill_1
XFILLER_6_146 VPWR VGND sg13g2_fill_1
X_1060_ net795 net677 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_77_175 VPWR VGND sg13g2_fill_2
XFILLER_77_120 VPWR VGND sg13g2_fill_1
X_0913_ net809 net735 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
X_0844_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit4.Q net230
+ net154 net147 net148 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit6.Q
+ _0279_ VPWR VGND sg13g2_mux4_1
X_0775_ VGND VPWR _0026_ _0214_ _0216_ _0215_ sg13g2_a21oi_1
X_1189_ net756 net739 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
X_1327_ net764 net681 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
X_1258_ net758 net704 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
Xoutput270 net270 BM_SRAM17 VPWR VGND sg13g2_buf_1
XFILLER_74_22 VPWR VGND sg13g2_fill_1
XFILLER_59_164 VPWR VGND sg13g2_decap_8
Xoutput292 net292 BM_SRAM9 VPWR VGND sg13g2_buf_1
Xoutput281 net281 BM_SRAM27 VPWR VGND sg13g2_buf_1
X_0560_ VGND VPWR _0013_ _0116_ _0120_ _0119_ sg13g2_a21oi_1
X_0491_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit27.Q net12
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG5 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG1
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG6 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit26.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG10 VPWR VGND sg13g2_mux4_1
XFILLER_2_182 VPWR VGND sg13g2_decap_8
XFILLER_31_6 VPWR VGND sg13g2_fill_1
X_1112_ net785 net666 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
X_1043_ net811 net687 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_119_136 VPWR VGND sg13g2_decap_8
XFILLER_9_94 VPWR VGND sg13g2_fill_2
X_0758_ net144 net182 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit8.Q
+ _0200_ VPWR VGND sg13g2_mux2_1
X_0827_ _0263_ net148 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit0.Q
+ VPWR VGND sg13g2_nand2_1
X_0689_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit23.Q net638
+ _0168_ VPWR VGND Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit22.Q
+ sg13g2_nand3b_1
XFILLER_71_126 VPWR VGND sg13g2_fill_2
XFILLER_107_2 VPWR VGND sg13g2_fill_1
XFILLER_85_87 VPWR VGND sg13g2_fill_2
XFILLER_85_54 VPWR VGND sg13g2_fill_2
XFILLER_47_178 VPWR VGND sg13g2_fill_1
X_1592_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG9 net448 VPWR
+ VGND sg13g2_buf_1
X_1661_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG6 net515 VPWR
+ VGND sg13g2_buf_1
X_0612_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit20.Q net145
+ net164 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG15 _0077_
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit21.Q Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S1BEG3
+ VPWR VGND sg13g2_mux4_1
X_0474_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit30.Q net10
+ net23 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG3 net628 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit31.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG12 VPWR VGND sg13g2_mux4_1
X_0543_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit16.Q VPWR
+ _0105_ VGND _0103_ _0104_ sg13g2_o21ai_1
X_1026_ net793 net685 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_53_159 VPWR VGND sg13g2_fill_1
XFILLER_61_192 VPWR VGND sg13g2_fill_1
XFILLER_111_30 VPWR VGND sg13g2_fill_2
XFILLER_55_79 VPWR VGND sg13g2_fill_1
XFILLER_112_0 VPWR VGND sg13g2_fill_1
XFILLER_121_164 VPWR VGND sg13g2_decap_8
X_1713_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG2 net573 VPWR
+ VGND sg13g2_buf_1
XFILLER_112_131 VPWR VGND sg13g2_fill_1
X_0526_ _0093_ net38 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit31.Q
+ VPWR VGND sg13g2_nand2b_1
X_1575_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb0 net429 VPWR
+ VGND sg13g2_buf_1
X_1644_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S1BEG1 net498 VPWR
+ VGND sg13g2_buf_1
X_0457_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit30.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END3
+ net250 net117 net137 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit31.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG11 VPWR VGND sg13g2_mux4_1
X_0388_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit30.Q net53
+ net45 net63 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit31.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG0 VPWR VGND sg13g2_mux4_1
XFILLER_26_115 VPWR VGND sg13g2_fill_2
X_1009_ net809 net697 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_25_27 VPWR VGND sg13g2_fill_1
XFILLER_26_159 VPWR VGND sg13g2_fill_2
XFILLER_103_186 VPWR VGND sg13g2_fill_2
XFILLER_32_107 VPWR VGND sg13g2_fill_2
XFILLER_40_173 VPWR VGND sg13g2_fill_1
X_1360_ net765 net673 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_56_8 VPWR VGND sg13g2_fill_2
X_0311_ VPWR _0014_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit24.Q
+ VGND sg13g2_inv_1
Xinput181 Tile_X0Y1_EE4END[1] net181 VPWR VGND sg13g2_buf_1
X_1291_ net211 net694 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
Xinput192 Tile_X0Y1_FrameData[11] net192 VPWR VGND sg13g2_buf_1
Xinput170 Tile_X0Y1_E6END[6] net170 VPWR VGND sg13g2_buf_1
X_1489_ net807 net334 VPWR VGND sg13g2_buf_1
X_1558_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N4BEG0 net403 VPWR
+ VGND sg13g2_buf_1
X_0509_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit30.Q net66
+ net80 net54 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit31.Q
+ net269 VPWR VGND sg13g2_mux4_1
X_1627_ net197 net472 VPWR VGND sg13g2_buf_1
XFILLER_117_95 VPWR VGND sg13g2_decap_8
XFILLER_13_151 VPWR VGND sg13g2_decap_4
X_0791_ net143 net178 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit9.Q
+ _0230_ VPWR VGND sg13g2_mux2_1
X_0860_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit4.Q _0293_
+ _0294_ _0295_ VPWR VGND sg13g2_nor3_1
XFILLER_3_41 VPWR VGND sg13g2_decap_8
X_1343_ net750 net684 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
X_1412_ net755 net659 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
X_1274_ net195 net704 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
X_0989_ net802 net712 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
Xoutput441 net441 Tile_X0Y0_W6BEG[2] VPWR VGND sg13g2_buf_1
Xoutput452 net452 Tile_X0Y0_WW4BEG[12] VPWR VGND sg13g2_buf_1
Xoutput430 net430 Tile_X0Y0_W2BEGb[1] VPWR VGND sg13g2_buf_1
Xoutput485 net485 Tile_X0Y1_FrameData_O[28] VPWR VGND sg13g2_buf_1
Xoutput474 net474 Tile_X0Y1_FrameData_O[18] VPWR VGND sg13g2_buf_1
Xoutput496 net496 Tile_X0Y1_FrameData_O[9] VPWR VGND sg13g2_buf_1
Xoutput463 net463 Tile_X0Y0_WW4BEG[8] VPWR VGND sg13g2_buf_1
XFILLER_63_46 VPWR VGND sg13g2_decap_4
XFILLER_10_143 VPWR VGND sg13g2_fill_1
Xfanout690 net691 net690 VPWR VGND sg13g2_buf_1
X_0912_ net87 net734 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
X_0843_ net327 _0274_ _0278_ _0270_ _0036_ VPWR VGND sg13g2_a22oi_1
X_0774_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit13.Q VPWR
+ _0215_ VGND _0212_ _0213_ sg13g2_o21ai_1
X_1326_ net763 net681 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_83_157 VPWR VGND sg13g2_fill_2
X_1188_ net755 net738 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
X_1257_ net757 net704 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_3_139 VPWR VGND sg13g2_decap_8
Xoutput260 net260 ADDR_SRAM9 VPWR VGND sg13g2_buf_1
Xoutput271 net271 BM_SRAM18 VPWR VGND sg13g2_buf_1
Xoutput282 net282 BM_SRAM28 VPWR VGND sg13g2_buf_1
Xoutput293 net293 CLK_SRAM VPWR VGND sg13g2_buf_1
XFILLER_74_157 VPWR VGND sg13g2_fill_2
XFILLER_74_89 VPWR VGND sg13g2_fill_1
X_0490_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit25.Q net11
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG6 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG2
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG5 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit24.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG9 VPWR VGND sg13g2_mux4_1
XFILLER_2_161 VPWR VGND sg13g2_decap_8
X_1111_ net111 net666 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_80_138 VPWR VGND sg13g2_fill_2
X_1042_ net810 net686 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_48_90 VPWR VGND sg13g2_decap_8
XFILLER_119_115 VPWR VGND sg13g2_decap_8
X_0688_ _0165_ VPWR net252 VGND Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit21.Q
+ _0167_ sg13g2_o21ai_1
X_0757_ _0198_ VPWR _0199_ VGND _0023_ _0159_ sg13g2_o21ai_1
X_0826_ _0262_ net147 _0035_ VPWR VGND sg13g2_nand2_1
X_1309_ net779 net692 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_44_26 VPWR VGND sg13g2_fill_2
XFILLER_118_192 VPWR VGND sg13g2_fill_1
XFILLER_118_181 VPWR VGND sg13g2_decap_8
XFILLER_114_4 VPWR VGND sg13g2_fill_2
XFILLER_70_182 VPWR VGND sg13g2_fill_2
X_1591_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG8 net447 VPWR
+ VGND sg13g2_buf_1
X_1660_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG5 net514 VPWR
+ VGND sg13g2_buf_1
X_0542_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit15.Q VPWR
+ _0104_ VGND Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit14.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG12 sg13g2_o21ai_1
X_0611_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit18.Q net144
+ net163 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG14 _0070_
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit19.Q Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S1BEG2
+ VPWR VGND sg13g2_mux4_1
X_0473_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit14.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END3
+ net250 net117 net137 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit15.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG3 VPWR VGND sg13g2_mux4_1
XFILLER_38_179 VPWR VGND sg13g2_fill_2
XFILLER_53_105 VPWR VGND sg13g2_fill_1
X_1025_ net792 net685 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
X_0809_ VGND VPWR _0239_ _0241_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S4BEG2
+ _0246_ sg13g2_a21oi_1
XFILLER_29_157 VPWR VGND sg13g2_fill_2
XFILLER_29_179 VPWR VGND sg13g2_fill_2
XFILLER_121_143 VPWR VGND sg13g2_decap_8
XFILLER_96_21 VPWR VGND sg13g2_fill_1
X_1712_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG1 net572 VPWR
+ VGND sg13g2_buf_1
XFILLER_6_52 VPWR VGND sg13g2_fill_2
X_1643_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S1BEG0 net497 VPWR
+ VGND sg13g2_buf_1
X_0525_ net46 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit30.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit31.Q _0092_ VPWR
+ VGND sg13g2_nor3_1
X_1574_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG7 net428 VPWR
+ VGND sg13g2_buf_1
X_0456_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit12.Q net13
+ net27 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG12 net626
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit13.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG3
+ VPWR VGND sg13g2_mux4_1
X_0387_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit28.Q net37
+ net63 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG15 _0073_
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit29.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1BEG3
+ VPWR VGND sg13g2_mux4_1
X_1008_ net808 net700 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_66_46 VPWR VGND sg13g2_fill_2
XFILLER_82_45 VPWR VGND sg13g2_fill_2
X_0310_ VPWR _0013_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit21.Q
+ VGND sg13g2_inv_1
Xinput160 Tile_X0Y1_E2MID[6] net160 VPWR VGND sg13g2_buf_1
Xinput182 Tile_X0Y1_EE4END[2] net182 VPWR VGND sg13g2_buf_1
X_1290_ net758 net694 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
Xinput171 Tile_X0Y1_E6END[7] net171 VPWR VGND sg13g2_buf_1
Xinput193 Tile_X0Y1_FrameData[12] net193 VPWR VGND sg13g2_buf_1
XFILLER_82_2 VPWR VGND sg13g2_fill_1
XFILLER_16_182 VPWR VGND sg13g2_fill_1
X_1626_ net775 net471 VPWR VGND sg13g2_buf_1
X_0508_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit28.Q net37
+ net79 net72 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG15 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit29.Q
+ net319 VPWR VGND sg13g2_mux4_1
X_1488_ net808 net333 VPWR VGND sg13g2_buf_1
X_0439_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit12.Q net13
+ net22 net628 net626 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit13.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG3 VPWR VGND sg13g2_mux4_1
X_1557_ Tile_X0Y0_IHP_SRAM_top.N4BEG_outbuf_11.A net402 VPWR VGND sg13g2_buf_1
XFILLER_14_108 VPWR VGND sg13g2_fill_2
XFILLER_117_74 VPWR VGND sg13g2_decap_8
XFILLER_89_130 VPWR VGND sg13g2_fill_1
XFILLER_77_78 VPWR VGND sg13g2_decap_4
XFILLER_61_7 VPWR VGND sg13g2_fill_2
X_0790_ _0228_ VPWR _0229_ VGND _0029_ _0160_ sg13g2_o21ai_1
XFILLER_95_144 VPWR VGND sg13g2_fill_1
X_1342_ net780 net680 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_3_97 VPWR VGND sg13g2_decap_4
XFILLER_3_20 VPWR VGND sg13g2_decap_8
X_1411_ net754 net659 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
X_1273_ net196 net704 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
X_0988_ net791 net710 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
Xoutput486 net486 Tile_X0Y1_FrameData_O[29] VPWR VGND sg13g2_buf_1
Xoutput475 net475 Tile_X0Y1_FrameData_O[19] VPWR VGND sg13g2_buf_1
Xoutput442 net442 Tile_X0Y0_W6BEG[3] VPWR VGND sg13g2_buf_1
Xoutput464 net464 Tile_X0Y0_WW4BEG[9] VPWR VGND sg13g2_buf_1
Xoutput453 net453 Tile_X0Y0_WW4BEG[13] VPWR VGND sg13g2_buf_1
Xoutput431 net431 Tile_X0Y0_W2BEGb[2] VPWR VGND sg13g2_buf_1
X_1609_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG14 net454 VPWR
+ VGND sg13g2_buf_1
Xoutput420 net420 Tile_X0Y0_W1BEG[3] VPWR VGND sg13g2_buf_1
XFILLER_103_32 VPWR VGND sg13g2_fill_1
Xoutput497 net497 Tile_X0Y1_S1BEG[0] VPWR VGND sg13g2_buf_1
XFILLER_27_200 VPWR VGND sg13g2_fill_1
XFILLER_63_25 VPWR VGND sg13g2_decap_4
XFILLER_92_136 VPWR VGND sg13g2_fill_2
XFILLER_77_199 VPWR VGND sg13g2_fill_2
XFILLER_77_177 VPWR VGND sg13g2_fill_1
Xfanout691 Tile_X0Y1_FrameStrobe[5] net691 VPWR VGND sg13g2_buf_1
Xfanout680 net681 net680 VPWR VGND sg13g2_buf_1
X_0911_ net88 net734 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
X_0842_ VGND VPWR _0035_ _0277_ _0278_ _0036_ sg13g2_a21oi_1
X_0773_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG7 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG11
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit11.Q _0214_ VPWR
+ VGND sg13g2_mux2_1
XFILLER_83_114 VPWR VGND sg13g2_fill_1
XFILLER_68_177 VPWR VGND sg13g2_fill_2
XFILLER_68_122 VPWR VGND sg13g2_decap_8
X_1325_ net762 net683 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
X_1256_ net190 net714 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
X_1187_ net754 net738 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_59_122 VPWR VGND sg13g2_decap_4
XFILLER_3_118 VPWR VGND sg13g2_decap_8
Xoutput261 net261 BM_SRAM0 VPWR VGND sg13g2_buf_1
Xoutput272 net272 BM_SRAM19 VPWR VGND sg13g2_buf_1
Xoutput283 net283 BM_SRAM29 VPWR VGND sg13g2_buf_1
Xoutput294 net294 DIN_SRAM0 VPWR VGND sg13g2_buf_1
XFILLER_114_75 VPWR VGND sg13g2_fill_2
XFILLER_2_140 VPWR VGND sg13g2_decap_8
X_1110_ net112 net666 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_65_125 VPWR VGND sg13g2_fill_1
X_1041_ net809 net686 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
X_0825_ VGND VPWR net241 _0035_ _0261_ _0260_ sg13g2_a21oi_1
X_0687_ VGND VPWR net147 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit20.Q
+ _0167_ _0166_ sg13g2_a21oi_1
X_0756_ VPWR _0198_ _0197_ VGND sg13g2_inv_1
XFILLER_71_128 VPWR VGND sg13g2_fill_1
X_1308_ net778 net695 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
X_1239_ net198 net714 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_56_103 VPWR VGND sg13g2_fill_1
XFILLER_100_44 VPWR VGND sg13g2_fill_2
XFILLER_118_160 VPWR VGND sg13g2_decap_8
XFILLER_85_12 VPWR VGND sg13g2_fill_2
XFILLER_69_79 VPWR VGND sg13g2_decap_4
XFILLER_85_89 VPWR VGND sg13g2_fill_1
XFILLER_18_61 VPWR VGND sg13g2_fill_1
XFILLER_109_171 VPWR VGND sg13g2_fill_1
X_0541_ net631 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit14.Q
+ _0103_ VPWR VGND sg13g2_nor2b_1
X_0472_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit28.Q net18
+ net22 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG4 net626 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit29.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG11 VPWR VGND sg13g2_mux4_1
X_1590_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG7 net446 VPWR
+ VGND sg13g2_buf_1
X_0610_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit16.Q net143
+ net173 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG13 _0063_
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit17.Q Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S1BEG1
+ VPWR VGND sg13g2_mux4_1
X_1024_ net790 net685 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
X_0808_ VGND VPWR _0032_ _0244_ _0246_ _0245_ sg13g2_a21oi_1
X_0739_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit3.Q VPWR
+ _0183_ VGND Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit2.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG12 sg13g2_o21ai_1
XFILLER_111_32 VPWR VGND sg13g2_fill_1
XFILLER_37_191 VPWR VGND sg13g2_fill_2
XFILLER_121_122 VPWR VGND sg13g2_decap_8
X_1642_ net757 net489 VPWR VGND sg13g2_buf_1
X_1711_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG0 net565 VPWR
+ VGND sg13g2_buf_1
XFILLER_112_166 VPWR VGND sg13g2_fill_2
X_0524_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit28.Q net37
+ net79 net72 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG15 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit29.Q
+ net286 VPWR VGND sg13g2_mux4_1
X_0455_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit0.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END0
+ net247 net114 net134 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit1.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG12 VPWR VGND sg13g2_mux4_1
X_1573_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG6 net427 VPWR
+ VGND sg13g2_buf_1
X_1007_ net807 net700 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
X_0386_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit6.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END3
+ net250 net117 net137 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit7.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG15 VPWR VGND sg13g2_mux4_1
XFILLER_34_161 VPWR VGND sg13g2_fill_1
XFILLER_103_100 VPWR VGND sg13g2_fill_2
XFILLER_103_188 VPWR VGND sg13g2_fill_1
Xinput161 Tile_X0Y1_E2MID[7] net161 VPWR VGND sg13g2_buf_1
Xinput183 Tile_X0Y1_EE4END[3] net183 VPWR VGND sg13g2_buf_1
Xinput150 Tile_X0Y1_E2END[4] net150 VPWR VGND sg13g2_buf_1
Xinput172 Tile_X0Y1_E6END[8] net172 VPWR VGND sg13g2_buf_1
Xinput194 Tile_X0Y1_FrameData[13] net194 VPWR VGND sg13g2_buf_1
X_1625_ net776 net470 VPWR VGND sg13g2_buf_1
X_1556_ Tile_X0Y0_IHP_SRAM_top.N4BEG_outbuf_10.A net401 VPWR VGND sg13g2_buf_1
X_1487_ net809 net332 VPWR VGND sg13g2_buf_1
X_0507_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit26.Q net36
+ net78 net71 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG14 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit27.Q
+ net318 VPWR VGND sg13g2_mux4_1
X_0369_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit28.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit29.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END2 _0065_ VPWR VGND sg13g2_nor3_1
X_0438_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit10.Q net12
+ net21 net629 net625 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit11.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG2 VPWR VGND sg13g2_mux4_1
XFILLER_117_53 VPWR VGND sg13g2_decap_8
XFILLER_9_146 VPWR VGND sg13g2_fill_1
XFILLER_9_135 VPWR VGND sg13g2_decap_8
XFILLER_9_113 VPWR VGND sg13g2_fill_1
XFILLER_26_61 VPWR VGND sg13g2_fill_2
X_1410_ net218 net662 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
X_1341_ net779 net680 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_3_76 VPWR VGND sg13g2_decap_8
X_1272_ net197 net707 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
X_0987_ net788 net711 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
Xoutput410 net410 Tile_X0Y0_N4BEG[4] VPWR VGND sg13g2_buf_1
Xoutput487 net487 Tile_X0Y1_FrameData_O[2] VPWR VGND sg13g2_buf_1
Xoutput476 net476 Tile_X0Y1_FrameData_O[1] VPWR VGND sg13g2_buf_1
Xoutput465 net465 Tile_X0Y1_FrameData_O[0] VPWR VGND sg13g2_buf_1
X_1608_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG13 net453 VPWR
+ VGND sg13g2_buf_1
Xoutput443 net443 Tile_X0Y0_W6BEG[4] VPWR VGND sg13g2_buf_1
Xoutput454 net454 Tile_X0Y0_WW4BEG[14] VPWR VGND sg13g2_buf_1
Xoutput432 net432 Tile_X0Y0_W2BEGb[3] VPWR VGND sg13g2_buf_1
Xoutput421 net421 Tile_X0Y0_W2BEG[0] VPWR VGND sg13g2_buf_1
X_1539_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb1 net393 VPWR
+ VGND sg13g2_buf_1
Xoutput498 net498 Tile_X0Y1_S1BEG[1] VPWR VGND sg13g2_buf_1
Xfanout670 net672 net670 VPWR VGND sg13g2_buf_1
Xfanout681 net684 net681 VPWR VGND sg13g2_buf_1
Xfanout692 net693 net692 VPWR VGND sg13g2_buf_1
X_0910_ net806 net737 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
X_0841_ VGND VPWR Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit1.Q
+ _0276_ _0275_ _0002_ _0277_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit2.Q
+ sg13g2_a221oi_1
X_0772_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit12.Q VPWR
+ _0213_ VGND Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit11.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG15 sg13g2_o21ai_1
XFILLER_68_112 VPWR VGND sg13g2_fill_2
XFILLER_68_101 VPWR VGND sg13g2_decap_8
XFILLER_83_159 VPWR VGND sg13g2_fill_1
X_1324_ net761 net683 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
X_1186_ net753 net740 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
X_1255_ net770 net715 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_58_26 VPWR VGND sg13g2_fill_2
XFILLER_58_15 VPWR VGND sg13g2_decap_8
Xoutput251 net251 ADDR_SRAM0 VPWR VGND sg13g2_buf_1
Xoutput262 net262 BM_SRAM1 VPWR VGND sg13g2_buf_1
Xoutput273 net273 BM_SRAM2 VPWR VGND sg13g2_buf_1
Xoutput284 net284 BM_SRAM3 VPWR VGND sg13g2_buf_1
Xoutput295 net295 DIN_SRAM1 VPWR VGND sg13g2_buf_1
XFILLER_74_159 VPWR VGND sg13g2_fill_1
X_1040_ net808 net685 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_2_196 VPWR VGND sg13g2_fill_1
XFILLER_48_81 VPWR VGND sg13g2_decap_4
X_0755_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit9.Q VPWR
+ _0197_ VGND net163 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit8.Q
+ sg13g2_o21ai_1
X_0824_ VGND VPWR _0260_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit2.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit1.Q sg13g2_or2_1
X_0686_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit20.Q net155
+ _0166_ VPWR VGND sg13g2_nor2b_1
X_1169_ net766 net738 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
X_1307_ net777 net693 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
X_1238_ net199 net717 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_60_49 VPWR VGND sg13g2_fill_1
XFILLER_114_6 VPWR VGND sg13g2_fill_1
XFILLER_85_68 VPWR VGND sg13g2_fill_2
XFILLER_85_35 VPWR VGND sg13g2_fill_2
XFILLER_62_129 VPWR VGND sg13g2_decap_8
X_0540_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG4 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG8
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit14.Q _0102_ VPWR
+ VGND sg13g2_mux2_1
X_0471_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit16.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END0
+ net247 net114 net134 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit17.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG4 VPWR VGND sg13g2_mux4_1
X_1023_ net789 net685 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
X_0738_ _0019_ _0043_ _0182_ VPWR VGND sg13g2_nor2_1
X_0807_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit14.Q VPWR
+ _0245_ VGND _0242_ _0243_ sg13g2_o21ai_1
X_0669_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit26.Q net243
+ net138 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG11 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG15
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit27.Q Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG0
+ VPWR VGND sg13g2_mux4_1
XFILLER_121_101 VPWR VGND sg13g2_decap_8
XFILLER_96_67 VPWR VGND sg13g2_fill_2
XFILLER_29_94 VPWR VGND sg13g2_fill_2
X_1572_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG5 net426 VPWR
+ VGND sg13g2_buf_1
XFILLER_61_92 VPWR VGND sg13g2_fill_2
XFILLER_61_81 VPWR VGND sg13g2_fill_1
X_1641_ net758 net488 VPWR VGND sg13g2_buf_1
XFILLER_6_54 VPWR VGND sg13g2_fill_1
X_1710_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG11 net555 VPWR
+ VGND sg13g2_buf_1
X_0523_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit26.Q net36
+ net78 net71 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG14 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit27.Q
+ net285 VPWR VGND sg13g2_mux4_1
X_0454_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit10.Q net12
+ net26 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG13 net625
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit11.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG2
+ VPWR VGND sg13g2_mux4_1
X_0385_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit17.Q net145
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG15 net171 _0077_
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit16.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END3
+ VPWR VGND sg13g2_mux4_1
X_1006_ net806 net698 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_110_0 VPWR VGND sg13g2_fill_2
Xinput140 Tile_X0Y0_S4END[6] net140 VPWR VGND sg13g2_buf_1
Xinput151 Tile_X0Y1_E2END[5] net151 VPWR VGND sg13g2_buf_1
Xinput162 Tile_X0Y1_E6END[0] net162 VPWR VGND sg13g2_buf_1
Xinput184 Tile_X0Y1_EE4END[4] net184 VPWR VGND sg13g2_buf_1
Xinput173 Tile_X0Y1_E6END[9] net173 VPWR VGND sg13g2_buf_1
Xinput195 Tile_X0Y1_FrameData[14] net195 VPWR VGND sg13g2_buf_1
X_0506_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit24.Q net35
+ net77 net70 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG13 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit25.Q
+ net316 VPWR VGND sg13g2_mux4_1
X_1555_ Tile_X0Y0_IHP_SRAM_top.N4BEG_outbuf_9.A net415 VPWR VGND sg13g2_buf_1
X_1624_ net194 net469 VPWR VGND sg13g2_buf_1
X_1486_ net810 net331 VPWR VGND sg13g2_buf_1
X_0368_ _0064_ net116 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit28.Q
+ VPWR VGND sg13g2_nand2b_1
X_0437_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit8.Q net11
+ net20 net630 net624 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit9.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG1 VPWR VGND sg13g2_mux4_1
X_0299_ VPWR _0002_ net128 VGND sg13g2_inv_1
XFILLER_52_39 VPWR VGND sg13g2_fill_2
XFILLER_117_32 VPWR VGND sg13g2_decap_8
XFILLER_89_198 VPWR VGND sg13g2_fill_2
XFILLER_77_47 VPWR VGND sg13g2_fill_1
X_1340_ net778 net680 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_95_157 VPWR VGND sg13g2_fill_1
XFILLER_3_55 VPWR VGND sg13g2_decap_8
X_1271_ net198 net707 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
Xoutput400 net400 Tile_X0Y0_N4BEG[0] VPWR VGND sg13g2_buf_1
Xoutput411 net411 Tile_X0Y0_N4BEG[5] VPWR VGND sg13g2_buf_1
X_0986_ net108 net710 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
Xoutput488 net488 Tile_X0Y1_FrameData_O[30] VPWR VGND sg13g2_buf_1
Xoutput477 net477 Tile_X0Y1_FrameData_O[20] VPWR VGND sg13g2_buf_1
Xoutput466 net466 Tile_X0Y1_FrameData_O[10] VPWR VGND sg13g2_buf_1
X_1607_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG12 net452 VPWR
+ VGND sg13g2_buf_1
Xoutput444 net444 Tile_X0Y0_W6BEG[5] VPWR VGND sg13g2_buf_1
Xoutput455 net455 Tile_X0Y0_WW4BEG[15] VPWR VGND sg13g2_buf_1
Xoutput433 net433 Tile_X0Y0_W2BEGb[4] VPWR VGND sg13g2_buf_1
Xoutput422 net422 Tile_X0Y0_W2BEG[1] VPWR VGND sg13g2_buf_1
Xoutput499 net499 Tile_X0Y1_S1BEG[2] VPWR VGND sg13g2_buf_1
X_1469_ net192 net642 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
X_1538_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb0 net392 VPWR
+ VGND sg13g2_buf_1
XFILLER_92_138 VPWR VGND sg13g2_fill_1
Xfanout671 net672 net671 VPWR VGND sg13g2_buf_1
Xfanout682 net684 net682 VPWR VGND sg13g2_buf_1
Xfanout693 net695 net693 VPWR VGND sg13g2_buf_1
Xfanout660 net661 net660 VPWR VGND sg13g2_buf_1
X_0840_ net149 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit1.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit2.Q _0276_ VPWR
+ VGND sg13g2_nor3_1
X_0771_ _0025_ _0080_ _0212_ VPWR VGND sg13g2_nor2_1
XFILLER_5_183 VPWR VGND sg13g2_fill_2
X_1323_ net760 net682 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
X_1254_ net212 net717 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
X_1185_ net752 net741 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
X_0969_ net800 net710 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
Xoutput252 net252 ADDR_SRAM1 VPWR VGND sg13g2_buf_1
XFILLER_74_138 VPWR VGND sg13g2_fill_2
Xoutput296 net296 DIN_SRAM10 VPWR VGND sg13g2_buf_1
Xoutput274 net274 BM_SRAM20 VPWR VGND sg13g2_buf_1
Xoutput263 net263 BM_SRAM10 VPWR VGND sg13g2_buf_1
Xoutput285 net285 BM_SRAM30 VPWR VGND sg13g2_buf_1
XFILLER_114_77 VPWR VGND sg13g2_fill_1
XFILLER_2_175 VPWR VGND sg13g2_decap_8
XFILLER_119_129 VPWR VGND sg13g2_decap_8
X_0754_ VGND VPWR _0189_ _0191_ Tile_X0Y0_IHP_SRAM_top.N4BEG_outbuf_9.A _0196_ sg13g2_a21oi_1
X_0685_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit21.Q _0078_
+ _0165_ VPWR VGND Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit20.Q
+ sg13g2_nand3b_1
X_0823_ _0259_ net229 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit0.Q
+ VPWR VGND sg13g2_nand2_1
X_1306_ net776 net695 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_71_119 VPWR VGND sg13g2_decap_8
X_1099_ net803 net663 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
X_1168_ net206 net742 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
X_1237_ net200 net717 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_100_46 VPWR VGND sg13g2_fill_1
XFILLER_47_116 VPWR VGND sg13g2_fill_2
X_0470_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit26.Q net17
+ net21 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG5 net625 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit27.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG10 VPWR VGND sg13g2_mux4_1
X_1022_ net813 net699 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
X_0668_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit24.Q net25
+ net9 _0161_ _0043_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit25.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG15 VPWR VGND sg13g2_mux4_1
X_0737_ VGND VPWR _0020_ _0180_ _0181_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit4.Q
+ sg13g2_a21oi_1
X_0806_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG6 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG10
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit12.Q _0244_ VPWR
+ VGND sg13g2_mux2_1
X_0599_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit29.Q VPWR
+ _0154_ VGND _0152_ _0153_ sg13g2_o21ai_1
XFILLER_71_27 VPWR VGND sg13g2_fill_1
XFILLER_52_196 VPWR VGND sg13g2_fill_1
XFILLER_121_157 VPWR VGND sg13g2_decap_8
X_1571_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG4 net425 VPWR
+ VGND sg13g2_buf_1
X_0522_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit24.Q net35
+ net77 net70 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG13 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit25.Q
+ net283 VPWR VGND sg13g2_mux4_1
XFILLER_6_99 VPWR VGND sg13g2_decap_4
X_1640_ net760 net486 VPWR VGND sg13g2_buf_1
XFILLER_112_168 VPWR VGND sg13g2_fill_1
X_0453_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit8.Q net11
+ net24 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG14 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG6
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit9.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG1
+ VPWR VGND sg13g2_mux4_1
X_0384_ VGND VPWR _0076_ _0075_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit31.Q
+ _0007_ _0077_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit30.Q
+ sg13g2_a221oi_1
X_1005_ net805 net698 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_34_141 VPWR VGND sg13g2_fill_2
XFILLER_103_102 VPWR VGND sg13g2_fill_1
XFILLER_17_119 VPWR VGND sg13g2_fill_1
XFILLER_40_199 VPWR VGND sg13g2_fill_2
XFILLER_103_0 VPWR VGND sg13g2_fill_2
Xinput141 Tile_X0Y0_S4END[7] net141 VPWR VGND sg13g2_buf_1
Xinput130 Tile_X0Y0_S2MID[4] net130 VPWR VGND sg13g2_buf_1
Xinput174 Tile_X0Y1_EE4END[0] net174 VPWR VGND sg13g2_buf_1
Xinput152 Tile_X0Y1_E2END[6] net152 VPWR VGND sg13g2_buf_1
Xinput185 Tile_X0Y1_EE4END[5] net185 VPWR VGND sg13g2_buf_1
Xinput163 Tile_X0Y1_E6END[10] net163 VPWR VGND sg13g2_buf_1
XFILLER_48_200 VPWR VGND sg13g2_fill_1
Xinput196 Tile_X0Y1_FrameData[15] net196 VPWR VGND sg13g2_buf_1
XFILLER_31_133 VPWR VGND sg13g2_fill_2
XFILLER_56_93 VPWR VGND sg13g2_fill_2
X_1485_ net811 net330 VPWR VGND sg13g2_buf_1
XFILLER_98_133 VPWR VGND sg13g2_fill_1
XFILLER_98_111 VPWR VGND sg13g2_fill_1
X_0436_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit6.Q net10
+ net19 net631 net623 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit7.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG0 VPWR VGND sg13g2_mux4_1
X_0505_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit22.Q net34
+ net76 net69 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG12 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit23.Q
+ net315 VPWR VGND sg13g2_mux4_1
X_1554_ Tile_X0Y0_IHP_SRAM_top.N4BEG_outbuf_8.A net414 VPWR VGND sg13g2_buf_1
XFILLER_39_200 VPWR VGND sg13g2_fill_1
X_1623_ net193 net468 VPWR VGND sg13g2_buf_1
.ends

